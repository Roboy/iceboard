// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Oct 29 10:19:13 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    inout PIN_9 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    inout PIN_10 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    inout PIN_11 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_1, PIN_2_c_0, PIN_6_c_0, PIN_7_c_1, 
        PIN_8_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, PIN_22_c, 
        PIN_23_c;
    wire [31:0]communication_counter;   // verilog/TinyFPGA_B.v(67[9:30])
    wire [23:0]color;   // verilog/TinyFPGA_B.v(68[12:17])
    
    wire blink, hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(151[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(152[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(189[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(190[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(191[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(192[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(193[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(194[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(196[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(197[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(198[22:35])
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(200[22:34])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(225[22:33])
    
    wire n28485, n5869, n5868, n5867, n5866, n5865;
    wire [7:0]color_23__N_164;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n28484, n1169, n1163, n5864, n5863, n5886, n5885, n5884, 
        n1158, n1157, n1156, n1155, n41522, n672, n671, n670, 
        n669, n668, blink_N_255;
    wire [22:0]pwm_setpoint_22__N_57;
    
    wire PIN_13_N_105, n5883, n5882, n5881, n41799;
    wire [31:0]motor_state_23__N_106;
    wire [24:0]displacement_23__N_229;
    wire [23:0]displacement_23__N_80;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n5880, n5879, n5878, n28483, n28482, n28481;
    wire [3:0]state_3__N_362;
    wire [31:0]one_wire_N_513;
    
    wire n1251, n28480, n5847, n5839, n15573, n2, n5870, n63, 
        n28479, n5909, n2954, n2953, n2952, n4385, n98, n99, 
        n2718, n2720, n2716, n2714, n2712, n2710, n2708, n2906_adj_4319, 
        n5845, n15, n17, n13, n24, n19, n20, n8, n33325, n15_adj_4320, 
        n2951, n2950, n1154, n1153, n47, n46, n4591, n28478, 
        n15_adj_4321, n16754, n4613, n6, n87, n90, n89, n88, 
        n86, n85, n84, n60, n91, n92, n43, n2949, n2948, n2947, 
        n2946, n2945, n18, n2944, n2943, n2942, n2941, n42, 
        n15_adj_4322, n1152, n1151, n96, n40, n39, n28477, n5, 
        n38, n97, n95, n94, n93, n83, n82, n81, n80, n79, 
        n66, n65, n2914, n2913, n2912, n2911, n6_adj_4323, n2910, 
        n2909, n2908, n2907, n2906, n2905, n2904, n2903, n2902, 
        n2901, n2900, n2899, n2898, n2897, n2896, n2895, n2894, 
        n2893, n2892, n2891, n63_adj_4324, n28476, n667, n666, 
        n665, n664, n663, n662, n661, n660, n659, n658, n657, 
        n656, n655, n654, n653, n652, n651, n650, n649, n648, 
        n15564, n15561, n31, n1125, n1124, n1123, n1122, n5985, 
        n5984, n5983, n5982, n6012, n6011, n6010, n6009, n6008, 
        n6007, n6006, n6005, n6004, n6003, n6032, n6031, n6030, 
        n6029, n6028, n6027, n1121, n33327, n64, n1120, n78;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n5844, n5843, n4, n5892, n5922, n5921, n5920, n4_adj_4325, 
        n5919, n5918, n77, n75, n73, n72, n71, n68, n1257, 
        n10, n3, n4_adj_4326, n5_adj_4327, n6_adj_4328, n7, n8_adj_4329, 
        n9, n10_adj_4330, n11, n12, n13_adj_4331, n14, n15_adj_4332, 
        n16, n17_adj_4333, n18_adj_4334, n19_adj_4335, n20_adj_4336, 
        n21, n22, n23, n24_adj_4337, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    
    wire n15558, n15555, n15549;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n5986, n5987, n5988, n5989, n5990, n5991, n5992, n28475, 
        n122, n28474;
    wire [31:0]\FRAME_MATCHER.state_31__N_2426 ;
    
    wire n15546, n28473, n28472, n28471, n28470, n28469, n28468, 
        n28467, n28466, n15535, n61, n59, n70, n28465, n28464, 
        n28463, n28462, n28461, n35555, n737, n41223, n28460, 
        n42332, n28459, n26602, n35315, n26612, n28458, n28650, 
        n34, n28649, n28648, n28647, n28646, n15_adj_4338, n28645, 
        n27989, n15530, n28644, n28643, n27988, n31_adj_4339, n30, 
        n41217, n28457, n28456, n28, n15526, n15522, n22_adj_4340, 
        n28642, n28455, n21_adj_4341, n41215, n28641, n28454, n28640, 
        n28639, n27987, n28638, n28453, n28637, n28636, n28635, 
        n28634, n28452, n28451, n28450, n28449, n28633, n28448, 
        n35558, n15517, n28447, n28446, n28445, n28444, n28443, 
        n28442, n28441, n28440, n28439, n28438, n28632, n27986, 
        n27985, n40570, n24014, n35615, n27984, n41203, n41201, 
        n41199, n28437, n27983, n28436, n28631, n27982, n27981, 
        n28630, n28435, n2_adj_4342, n28629, n28628, n15508, n28434, 
        n28627, n28433, n28626, n28432, n28625, n28431, n28624, 
        n28623, n28430, n28622, n41191, n15504, n15501, n28429, 
        n15498, n15494, n28621, n28620, n35665, n28619, n28618, 
        n28617, n28428, n15491, n27980, n28427, n69, n67, n28616, 
        n5935, n5934, n5933, n5932, n41786, n2855, n41772, n41189, 
        n28426, n28425, n41185, n28424, n41183, n28423, n27979, 
        n5930, n5929, n5_adj_4343, n11_adj_4344, n12_adj_4345, n27978, 
        n28615, n28422, n28614, n18962, n28421, n28613, n28420, 
        n28612, n28611, n28610, n15454, n41173, n28609, n28608, 
        n28419, n28607, n28418, n28606, n29, n28605, n28604, n28417, 
        n28416, n27977, n27976, n27975, n27974, n28415, n28414, 
        n28603, n41795, n28602, n28601, n28413, n28600, n28412, 
        n30_adj_4346, n28599, n28411, n30_adj_4347, n29_adj_4348, 
        n41620, n35528, n28_adj_4349, n27, n28598, n28410, n18_adj_4350, 
        n41169, n19_adj_4351, n18_adj_4352, n12_adj_4353, n41542, 
        n15_adj_4354, n41152, n5927, n5926, n28409, n28408, n28597, 
        n28407, n16772, n28406, n28405, \FRAME_MATCHER.i_31__N_2386 , 
        \FRAME_MATCHER.i_31__N_2390 , n17303, n17302, n41546, n17301, 
        n17300, n17299, n17298, n17297, n17295, n17294, n17293, 
        n17292, n17291, n17290, n17289, n17288, n17287, n17286, 
        n17285, n17284, n17283, n17282, n17281, n17280, n17279, 
        n17278, n17277, n17276, n17275, n17274, n17273, n17272, 
        n17271, n17270, n17269, n17268, n17267, n17266, n17265, 
        n17264, n17263, n17262, n17261, n17260, n17259, n17258, 
        n17257, n17256, n17255, n17254, n17253, n17252, n17251, 
        n17250, n17249, n17248, n17247, n17246, n17245, n17244, 
        n17243, n17242, n17241, n17240, n17239, n17238, n17237, 
        n17236, n17235, n17234, n17233, n17232, n17231, n17230, 
        n17229, n17228, n17227, n17226, n17225, n17224, n17223, 
        n17222, n17221, n17220, n17219, n17218, n17217, n17216, 
        n17215, n17214, n17213, n17212, n17211, n17210, n17209, 
        n17208, n17207, n17206, n17205, n17204, n17203, n17202, 
        n17201, n17200, n17199, n17198, n17197, n17196, n17195, 
        n17194, n17193, n17192, n17191, n17190, n17189, n17188, 
        n17187, n17186, n17185, n17184, n17183, n17182, n17181, 
        n17180, n17179, n17178, n17177, n17176, n17175, n17174, 
        n17173, n17172, n17171, n17170, n17169, n17165, n17164, 
        n17163, n17162, n17161, n17160, n17159, n17158, n17157, 
        n17155, n17154, n17153, n17151, n17149, n17147, n17146, 
        n17145, n17144, n17143, n17142, n17141, n17139, n17138, 
        n17137, n17136, n17135, n17134, n17133, n17132, n17131, 
        n17130, n17129, n17128, n17127, n17126, n17125, n17124, 
        n17123, n17122, n17121, n17120, n17119, n17118, n17117, 
        n17116, n17115, n17114, n17113, n17112, n17111, n17110, 
        n17109, n17108, n17107, n17106, n17105, n17104, n17103, 
        n17102, n17101, n17100, n17099, n17098, n17097, n17096, 
        n17095, n17094, n558, n14_adj_4355, n534, n533, n6048, 
        n6049, n6050, n6051, n6052, n6025, n6026, n511, n510, 
        n1085, n41784, n1382, n1058, n1057, n1056, n1055, n1054, 
        n1053, n1052, n5831, n5830, n5829, n5828, n5827, n5860, 
        n393, n392, n1358, n1357, n1356, n1355, n1354, n1353, 
        n17093, n369, n1025, n1024, n1023, n1022, n1352, n1351, 
        n1350, n1349, n17092, n17091, n17090, n17089, n17088, 
        n17087, n17086, n17085, n17084, n17083, n17082, n17081, 
        n17080, n17079, n17078, n17077, n1021, n4_adj_4356, n28404, 
        n28596, n28403, n33975, n28595, n28402, n28401, n28400, 
        n22_adj_4357, n25_adj_4358, n28594, n28593, n9_adj_4359, n5840, 
        n5841, n28592, n28591, n28590, n28589, n28399, n28588, 
        n28398, n28397, n28587, n28396, n35536, n4315, n4314, 
        n4313, n4312, n4311, n4310, n4309, n4308, n4307, n4306, 
        n4305, n4304, n4303, n4302, n4301, n4300, n4299, n4298, 
        n4297, n4296, n4295, n4294, n4293, n4292, n986, n5874, 
        n5873, n5872, n24_adj_4360, n35627, n21_adj_4361, n20_adj_4362, 
        n17_adj_4363, n42326, n17076, n17075, n17074, n17072, n17071, 
        n17070, n17069, n17068, n17067, n17066, n17065, n17064, 
        n17063, n17062, n17061, n17060, n17059, n17058, n17057, 
        n17056, n17055, n17054, n17053, n17052, n17051, n17050, 
        n17049, n11_adj_4364, quadA_debounced, quadB_debounced, count_enable, 
        n53, n54, n56, n57, n58, n55, n62, n10_adj_4365, n28586, 
        n9_adj_4366, n6_adj_4367, n6_adj_4368, n8_adj_4369, n7_adj_4370, 
        n249, n248, n6_adj_4371, n28585, quadA_debounced_adj_4372, 
        quadB_debounced_adj_4373, count_enable_adj_4374, n17048, n17047, 
        n42325, n17046, n4_adj_4375, n17045, n17044, n17043, n17042, 
        n28395, n1254, n42320, n7_adj_4376, n28584, n2964, n2963, 
        n2962, n2961, n2960, n2959, n2958, n2957, n2956, n2955, 
        n1283, n224, n42317, n14_adj_4377, n16_adj_4378, n4_adj_4379, 
        n28583, n28258, n28582, n3_adj_4380, n28394, n28257, n42312, 
        n8_adj_4381, n3_adj_4382, n28393, n28581, n28256, n28392, 
        n28580, n28255, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n5871, n33329, n33331, n42173, n17029, n28391, n28254, 
        n28390, n28389, n42331, n28579, n28388, n28387, n219, 
        n220, n223, n225, n17017, n33343, n28253, n28578, n28386, 
        n28577, n17012, n17011, n17010, n17009, n17008, n17007;
    wire [2:0]r_SM_Main_adj_5053;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_5054;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_5055;   // verilog/uart_tx.v(33[16:27])
    
    wire n28252, n41410, n313, n314, n5842, n17006, n17005, n17002, 
        n6_adj_4389, n28576, n28575, n16990, n33349, n28574, n316, 
        n318, n320;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n16986, n28385, n33351, n28573;
    wire [1:0]reg_B_adj_5064;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n16982, n16981, n16979, n33353, n1252, n5915, n5846, 
        n33355, n1258, n1253, n28251, n28384, n16971, n16970, 
        n16968, n16967, n16965, n958, n5937, n957, n5936, n5931, 
        n16964, n16963, n16962, n16961, n956, n5908, n33357, n33359, 
        n955, n5913, n5912, n5911, n5910, n33361, n954, n5914, 
        n1220, n28572, n33363, n33365, n1256, n953, n5916, n33367, 
        n21_adj_4392, n1224, n5917, n1225, n33369, n1255, n23_adj_4393, 
        n1223, n1325, n1324, n29111, n29110, n29109, n33371, n29108, 
        n29107, n29106, n29105, n1221, n1222, n29104, n1323, n29103, 
        n1322, n33373, n29102, n1219, n29101, n42336, n1321, n29100, 
        n1320, n1319, n1318, n4_adj_4394, n29099, n29098, n29097, 
        n29096, n29095, n29094, n29093, n29092, n29091, n29090, 
        n29089, n29088, n29087, n29086, n28571, n28570, n74, n29085, 
        n29084, n29083, n5928, n29082, n28569, n29081, n16918, 
        n42299, n16915, n29080, n29079, n28383, n29078, n29077, 
        n29076, n12_adj_4395, n13_adj_4396, n14_adj_4397, n15_adj_4398, 
        n16_adj_4399, n17_adj_4400, n18_adj_4401, n19_adj_4402, n20_adj_4403, 
        n21_adj_4404, n22_adj_4405, n23_adj_4406, n24_adj_4407, n25_adj_4408, 
        n29075, n42295, n41785, n783, n784, n785, n806, n807, 
        n884, n42287, n914, n915, n916, n917, n918, n35678, 
        n15576, n938, n939, n41780, n855, n852, n10283, n1043, 
        n1044, n1045, n1046, n1047, n1048, n1067, n1068, n41073, 
        n15567, n15570, n1169_adj_4409, n1170, n1171, n1172, n1173, 
        n1174, n1175, n1193, n1194, n5833, n5834, n5835, n1292, 
        n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1316, 
        n1317, n42319, n749, n748, n746, n42294, n1412, n1413, 
        n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1436, 
        n1437, n42258, n42256, n42255, n42252, n5850, n5851, n5852, 
        n5853, n5854, n5855, n5856, n5857, n5858, n5859, n1529, 
        n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
        n1538, n40507, n1553, n1554, n28568, n29074, n42248, n43025, 
        n43028, n43031, n43034, n43037, n3459, n3458, n3457, n3456, 
        n42247, n42210, n3452, n3453, n3454, n3455, n28382, n1643, 
        n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, 
        n1652, n1653, n29073, n1667, n1668, n29072, n29071, n6_adj_4410, 
        n41055, n5887, n5888, n5889, n29070, n1754, n1755, n1756, 
        n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
        n1765, n1778, n1779, n28567, n29069, n5893, n5894, n5895, 
        n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, 
        n5904, n5905, n29068, n1862, n1863, n1864, n1865, n1866, 
        n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, 
        n3362, n1886, n1887, n42234, n3358, n3357, n3356, n3355, 
        n3354, n3353, n3352, n3351, n3350, n18_adj_4411, n16_adj_4412, 
        n3342, n3344, n3346, n13_adj_4413, n1967, n1968, n1969, 
        n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
        n1978, n1979, n1980, n3340, n3339, n3338, n3337, n1991, 
        n1992, n3325, n3324, n3323, n3322, n3321, n5938, n5939, 
        n5940, n5959, n5979, n3313, n3314, n3315, n3316, n3317, 
        n3318, n3319, n3320, n2069, n2070, n2071, n2072, n2073, 
        n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, 
        n2082, n2083, n3312, n3311, n3310, n3309, n3308, n3307, 
        n3306, n3305, n3304, n2093, n2094, n3302, n3301, n3300, 
        n3299, n3298, n5943, n5944, n5945, n5946, n5947, n5948, 
        n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, 
        n5957, n5958, n29067, n2168, n2169, n2170, n2171, n2172, 
        n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, 
        n2181, n2182, n2183, n2192, n2193, n41043, n5962, n5963, 
        n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, 
        n5972, n5973, n5974, n5975, n5976, n5977, n5978, n39_adj_4414, 
        n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, 
        n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, 
        n2280, n3263, n37, n3258, n2288, n2289, n36, n34_adj_4415, 
        n28381, n3256, n3255, n3254, n3253, n3252, n3251, n33, 
        n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, 
        n28_adj_4416, n3246, n3247, n3248, n3249, n3250, n28566, 
        n29066, n28380, n28379, n2357, n2358, n2359, n2360, n2361, 
        n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
        n2370, n2371, n2372, n2373, n2374, n3245, n3244, n3243, 
        n3242, n3241, n3240, n2381, n2382, n22_adj_4417, n3238, 
        n3237, n3236, n3235, n3234, n6013, n6014, n6015, n6016, 
        n6017, n6018, n6019, n6020, n6021, n6022, n3230, n3231, 
        n3232, n3233, n28378, n2447, n2448, n2449, n2450, n2451, 
        n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, 
        n2460, n2461, n2462, n2463, n2464, n2465, n28377, n3225, 
        n2471, n2472, n3223, n3222, n3221, n3220, n6033, n6034, 
        n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, 
        n6043, n6044, n6045, n41566, n41792, n3217, n3218, n3219, 
        n29065, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
        n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
        n2549, n2550, n2551, n2552, n2553, n3216, n3215, n3214, 
        n3213, n2558, n2559, n29064, n3211, n3210, n3209, n6053, 
        n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
        n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, 
        n3207, n3208, n2618, n2619, n2620, n2621, n2622, n2623, 
        n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
        n2632, n2633, n2634, n2635, n2636, n2637, n2638, n3206, 
        n3205, n3204, n2642, n2643, n29063, n28243, n3202, n3201, 
        n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, 
        n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, 
        n6089, n6090, n6091, n6092, n6093, n6094, n3200, n2699, 
        n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, 
        n2708_adj_4418, n2709, n2710_adj_4419, n2711, n2712_adj_4420, 
        n2713, n2714_adj_4421, n2715, n2716_adj_4422, n2717, n2718_adj_4423, 
        n2719, n2720_adj_4424, n3199, n2723, n2724, n29062, n2777, 
        n2798, n2799, n2801, n2802, n29061, n29060, n35699, n29059, 
        n35580, n28565, n29058, n28564, n29057, n28563, n35597, 
        n28376, n28375, n29056, n3164, n29055, n28562, n3158, 
        n3157, n3156, n3155, n3154, n3153, n3152, n3151, n3150, 
        n3149, n3148, n3147, n3146, n3145, n3144, n3143, n3142, 
        n3141, n3140, n3139, n3138, n3137, n3136, n3135, n3134, 
        n3133, n3132, n3131, n29054, n40505, n46_adj_4425, n3125, 
        n3124, n3123, n3122, n3121, n3120, n3119, n3118, n3117, 
        n3116, n3115, n3114, n3113, n3112, n3111, n28242, n3110, 
        n3109, n3108, n3107, n3106, n28374, n17597, n17596, n29053, 
        n3105, n3104, n3103, n28373, n42188, n3102, n3101, n28241, 
        n3100, n28372, n28371, n17595, n28561, n17594, n17593, 
        n17592, n17591, n17590, n17589, n17588, n17587, n17586, 
        n17585, n17584, n17583, n17582, n17581, n17580, n17579, 
        n17578, n17577, n17576, n17575, n17574, n17573, n17572, 
        n17570, n17569, n17568, n17567, n17566, n33319, n17562, 
        n28240, n28239, n28560, n42184, n28559, n17561, n17560, 
        n33321, n33323, n17553, n17551, n17550, n17548, n17547, 
        n17546, n17545, n17544, n17543, n17542, n17541, n17540, 
        n17539, n17538, n17537, n17536, n17535, n17534, n17533, 
        n17532, n42182, n28558, n28557, n3065, n17531, n28556, 
        n29052, n17530, n28370, n17529, n3058, n17528, n17527, 
        n17526, n17524, n17523, n17522, n17521, n17520, n17519, 
        n17518, n17517, n17516, n17515, n17514, n17513, n17512, 
        n17511, n17510, n17509, n17508, n17507, n17506, n17505, 
        n17504, n17503, n17502, n17501, n17500, n17499, n17498, 
        n42180, n3057, n3056, n17497, n3055, n17496, n3054, n17495, 
        n3053, n17494, n3052, n17493, n3051, n17492, n3050, n17491, 
        n3049, n17490, n3048, n17489, n3047, n17488, n3046, n17487, 
        n3045, n17486, n3044, n17485, n3043, n17484, n3042, n17483, 
        n3041, n17482, n3040, n17481, n3039, n17480, n3038, n17479, 
        n3037, n3036, n3035, n3034, n3033, n3032, n1250, n3025, 
        n3024, n3023, n3022, n3021, n3020, n3019, n3018, n3017, 
        n3016, n3015, n3014, n3013, n3012, n3011, n3010, n3009, 
        n3008, n3007, n3006, n3005, n3004, n3003, n3002, n3001, 
        n16911, n15543, n1184, n42179, n29051, n28555, n28554, 
        n16905, n28369, n28368, n28553, n28552, n28551, n16899, 
        n16641, n28367, n28550, n2966, n28238, n16635, n28549, 
        n2958_adj_4426, n2957_adj_4427, n2956_adj_4428, n2955_adj_4429, 
        n2954_adj_4430, n2953_adj_4431, n2952_adj_4432, n2951_adj_4433, 
        n2950_adj_4434, n2949_adj_4435, n2948_adj_4436, n2947_adj_4437, 
        n2946_adj_4438, n2945_adj_4439, n2944_adj_4440, n2943_adj_4441, 
        n2942_adj_4442, n2941_adj_4443, n2940, n2939, n2938, n28548, 
        n28547, n28366, n2937, n2936, n2935, n2934, n2933, n29050, 
        n2925, n2924, n2923, n2922, n2921, n2920, n2919, n2918, 
        n2917, n2916, n2915, n2914_adj_4444, n2913_adj_4445, n2912_adj_4446, 
        n2911_adj_4447, n2910_adj_4448, n2909_adj_4449, n2908_adj_4450, 
        n28546, n16746, n16893, n28365, n28545, n29049, n29048, 
        n29047, n41862, n29046, n40487, n28544, n28543, n28542, 
        n41798, n16890, n40479, n42172, n16887, n16530, n28541, 
        n41570, n28540, n28364, n29045, n2907_adj_4451, n28539, 
        n29044, n28538, n28363, n29043, n29042, n29041, n29040, 
        n29039, n29038, n29037, n29036, n29035, n29034, n28362, 
        n41017, n29033, n28361, n29032, n42166, n33_adj_4452, n32, 
        n31_adj_4453, n30_adj_4454, n29_adj_4455, n28_adj_4456, n27_adj_4457, 
        n26, n25_adj_4458, n24_adj_4459, n23_adj_4460, n22_adj_4461, 
        n21_adj_4462, n20_adj_4463, n19_adj_4464, n18_adj_4465, n17_adj_4466, 
        n16_adj_4467, n15_adj_4468, n14_adj_4469, n2905_adj_4470, n2904_adj_4471, 
        n2903_adj_4472, n2902_adj_4473, n35585, n2867, n28537, n2858, 
        n2857, n2856, n2855_adj_4474, n2854, n2853, n2852, n2851, 
        n2850, n2849, n2848, n2847, n2846, n2845, n2844, n2843, 
        n2842, n2841, n2840, n2839, n2838, n2837, n2836, n2835, 
        n2834, n6_adj_4475, n29031, n4_adj_4476, n2825, n2824, n2823, 
        n2822, n2821, n42237, n42160, n2820, n2819, n35596, n2818, 
        n2817, n2816, n2815, n2814, n2813, n2812, n2811, n2810, 
        n2809, n42158, n2808, n2807, n2806, n2805, n2804, n2803, 
        n28360, n28359, n28536, n41598, n2768, n2758, n2757, n2756, 
        n2755, n2754, n2753, n2752, n2751, n2750, n2749, n2748, 
        n2747, n2746, n2745, n2744, n2743, n2742, n2741, n2740, 
        n2739, n2738, n2737, n2736, n2735, n7_adj_4477, n2725, 
        n2724_adj_4478, n2723_adj_4479, n2722, n29030, n2721, n29029, 
        n2719_adj_4480, n29028, n2717_adj_4481, n29027, n2715_adj_4482, 
        n29026, n2713_adj_4483, n29025, n2711_adj_4484, n29024, n2709_adj_4485, 
        n5832, n2707_adj_4486, n2706_adj_4487, n2705_adj_4488, n2704_adj_4489, 
        n2669, n29023, n29022, n28535, n2658, n2657, n2656, n2655, 
        n2654, n2653, n2652, n2651, n2650, n2649, n2648, n2647, 
        n2646, n2645, n2644, n2643_adj_4490, n2642_adj_4491, n2641, 
        n2640, n2639, n2638_adj_4492, n2637_adj_4493, n29021, n28534, 
        n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
        n1753, n1754_adj_4494, n1755_adj_4495, n1756_adj_4496, n1757_adj_4497, 
        n29020, n1758_adj_4498, n29019, n16_adj_4499, n29018, n1778_adj_4500, 
        n1813, n1814, n1815, n11_adj_4501, n1816, n1817, n1818, 
        n1819, n2636_adj_4502, n134, n135, n136, n137, n138, n139, 
        n140, n141, n142, n143, n144, n145, n146, n147, n148, 
        n149, n150, n151, n152, n153, n154, n155, n156, n157, 
        n158, n159, n160, n161, n162, n163, n164, n165, n10_adj_4503, 
        n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, 
        n1722, n1723, n1724, n1725, n29017, n29016, n29015, n28132, 
        n1679, n13_adj_4504, n12_adj_4505, n11_adj_4506, n10_adj_4507, 
        n9_adj_4508, n8_adj_4509, n7_adj_4510, n6_adj_4511, n5_adj_4512, 
        n4_adj_4513, n3_adj_4514, n24853, n28_adj_4515, n28533, n29014, 
        n29013, n2625_adj_4516, n2624_adj_4517, n2623_adj_4518, n2622_adj_4519, 
        n2621_adj_4520, n2620_adj_4521, n2619_adj_4522, n2618_adj_4523, 
        n2617, n2616, n26_adj_4524, n2615, n2614, n29012, n2613, 
        n2612, n2611, n2610, n2609, n2608, n2607, n2606, n2605, 
        n24867, n28131, n29011, n1580, n28130, n40999, n1646_adj_4525, 
        n1615, n1647_adj_4526, n1616, n1648_adj_4527, n1617, n1649_adj_4528, 
        n1618, n1650_adj_4529, n1619, n1651_adj_4530, n1620, n1652_adj_4531, 
        n1621, n1653_adj_4532, n1622, n1654, n1623, n1655, n1624, 
        n1656, n1625, n1657, n1658, n28532, n29010, n1547, n1548, 
        n1549, n1550, n1551, n1552, n1553_adj_4533, n1554_adj_4534, 
        n1555, n1556, n1557, n1558, n1516, n1517, n1518, n1519, 
        n1520, n1521, n1522, n1523, n1524, n1525, n28358, n1481, 
        n40456, n33333, n33335, n16832, n16831, n28531, n28530, 
        n16881, n28529, n28528, n42127, n24_adj_4535, n1448, n1449, 
        n1450, n1451, n1452, n1453, n1454, n1455, n29009, n1456, 
        n1457, n1458, n29008, n42123, n29007, n28527, n29006, 
        n1417_adj_4536, n1418_adj_4537, n1419_adj_4538, n1420_adj_4539, 
        n1421, n1422, n1423, n1424, n1425, n16872, n16869, n33375, 
        n33377, n33379, n33381, n33383, n33385, n33387, n29005, 
        n2570, n29004, n2558_adj_4540, n2557, n2556, n2555, n2554, 
        n2553_adj_4541, n2552_adj_4542, n2551_adj_4543, n2550_adj_4544, 
        n2549_adj_4545, n2548_adj_4546, n2547_adj_4547, n2546_adj_4548, 
        n2545_adj_4549, n2544_adj_4550, n2543_adj_4551, n2542_adj_4552, 
        n2541_adj_4553, n2540_adj_4554, n2539_adj_4555, n2538_adj_4556, 
        n2537_adj_4557, n28526, n29003, n42111, n42104, n2471_adj_4558, 
        n2_adj_4559, n29002, n29001, n2458_adj_4560, n2457_adj_4561, 
        n2456_adj_4562, n2455_adj_4563, n2454_adj_4564, n2453_adj_4565, 
        n2452_adj_4566, n29000, n2451_adj_4567, n2450_adj_4568, n2449_adj_4569, 
        n2448_adj_4570, n2447_adj_4571, n2446, n28999, n2445, n2444, 
        n2443, n2442, n2441, n42103, n2440, n2439, n2438, n2_adj_4572, 
        n3_adj_4573, n4_adj_4574, n5_adj_4575, n6_adj_4576, n7_adj_4577, 
        n8_adj_4578, n9_adj_4579, n10_adj_4580, n11_adj_4581, n12_adj_4582, 
        n13_adj_4583, n14_adj_4584, n15_adj_4585, n16_adj_4586, n17_adj_4587, 
        n18_adj_4588, n19_adj_4589, n20_adj_4590, n21_adj_4591, n22_adj_4592, 
        n23_adj_4593, n24_adj_4594, n25_adj_4595, n2_adj_4596, n3_adj_4597, 
        n4_adj_4598, n5_adj_4599, n6_adj_4600, n7_adj_4601, n8_adj_4602, 
        n9_adj_4603, n10_adj_4604, n11_adj_4605, n12_adj_4606, n13_adj_4607, 
        n14_adj_4608, n15_adj_4609, n16_adj_4610, n17_adj_4611, n18_adj_4612, 
        n19_adj_4613, n20_adj_4614, n21_adj_4615, n22_adj_4616, n23_adj_4617, 
        n24_adj_4618, n25_adj_4619, n28998, n28525, n28357, n2425, 
        n2424, n2423, n2422, n2421, n2420, n2419, n2418, n2417, 
        n2416, n2415, n2414, n2413, n2412, n2411, n2410, n2409, 
        n2408, n2407, n28997, n44, n41590, n28996, n2372_adj_4620, 
        n28995, n19_adj_4621, n28994, n28356, n2358_adj_4622, n2357_adj_4623, 
        n2356, n2355, n2354, n2353, n2352, n2351, n2350, n2349, 
        n2348, n2347, n2346, n2345, n2344, n2343, n2342, n2341, 
        n2340, n2339, n28993, n42_adj_4624, n2325, n2324, n2323, 
        n2322, n2321, n2320, n2319, n2318, n2317, n2316, n2315, 
        n2314, n2313, n2312, n2311, n2310, n2309, n2308, n16_adj_4625, 
        n28992, n28991, n40_adj_4626, n42_adj_4627, n44_adj_4628, 
        n45, n2273_adj_4629, n28355, n28129, n28990, n2258, n2257, 
        n2256, n2255, n2254, n2253, n2252, n2251, n2250, n2249, 
        n2248, n2247, n2246, n2245, n2244, n2243, n2242, n2241, 
        n2240, n28354, n2_adj_4630, n28989, n40415, n38_adj_4631, 
        n40_adj_4632, n42_adj_4633, n43_adj_4634, n42175, n28353, 
        n28352, n2225, n2224, n2223, n2222, n2221, n2220, n2219, 
        n2218, n2217, n2216, n2215, n2214, n2213, n2212, n2211, 
        n2210, n2209, n28988, n40413, n36_adj_4635, n38_adj_4636, 
        n40_adj_4637, n41, n2174_adj_4638, n28987, n28524, n28128, 
        n28229, n2158, n2157, n2156, n2155, n2154, n2153, n2152, 
        n2151, n2150, n2149, n2148, n2147, n2146, n2145, n2144, 
        n2143, n2142, n2141, n28351, n28986, n40411, n34_adj_4639, 
        n36_adj_4640, n38_adj_4641, n39_adj_4642, n41_adj_4643, n43_adj_4644, 
        n44_adj_4645, n45_adj_4646, n41600, n28985, n28350, n2125, 
        n2124, n2123, n2122, n2121, n2120, n2119, n2118, n2117, 
        n2116, n2115, n2114, n2113, n2112, n2111, n2110, n28984, 
        n32_adj_4647, n34_adj_4648, n37_adj_4649, n39_adj_4650, n41_adj_4651, 
        n42040, n43_adj_4652, n41602, n28983, n2075_adj_4653, n28982, 
        n28981, n28349, n28228, n2058, n2057, n28980, n30_adj_4654, 
        n31_adj_4655, n32_adj_4656, n33_adj_4657, n34_adj_4658, n35, 
        n37_adj_4659, n39_adj_4660, n41_adj_4661, n42_adj_4662, n43_adj_4663, 
        n45_adj_4664, n42068, n2056, n2055, n2054, n2053, n2052, 
        n2051, n2050, n2049, n2048, n2047, n2046, n2045, n2044, 
        n2043, n2042, n28979, n42245, n2025, n2024, n2023, n2022, 
        n2021, n28978, n40402, n28_adj_4665, n29_adj_4666, n30_adj_4667, 
        n31_adj_4668, n32_adj_4669, n33_adj_4670, n35_adj_4671, n37_adj_4672, 
        n42030, n39_adj_4673, n40_adj_4674, n41_adj_4675, n43_adj_4676, 
        n42169, n2020, n2019, n2018, n2017, n2016, n2015, n2014, 
        n2013, n2012, n2011, n28977, n28976, n28975, n40400, n26_adj_4677, 
        n27_adj_4678, n28_adj_4679, n29_adj_4680, n30_adj_4681, n31_adj_4682, 
        n33_adj_4683, n35_adj_4684, n42028, n37_adj_4685, n38_adj_4686, 
        n39_adj_4687, n41_adj_4688, n41856, n1976_adj_4689, n28974, 
        n28973, n28972, n28227, n28971, n1958, n1957, n28970, 
        n24_adj_4690, n25_adj_4691, n26_adj_4692, n27_adj_4693, n28_adj_4694, 
        n29_adj_4695, n30_adj_4696, n31_adj_4697, n32_adj_4698, n33_adj_4699, 
        n35_adj_4700, n36_adj_4701, n37_adj_4702, n39_adj_4703, n41858, 
        n1956, n1955, n1954, n1953, n1952, n1951, n1950, n1949, 
        n28523, n1948, n1947, n1946, n1945, n1944, n1943, n28969, 
        n28522, n28968, n28967, n28966, n40396, n22_adj_4704, n23_adj_4705, 
        n24_adj_4706, n25_adj_4707, n26_adj_4708, n27_adj_4709, n28_adj_4710, 
        n29_adj_4711, n30_adj_4712, n31_adj_4713, n33_adj_4714, n34_adj_4715, 
        n35_adj_4716, n37_adj_4717, n39_adj_4718, n41_adj_4719, n43_adj_4720, 
        n41866, n42076, n28965, n28964, n28963, n28962, n3330, 
        n28961, n20_adj_4721, n21_adj_4722, n22_adj_4723, n23_adj_4724, 
        n24_adj_4725, n25_adj_4726, n26_adj_4727, n27_adj_4728, n28_adj_4729, 
        n29_adj_4730, n31_adj_4731, n32_adj_4732, n33_adj_4733, n35_adj_4734, 
        n37_adj_4735, n42174, n39_adj_4736, n41_adj_4737, n3303, n28960, 
        n28959, n18_adj_4738, n19_adj_4739, n20_adj_4740, n21_adj_4741, 
        n22_adj_4742, n23_adj_4743, n24_adj_4744, n25_adj_4745, n26_adj_4746, 
        n27_adj_4747, n29_adj_4748, n30_adj_4749, n31_adj_4750, n33_adj_4751, 
        n35_adj_4752, n37_adj_4753, n39_adj_4754, n41_adj_4755, n43_adj_4756, 
        n45_adj_4757, n41868, n1877, n28958, n28957, n28521, n28348, 
        n28956, n42082, n28955, n28954, n16_adj_4758, n17_adj_4759, 
        n18_adj_4760, n19_adj_4761, n20_adj_4762, n21_adj_4763, n22_adj_4764, 
        n23_adj_4765, n25_adj_4766, n27_adj_4767, n28_adj_4768, n29_adj_4769, 
        n31_adj_4770, n33_adj_4771, n35_adj_4772, n41802, n37_adj_4773, 
        n39_adj_4774, n41_adj_4775, n43_adj_4776, n42296, n42080, 
        n28520, n28953, n3257, n1858, n1857, n1856, n1855, n1854, 
        n1853, n1852, n1851, n28952, n14_adj_4777, n16_adj_4778, 
        n17_adj_4779, n18_adj_4780, n19_adj_4781, n20_adj_4782, n21_adj_4783, 
        n22_adj_4784, n23_adj_4785, n25_adj_4786, n26_adj_4787, n27_adj_4788, 
        n29_adj_4789, n31_adj_4790, n33_adj_4791, n35_adj_4792, n37_adj_4793, 
        n42021, n39_adj_4794, n40_adj_4795, n41_adj_4796, n43_adj_4797, 
        n45_adj_4798, n42078, n1850, n1849, n1848, n1847, n1846, 
        n3239, n1845, n1844, n28951, n28950, n28949, n40386, n12_adj_4799, 
        n14_adj_4800, n15_adj_4801, n16_adj_4802, n17_adj_4803, n18_adj_4804, 
        n19_adj_4805, n20_adj_4806, n21_adj_4807, n23_adj_4808, n24_adj_4809, 
        n25_adj_4810, n27_adj_4811, n29_adj_4812, n31_adj_4813, n42239, 
        n33_adj_4814, n35_adj_4815, n42017, n37_adj_4816, n38_adj_4817, 
        n39_adj_4818, n41_adj_4819, n43_adj_4820, n42015, n3224, n28948, 
        n10_adj_4821, n12_adj_4822, n13_adj_4823, n14_adj_4824, n15_adj_4825, 
        n16_adj_4826, n17_adj_4827, n18_adj_4828, n19_adj_4829, n21_adj_4830, 
        n22_adj_4831, n23_adj_4832, n25_adj_4833, n27_adj_4834, n29_adj_4835, 
        n42241, n31_adj_4836, n33_adj_4837, n42011, n35_adj_4838, 
        n36_adj_4839, n37_adj_4840, n39_adj_4841, n41_adj_4842, n42183, 
        n42243, n3212, n1825, n1824, n28947, n8_adj_4843, n10_adj_4844, 
        n11_adj_4845, n12_adj_4846, n13_adj_4847, n14_adj_4848, n15_adj_4849, 
        n16_adj_4850, n17_adj_4851, n19_adj_4852, n20_adj_4853, n21_adj_4854, 
        n23_adj_4855, n25_adj_4856, n42005, n27_adj_4857, n29_adj_4858, 
        n31_adj_4859, n42003, n33_adj_4860, n34_adj_4861, n35_adj_4862, 
        n37_adj_4863, n39_adj_4864, n41891, n41_adj_4865, n43_adj_4866, 
        n44_adj_4867, n45_adj_4868, n41893, n41895, n1823, n1822, 
        n3203, n1821, n6_adj_4869, n8_adj_4870, n9_adj_4871, n10_adj_4872, 
        n11_adj_4873, n12_adj_4874, n13_adj_4875, n14_adj_4876, n15_adj_4877, 
        n17_adj_4878, n19_adj_4879, n21_adj_4880, n23_adj_4881, n41794, 
        n25_adj_4882, n27_adj_4883, n29_adj_4884, n31_adj_4885, n32_adj_4886, 
        n33_adj_4887, n35_adj_4888, n37_adj_4889, n41793, n1820, n28946, 
        n4_adj_4890, n6_adj_4891, n7_adj_4892, n8_adj_4893, n9_adj_4894, 
        n10_adj_4895, n11_adj_4896, n12_adj_4897, n13_adj_4898, n15_adj_4899, 
        n16_adj_4900, n17_adj_4901, n19_adj_4902, n21_adj_4903, n41787, 
        n23_adj_4904, n24_adj_4905, n25_adj_4906, n27_adj_4907, n29_adj_4908, 
        n30_adj_4909, n31_adj_4910, n33_adj_4911, n43083, n35_adj_4912, 
        n37_adj_4913, n42298, n39_adj_4914, n41_adj_4915, n43_adj_4916, 
        n45_adj_4917, n42212, n28945, n28519, n28226, n5818, n5819, 
        n5820, n5821, n5822, n5823, n5824, n5808, n5809, n5810, 
        n5811, n5812, n5813, n5814, n28944, n28943, n28518, n28942, 
        n28941, n5801, n5802, n5803, n5804, n5805, n35530, n15459, 
        n28940, n28939, n42161, n28517, n28347, n28516, n28346, 
        n28938, n28937, n40961, n29951, n29950, n43021, n13_adj_4918, 
        n11_adj_4919, n28936, n28935, n29949, n28515, n28514, n28225, 
        n28934, n35524, n28933, n28932, n28513, n42069, n29948, 
        n29947, n28512, n28931, n28930, n28511, n28510, n28509, 
        n28929, n28345, n28928, n28927, n28926, n29946, n29945, 
        n28925, n28924, n28127, n28344, n28343, n28224, n28923, 
        n42334, n28126, n28922, n28921, n29944, n28920, n28223, 
        n28222, n28919, n28918, n29943, n28917, n28221, n28916, 
        n42066, n28915, n29942, n28914, n28220, n28125, n28124, 
        n35602, n28913, n28912, n29941, n28911, n28342, n28910, 
        n28909, n42061, n29940, n28908, n28123, n28219, n28508, 
        n28907, n29939, n28906, n28507, n28506, n28341, n28905, 
        n28904, n42060, n29938, n28903, n28340, n28218, n42057, 
        n28902, n28901, n28900, n42056, n42171, n29937, n40361, 
        n40359, n28339, n28122, n28899, n28898, n33347, n33341, 
        n28897, n40346, n40339, n19_adj_4920, n28896, n42049, n40332, 
        n11_adj_4921, n35361, n33317, n29936, n40915, n40908, n42047, 
        n28895, n42012, n40_adj_4922, n8_adj_4923, n28894, n43272, 
        n41580, n42043, n42041, n40897, n28893, n40893, n12_adj_4924, 
        n40891, n5_adj_4925, n42039, n42038, n28892, n40882, n28217, 
        n42035, n28891, n42034, n41584, n28890, n42_adj_4926, n41_adj_4927, 
        n40_adj_4928, n39_adj_4929, n37_adj_4930, n36_adj_4931, n28338, 
        n28889, n30_adj_4932, n42031, n28888, n28887, n28886, n42025, 
        n42022, n22_adj_4933, n19_adj_4934, n18_adj_4935, n15_adj_4936, 
        n28337, n42018, n28885, n39_adj_4937, n38_adj_4938, n37_adj_4939, 
        n35_adj_4940, n34_adj_4941, n28884, n41586, n28883, n28882, 
        n27_adj_4942, n28881, n28880, n24907, n8849, n29935, n29934, 
        n29933, n29932, n29931, n29930, n29929, n29928, n29927, 
        n28879, n29926, n28878, n28877, n40322, n28876, n28875, 
        n29925, n29924, n41999, n29923, n29922, n41897, n41888, 
        n41886, n29921, n40861, n40859, n28874, n10087, n40857, 
        n40854, n10086, n10085, n10084, n10083, n10082, n41882, 
        n40849, n40845, n42004, n28336, n41876, n41853, n42235, 
        n41872, n40318, n42181, n28873, n41869, n40316, n28872, 
        n41847, n41845, n41841, n42042, n28871, n28870, n35686, 
        n28869, n28121, n41810, n35564, n28868, n40807, n41634, 
        n40801, n41640, n40799, n42008, n34657, n42006, n44_adj_4943, 
        n43_adj_4944, n42_adj_4945, n41_adj_4946, n40793, n40_adj_4947, 
        n38_adj_4948, n40789, n41508, n41292, n30_adj_4949, n26_adj_4950, 
        n10_adj_4951, n42333, n41290, n40777, n41266, n41336, n28867, 
        n42240, n13195, n28505, n28120, n28866, n40763, n28865, 
        n28864, n28863, n28504, n28862, n28503, n40755, n3_adj_4952, 
        n28861, n40751, n40747, n28860, n40739, n28859, n28858, 
        n41935, n28119, n28857, n40737, n28856, n28855, n28854, 
        n42238, n28853, n28852, n28851, n40729, n28850, n36606, 
        n28849, n28848, n28847, n28118, n28846, n28845, n28502, 
        n40709, n28844, n28843, n40703, n28842, n28841, n28840, 
        n41996, n40701, n40699, n42225, n40693, n40691, n5800, 
        n5817, n40687, n41398, n28839, n28838, n5838, n5877, n37954, 
        n26_adj_4953, n5925, n37950, n24_adj_4954, n6072, n37_adj_4955, 
        n22_adj_4956, n35_adj_4957, n34_adj_4958, n32_adj_4959, n31_adj_4960, 
        n18_adj_4961, n25_adj_4962, n40299, n40297, n40293, n40285, 
        n28837, n40279, n40277, n40275, n40273, n40261, n40259, 
        n40255, n35648, n41945, n42218, n40203, n40201, n41696, 
        n40199, n40198, n40197, n28335, n40196, n28836, n16695, 
        n28334, n28835, n28834, n40195, n28117, n40194, n40193, 
        n42224, n40192, n28833, n28832, n28831, n40191, n28830, 
        n28116, n28829, n28828, n40190, n40189, n40188, n13_adj_4963, 
        n40187, n11_adj_4964, n40186, n2_adj_4965, n3_adj_4966, n4_adj_4967, 
        n5_adj_4968, n6_adj_4969, n7_adj_4970, n8_adj_4971, n9_adj_4972, 
        n10_adj_4973, n11_adj_4974, n12_adj_4975, n13_adj_4976, n14_adj_4977, 
        n15_adj_4978, n16_adj_4979, n17_adj_4980, n18_adj_4981, n19_adj_4982, 
        n20_adj_4983, n21_adj_4984, n22_adj_4985, n23_adj_4986, n24_adj_4987, 
        n25_adj_4988, n26_adj_4989, n27_adj_4990, n28_adj_4991, n29_adj_4992, 
        n30_adj_4993, n31_adj_4994, n32_adj_4995, n33_adj_4996, n28827, 
        n28826, n28825, n41989, n28115, n28824, n28823, n28333, 
        n28822, n28821, n28820, n28332, n42222, n40185, n40184, 
        n28819, n28501, n28818, n40183, n28817, n28816, n28500, 
        n28815, n28814, n35534, n40182, n28813, n28499, n40181, 
        n28812, n28811, n28810, n28498, n40180, n28809, n28808, 
        n28807, n28331, n28806, n28330, n35660, n28216, n28805, 
        n28114, n40179, n40178, n28804, n28803, n28802, n28801, 
        n40177, n28800, n28497, n28799, n28329, n28798, n28797, 
        n28796, n28795, n28794, n28793, n28113, n40176, n28215, 
        n28328, n28792, n28112, n28327, n28791, n28790, n28789, 
        n35632, n28788, n28787, n28786, n28326, n28785, n28784, 
        n28783, n28782, n40175, n28781, n28325, n28780, n28214, 
        n28779, n28324, n40174, n40173, n28778, n28777, n28776, 
        n40172, n40171, n40170, n28496, n40169, n40168, n28775, 
        n28774, n28773, n28772, n28771, n28770, n28769, n28768, 
        n28767, n28213, n28766, n28765, n28764, n28495, n28763, 
        n28762, n28761, n28760, n28759, n28323, n28494, n28493, 
        n41953, n28758, n28757, n28756, n28755, n28754, n28753, 
        n28322, n28752, n28751, n28750, n28749, n28748, n28747, 
        n28212, n28746, n28745, n28744, n28743, n41961, n42232, 
        n28111, n28211, n28210, n40245, n35694, n28321, n41803, 
        n28209, n28719, n28718, n28717, n28716, n28715, n28714, 
        n28713, n28712, n28711, n28208, n28710, n28492, n28207, 
        n28709, n28708, n28320, n28707, n28706, n28705, n28704, 
        n28206, n28703, n28319, n28702, n28701, n28700, n28699, 
        n28318, n28205, n35642, n28698, n28697, n28204, n28491, 
        n35572, n28696, n28695, n28694, n28693, n28692, n28490, 
        n28489, n28203, n28317, n35481, n28488, n15464, n37700, 
        n37696, n28316, n28487, n37690, n28315, n40239, n28202, 
        n28314, n28313, n37686, n28486, n43071, n37658, n37656, 
        n37650, n37648, n34_adj_4997, n33_adj_4998, n32_adj_4999, 
        n31_adj_5000, n30_adj_5001, n41342, n35317, n35307, n40121, 
        n37588, n8_adj_5002, n7_adj_5003, n42228, n42337, n42233, 
        n42338, n37586, n37584, n37578, n37576, n47_adj_5004, n46_adj_5005, 
        n4_adj_5006, n37558, n36_adj_5007, n37554, n37550, n28_adj_5008, 
        n36885, n3_adj_5009, n43089, n43079, n37092, n37992, n37462, 
        n37460, n41963, n42229, n28_adj_5010, n27_adj_5011, n26_adj_5012, 
        n25_adj_5013, n40227, n36839, n36917, n37155, n41516;
    
    VCC i2 (.Y(VCC_net));
    SB_IO ID1_input (.PACKAGE_PIN(PIN_10), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID1_input.PIN_TYPE = 6'b000001;
    defparam ID1_input.PULLUP = 1'b1;
    defparam ID1_input.NEG_TRIGGER = 1'b0;
    defparam ID1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO ID2_input (.PACKAGE_PIN(PIN_11), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID2_input.PIN_TYPE = 6'b000001;
    defparam ID2_input.PULLUP = 1'b1;
    defparam ID2_input.NEG_TRIGGER = 1'b0;
    defparam ID2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY rem_4_add_1251_8 (.CI(n29052), .I0(n1853), .I1(n1877), .CO(n29053));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[0]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 div_46_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4643));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_DFF h2_56 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_80[0]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_57 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF dir_61 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 rem_4_add_1251_7_lut (.I0(n1854), .I1(n1854), .I2(n43071), 
            .I3(n29051), .O(n1953)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_7_lut.LUT_INIT = 16'hA3AC;
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_6_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b000001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.VCC_net(VCC_net), .timer({timer}), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .bit_ctr({bit_ctr}), .n40170(n40170), 
            .GND_net(GND_net), .n11(n11_adj_4921), .n33373(n33373), .n33375(n33375), 
            .n33361(n33361), .n33363(n33363), .n33365(n33365), .n33367(n33367), 
            .n33369(n33369), .n33335(n33335), .n33377(n33377), .n33379(n33379), 
            .n33381(n33381), .n33383(n33383), .n33385(n33385), .n33323(n33323), 
            .n33371(n33371), .n33353(n33353), .n33355(n33355), .n33357(n33357), 
            .n33359(n33359), .n33341(n33341), .n33343(n33343), .n33347(n33347), 
            .n33349(n33349), .n33351(n33351), .n33331(n33331), .n33333(n33333), 
            .n33329(n33329), .n33327(n33327), .n33317(n33317), .n33319(n33319), 
            .n33321(n33321), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n40197(n40197), .n19(n19_adj_4920), .n40169(n40169), .n40168(n40168), 
            .n40196(n40196), .n40181(n40181), .n40180(n40180), .n40195(n40195), 
            .n40179(n40179), .\state_3__N_362[1] (state_3__N_362[1]), .\state[1] (state[1]), 
            .n1163(n1163), .\state[0] (state[0]), .n4385(n4385), .n40176(n40176), 
            .\one_wire_N_513[10] (one_wire_N_513[10]), .\one_wire_N_513[8] (one_wire_N_513[8]), 
            .\one_wire_N_513[5] (one_wire_N_513[5]), .\one_wire_N_513[11] (one_wire_N_513[11]), 
            .\one_wire_N_513[7] (one_wire_N_513[7]), .\one_wire_N_513[9] (one_wire_N_513[9]), 
            .\one_wire_N_513[6] (one_wire_N_513[6]), .start(start), .n15464(n15464), 
            .n35361(n35361), .n24867(n24867), .n33325(n33325), .n17072(n17072), 
            .n17071(n17071), .n17070(n17070), .n17069(n17069), .n17068(n17068), 
            .n17067(n17067), .n17066(n17066), .n17065(n17065), .n17064(n17064), 
            .n17063(n17063), .n17062(n17062), .n17061(n17061), .n17060(n17060), 
            .n17059(n17059), .n17058(n17058), .n17057(n17057), .n17056(n17056), 
            .n17055(n17055), .n35481(n35481), .n40194(n40194), .n17054(n17054), 
            .n17053(n17053), .n24907(n24907), .n17052(n17052), .n17051(n17051), 
            .n17050(n17050), .n17049(n17049), .n17048(n17048), .n17047(n17047), 
            .n17046(n17046), .n37092(n37092), .n17045(n17045), .n17044(n17044), 
            .n17043(n17043), .n17042(n17042), .n40175(n40175), .n16530(n16530), 
            .n16754(n16754), .PIN_8_c(PIN_8_c), .n36917(n36917), .n40172(n40172), 
            .n40192(n40192), .n40191(n40191), .n40190(n40190), .n40189(n40189), 
            .n40188(n40188), .n40187(n40187), .n40186(n40186), .n40193(n40193), 
            .n40185(n40185), .n40171(n40171), .n40184(n40184), .n40199(n40199), 
            .n33387(n33387), .n16831(n16831), .n17017(n17017), .n40183(n40183), 
            .n40177(n40177), .n40198(n40198), .n40182(n40182), .n40178(n40178), 
            .n40174(n40174), .n40173(n40173), .n24853(n24853), .\color[2] (color[2]), 
            .\color[3] (color[3]), .\color[4] (color[4]), .\color[1] (color[1])) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(98[10] 104[2])
    SB_IO ID0_input (.PACKAGE_PIN(PIN_9), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID0_input.PIN_TYPE = 6'b000001;
    defparam ID0_input.PULLUP = 1'b1;
    defparam ID0_input.NEG_TRIGGER = 1'b0;
    defparam ID0_input.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY rem_4_add_1251_7 (.CI(n29051), .I0(n1854), .I1(n43071), .CO(n29052));
    SB_CARRY rem_4_add_1921_3 (.CI(n28796), .I0(n2858), .I1(GND_net), 
            .CO(n28797));
    SB_LUT4 rem_4_add_1251_6_lut (.I0(n1855), .I1(n1855), .I2(n43071), 
            .I3(n29050), .O(n1954)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1921_2 (.CI(VCC_net), .I0(n2958_adj_4426), .I1(VCC_net), 
            .CO(n28796));
    SB_LUT4 rem_4_add_1988_28_lut (.I0(n2966), .I1(n2933), .I2(VCC_net), 
            .I3(n28795), .O(n3032)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1251_6 (.CI(n29050), .I0(n1855), .I1(n43071), .CO(n29051));
    SB_LUT4 div_46_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n655));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1251_5_lut (.I0(n1856), .I1(n1856), .I2(n1877), 
            .I3(n29049), .O(n1955)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1251_5 (.CI(n29049), .I0(n1856), .I1(n1877), .CO(n29050));
    SB_LUT4 rem_4_add_1251_4_lut (.I0(n1857), .I1(n1857), .I2(n1877), 
            .I3(n29048), .O(n1956)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1988_27_lut (.I0(GND_net), .I1(n2934), .I2(VCC_net), 
            .I3(n28794), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_4 (.CI(n29048), .I0(n1857), .I1(n1877), .CO(n29049));
    SB_LUT4 rem_4_add_1251_3_lut (.I0(n1858), .I1(n1858), .I2(n43071), 
            .I3(n29047), .O(n1957)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1988_27 (.CI(n28794), .I0(n2934), .I1(VCC_net), 
            .CO(n28795));
    SB_CARRY rem_4_add_1251_3 (.CI(n29047), .I0(n1858), .I1(n43071), .CO(n29048));
    SB_LUT4 div_46_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1988_26_lut (.I0(GND_net), .I1(n2935), .I2(VCC_net), 
            .I3(n28793), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_2 (.CI(VCC_net), .I0(n1958), .I1(VCC_net), 
            .CO(n29047));
    SB_CARRY rem_4_add_1988_26 (.CI(n28793), .I0(n2935), .I1(VCC_net), 
            .CO(n28794));
    SB_LUT4 rem_4_add_1318_18_lut (.I0(n1976_adj_4689), .I1(n1943), .I2(VCC_net), 
            .I3(n29046), .O(n2042)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1988_25_lut (.I0(GND_net), .I1(n2936), .I2(VCC_net), 
            .I3(n28792), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_17_lut (.I0(GND_net), .I1(n1944), .I2(VCC_net), 
            .I3(n29045), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_25 (.CI(n28792), .I0(n2936), .I1(VCC_net), 
            .CO(n28793));
    SB_CARRY rem_4_add_1988_2 (.CI(VCC_net), .I0(n3058), .I1(VCC_net), 
            .CO(n28770));
    SB_CARRY rem_4_add_1318_17 (.CI(n29045), .I0(n1944), .I1(VCC_net), 
            .CO(n29046));
    SB_LUT4 rem_4_add_1988_24_lut (.I0(GND_net), .I1(n2937), .I2(VCC_net), 
            .I3(n28791), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_16_lut (.I0(GND_net), .I1(n1945), .I2(VCC_net), 
            .I3(n29044), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_16 (.CI(n29044), .I0(n1945), .I1(VCC_net), 
            .CO(n29045));
    SB_LUT4 rem_4_add_1318_15_lut (.I0(GND_net), .I1(n1946), .I2(VCC_net), 
            .I3(n29043), .O(n2013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_24 (.CI(n28791), .I0(n2937), .I1(VCC_net), 
            .CO(n28792));
    SB_LUT4 rem_4_add_1988_23_lut (.I0(GND_net), .I1(n2938), .I2(VCC_net), 
            .I3(n28790), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_15 (.CI(n29043), .I0(n1946), .I1(VCC_net), 
            .CO(n29044));
    SB_CARRY rem_4_add_1988_23 (.CI(n28790), .I0(n2938), .I1(VCC_net), 
            .CO(n28791));
    SB_LUT4 rem_4_add_2055_29_lut (.I0(n3065), .I1(n3032), .I2(VCC_net), 
            .I3(n28769), .O(n3131)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_2055_28_lut (.I0(GND_net), .I1(n3033), .I2(VCC_net), 
            .I3(n28768), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_14_lut (.I0(GND_net), .I1(n1947), .I2(VCC_net), 
            .I3(n29042), .O(n2014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_22_lut (.I0(GND_net), .I1(n2939), .I2(VCC_net), 
            .I3(n28789), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_14 (.CI(n29042), .I0(n1947), .I1(VCC_net), 
            .CO(n29043));
    SB_CARRY rem_4_add_1988_22 (.CI(n28789), .I0(n2939), .I1(VCC_net), 
            .CO(n28790));
    SB_LUT4 rem_4_add_1318_13_lut (.I0(GND_net), .I1(n1948), .I2(VCC_net), 
            .I3(n29041), .O(n2015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_21_lut (.I0(GND_net), .I1(n2940), .I2(VCC_net), 
            .I3(n28788), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_28 (.CI(n28768), .I0(n3033), .I1(VCC_net), 
            .CO(n28769));
    SB_LUT4 rem_4_add_2055_27_lut (.I0(GND_net), .I1(n3034), .I2(VCC_net), 
            .I3(n28767), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_27 (.CI(n28767), .I0(n3034), .I1(VCC_net), 
            .CO(n28768));
    SB_LUT4 rem_4_add_715_8_lut (.I0(n1085), .I1(n1052), .I2(VCC_net), 
            .I3(n28243), .O(n1151)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_825_i34_4_lut (.I0(n655), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34_adj_4639));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY rem_4_add_1318_13 (.CI(n29041), .I0(n1948), .I1(VCC_net), 
            .CO(n29042));
    SB_CARRY rem_4_add_1988_21 (.CI(n28788), .I0(n2940), .I1(VCC_net), 
            .CO(n28789));
    SB_LUT4 rem_4_add_1318_12_lut (.I0(GND_net), .I1(n1949), .I2(VCC_net), 
            .I3(n29040), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_20_lut (.I0(GND_net), .I1(n2941_adj_4443), .I2(VCC_net), 
            .I3(n28787), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_20 (.CI(n28787), .I0(n2941_adj_4443), .I1(VCC_net), 
            .CO(n28788));
    SB_CARRY rem_4_add_1318_12 (.CI(n29040), .I0(n1949), .I1(VCC_net), 
            .CO(n29041));
    SB_LUT4 rem_4_add_1318_11_lut (.I0(GND_net), .I1(n1950), .I2(VCC_net), 
            .I3(n29039), .O(n2017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_19_lut (.I0(GND_net), .I1(n2942_adj_4442), .I2(VCC_net), 
            .I3(n28786), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_11 (.CI(n29039), .I0(n1950), .I1(VCC_net), 
            .CO(n29040));
    SB_LUT4 i35278_3_lut (.I0(n34_adj_4639), .I1(n95), .I2(n41_adj_4643), 
            .I3(GND_net), .O(n42042));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35278_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35279_3_lut (.I0(n42042), .I1(n94), .I2(n43_adj_4644), .I3(GND_net), 
            .O(n42043));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35279_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34291_4_lut (.I0(n43_adj_4644), .I1(n41_adj_4643), .I2(n39_adj_4642), 
            .I3(n40359), .O(n41055));
    defparam i34291_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i12613_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n13195), .I3(GND_net), .O(n17295));   // verilog/coms.v(126[12] 289[6])
    defparam i12613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_825_i38_3_lut (.I0(n36_adj_4640), .I1(n96), 
            .I2(n39_adj_4642), .I3(GND_net), .O(n38_adj_4641));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35075_3_lut (.I0(n42043), .I1(n93), .I2(n45_adj_4646), .I3(GND_net), 
            .O(n44_adj_4645));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35075_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_2055_26_lut (.I0(GND_net), .I1(n3035), .I2(VCC_net), 
            .I3(n28766), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_10_lut (.I0(GND_net), .I1(n1951), .I2(VCC_net), 
            .I3(n29038), .O(n2018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34834_4_lut (.I0(n44_adj_4645), .I1(n38_adj_4641), .I2(n45_adj_4646), 
            .I3(n41055), .O(n41598));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34834_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut (.I0(n41598), .I1(n15561), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_CARRY rem_4_add_1988_19 (.CI(n28786), .I0(n2942_adj_4442), .I1(VCC_net), 
            .CO(n28787));
    SB_CARRY rem_4_add_2055_26 (.CI(n28766), .I0(n3035), .I1(VCC_net), 
            .CO(n28767));
    SB_LUT4 div_46_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_715_7_lut (.I0(GND_net), .I1(n1053), .I2(VCC_net), 
            .I3(n28242), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4359), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n654));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i744_1_lut.LUT_INIT = 16'h5555;
    SB_DFF color__i4 (.Q(color[4]), .C(LED_c), .D(n17562));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_DFF color__i2 (.Q(color[2]), .C(LED_c), .D(n17560));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_DFF color__i3 (.Q(color[3]), .C(LED_c), .D(n17561));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_DFF color__i1 (.Q(color[1]), .C(LED_c), .D(n17553));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_LUT4 div_46_LessThan_742_i36_4_lut (.I0(n654), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36_adj_4635));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY rem_4_add_715_7 (.CI(n28242), .I0(n1053), .I1(VCC_net), .CO(n28243));
    SB_LUT4 rem_4_add_715_6_lut (.I0(GND_net), .I1(n1054), .I2(GND_net), 
            .I3(n28241), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_6 (.CI(n28241), .I0(n1054), .I1(GND_net), .CO(n28242));
    SB_LUT4 rem_4_add_715_5_lut (.I0(GND_net), .I1(n1055), .I2(GND_net), 
            .I3(n28240), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_5 (.CI(n28240), .I0(n1055), .I1(GND_net), .CO(n28241));
    SB_LUT4 rem_4_add_715_4_lut (.I0(GND_net), .I1(n1056), .I2(VCC_net), 
            .I3(n28239), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_742_i40_3_lut (.I0(n38_adj_4636), .I1(n96), 
            .I2(n41), .I3(GND_net), .O(n40_adj_4637));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35469_4_lut (.I0(n40_adj_4637), .I1(n36_adj_4635), .I2(n41), 
            .I3(n40386), .O(n42233));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35469_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35470_3_lut (.I0(n42233), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n42234));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35470_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY rem_4_add_715_4 (.CI(n28239), .I0(n1056), .I1(VCC_net), .CO(n28240));
    SB_LUT4 i35402_3_lut (.I0(n42234), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n42166));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35402_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_2055_25_lut (.I0(GND_net), .I1(n3036), .I2(VCC_net), 
            .I3(n28765), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1589 (.I0(n42166), .I1(n15504), .I2(n93), .I3(n1169_adj_4409), 
            .O(n1193));
    defparam i1_4_lut_adj_1589.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4634));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2055_25 (.CI(n28765), .I0(n3036), .I1(VCC_net), 
            .CO(n28766));
    SB_LUT4 rem_4_add_2055_24_lut (.I0(GND_net), .I1(n3037), .I2(VCC_net), 
            .I3(n28764), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4381), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n653));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_18_lut (.I0(GND_net), .I1(n2943_adj_4441), .I2(VCC_net), 
            .I3(n28785), .O(n3010)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i659_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1318_10 (.CI(n29038), .I0(n1951), .I1(VCC_net), 
            .CO(n29039));
    SB_LUT4 div_46_LessThan_657_i38_4_lut (.I0(n653), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38_adj_4631));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_657_i42_3_lut (.I0(n40_adj_4632), .I1(n96), 
            .I2(n43_adj_4634), .I3(GND_net), .O(n42_adj_4633));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35296_4_lut (.I0(n42_adj_4633), .I1(n38_adj_4631), .I2(n43_adj_4634), 
            .I3(n40402), .O(n42060));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35296_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_add_1318_9_lut (.I0(GND_net), .I1(n1952), .I2(VCC_net), 
            .I3(n29037), .O(n2019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35297_3_lut (.I0(n42060), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n42061));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35297_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY rem_4_add_1988_18 (.CI(n28785), .I0(n2943_adj_4441), .I1(VCC_net), 
            .CO(n28786));
    SB_LUT4 i1_4_lut_adj_1590 (.I0(n42061), .I1(n15558), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1590.LUT_INIT = 16'hceef;
    SB_LUT4 mux_71_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[4]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_106[4]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_24 (.CI(n28764), .I0(n3037), .I1(VCC_net), 
            .CO(n28765));
    SB_LUT4 rem_4_add_2055_23_lut (.I0(GND_net), .I1(n3038), .I2(VCC_net), 
            .I3(n28763), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_71_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[5]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_106[5]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_17_lut (.I0(GND_net), .I1(n2944_adj_4440), .I2(VCC_net), 
            .I3(n28784), .O(n3011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_17 (.CI(n28784), .I0(n2944_adj_4440), .I1(VCC_net), 
            .CO(n28785));
    SB_LUT4 i22897_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4323), .I3(GND_net), 
            .O(n8));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22897_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i22889_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4325), .I3(GND_net), 
            .O(n6_adj_4323));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22889_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 rem_4_add_715_3_lut (.I0(GND_net), .I1(n1057), .I2(VCC_net), 
            .I3(n28238), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4376), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22873_2_lut (.I0(n651), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4342));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22873_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_570_i40_4_lut (.I0(n652), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40_adj_4626));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_570_i44_3_lut (.I0(n42_adj_4627), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4628));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34826_4_lut (.I0(n44_adj_4628), .I1(n40_adj_4626), .I2(n45), 
            .I3(n40415), .O(n41590));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34826_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1591 (.I0(n41590), .I1(n15501), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1591.LUT_INIT = 16'hceef;
    SB_LUT4 i22857_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_4476), .I3(GND_net), 
            .O(n6_adj_4475));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22857_3_lut.LUT_INIT = 16'he8e8;
    SB_CARRY rem_4_add_2055_23 (.CI(n28763), .I0(n3038), .I1(VCC_net), 
            .CO(n28764));
    SB_LUT4 i22841_2_lut (.I0(n650), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4559));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22841_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4367), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n651));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_481_i42_4_lut (.I0(n651), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42_adj_4624));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35292_3_lut (.I0(n42_adj_4624), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n42056));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35292_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35293_3_lut (.I0(n42056), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n42057));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35293_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1592 (.I0(n42057), .I1(n15498), .I2(n96), .I3(n35317), 
            .O(n806));
    defparam i1_4_lut_adj_1592.LUT_INIT = 16'hefce;
    SB_LUT4 i22817_2_lut (.I0(n511), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22817_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4343), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n650));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_390_i44_4_lut (.I0(n650), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i34822_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n41586));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34822_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_2055_22_lut (.I0(GND_net), .I1(n3039), .I2(VCC_net), 
            .I3(n28762), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1593 (.I0(n41586), .I1(n15494), .I2(n97), .I3(n35315), 
            .O(n671));
    defparam i1_4_lut_adj_1593.LUT_INIT = 16'hefce;
    SB_LUT4 i22972_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4630));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22972_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4356), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i299_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1318_9 (.CI(n29037), .I0(n1952), .I1(VCC_net), 
            .CO(n29038));
    SB_LUT4 div_46_LessThan_297_i46_4_lut (.I0(n511), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46_adj_4425));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1594 (.I0(n46_adj_4425), .I1(n15555), .I2(n98), 
            .I3(n35307), .O(n533));
    defparam i1_4_lut_adj_1594.LUT_INIT = 16'hefce;
    SB_LUT4 i1_4_lut_adj_1595 (.I0(n224), .I1(n99), .I2(n15491), .I3(n558), 
            .O(n5_adj_4925));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i1_4_lut_adj_1595.LUT_INIT = 16'h555d;
    SB_LUT4 div_46_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4382), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33688_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n40121));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33688_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1596 (.I0(n40121), .I1(n15491), .I2(n99), .I3(n5_adj_4925), 
            .O(n392));
    defparam i1_4_lut_adj_1596.LUT_INIT = 16'hefce;
    SB_LUT4 div_46_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n15549));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1597 (.I0(n81), .I1(n15543), .I2(GND_net), .I3(GND_net), 
            .O(n15535));
    defparam i1_2_lut_adj_1597.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_mux_3_i5_3_lut (.I0(communication_counter[4]), .I1(n29_adj_4455), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3158));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_715_3 (.CI(n28238), .I0(n1057), .I1(VCC_net), .CO(n28239));
    SB_LUT4 rem_4_add_715_2_lut (.I0(GND_net), .I1(n1058), .I2(GND_net), 
            .I3(VCC_net), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_22 (.CI(n28762), .I0(n3039), .I1(VCC_net), 
            .CO(n28763));
    SB_LUT4 rem_4_add_1988_16_lut (.I0(GND_net), .I1(n2945_adj_4439), .I2(VCC_net), 
            .I3(n28783), .O(n3012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_8_lut (.I0(GND_net), .I1(n1953), .I2(VCC_net), 
            .I3(n29036), .O(n2020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_8 (.CI(n29036), .I0(n1953), .I1(VCC_net), 
            .CO(n29037));
    SB_LUT4 rem_4_add_1318_7_lut (.I0(GND_net), .I1(n1954), .I2(GND_net), 
            .I3(n29035), .O(n2021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_16 (.CI(n28783), .I0(n2945_adj_4439), .I1(VCC_net), 
            .CO(n28784));
    SB_CARRY rem_4_add_715_2 (.CI(VCC_net), .I0(n1058), .I1(GND_net), 
            .CO(n28238));
    SB_LUT4 div_46_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1598 (.I0(n84), .I1(n15576), .I2(GND_net), .I3(GND_net), 
            .O(n15573));
    defparam i1_2_lut_adj_1598.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_add_1988_15_lut (.I0(GND_net), .I1(n2946_adj_4438), .I2(VCC_net), 
            .I3(n28782), .O(n3013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_21_lut (.I0(GND_net), .I1(n3040), .I2(VCC_net), 
            .I3(n28761), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_7 (.CI(n29035), .I0(n1954), .I1(GND_net), 
            .CO(n29036));
    SB_CARRY rem_4_add_1988_15 (.CI(n28782), .I0(n2946_adj_4438), .I1(VCC_net), 
            .CO(n28783));
    SB_LUT4 div_46_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2055_21 (.CI(n28761), .I0(n3040), .I1(VCC_net), 
            .CO(n28762));
    SB_LUT4 rem_4_add_1318_6_lut (.I0(GND_net), .I1(n1955), .I2(GND_net), 
            .I3(n29034), .O(n2022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_20_lut (.I0(GND_net), .I1(n3041), .I2(VCC_net), 
            .I3(n28760), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_20 (.CI(n28760), .I0(n3041), .I1(VCC_net), 
            .CO(n28761));
    SB_LUT4 rem_4_add_2055_19_lut (.I0(GND_net), .I1(n3042), .I2(VCC_net), 
            .I3(n28759), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_19 (.CI(n28759), .I0(n3042), .I1(VCC_net), 
            .CO(n28760));
    SB_LUT4 div_46_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1599 (.I0(n87), .I1(n15570), .I2(GND_net), .I3(GND_net), 
            .O(n15522));
    defparam i1_2_lut_adj_1599.LUT_INIT = 16'hdddd;
    SB_LUT4 rem_4_add_2055_18_lut (.I0(GND_net), .I1(n3043), .I2(VCC_net), 
            .I3(n28758), .O(n3110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_14_lut (.I0(GND_net), .I1(n2947_adj_4437), .I2(VCC_net), 
            .I3(n28781), .O(n3014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63_adj_4324), 
            .I2(gearBoxRatio[23]), .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_1988_14 (.CI(n28781), .I0(n2947_adj_4437), .I1(VCC_net), 
            .CO(n28782));
    SB_LUT4 rem_4_add_1988_13_lut (.I0(GND_net), .I1(n2948_adj_4436), .I2(VCC_net), 
            .I3(n28780), .O(n3015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_6 (.CI(n29034), .I0(n1955), .I1(GND_net), 
            .CO(n29035));
    SB_CARRY rem_4_add_1988_13 (.CI(n28780), .I0(n2948_adj_4436), .I1(VCC_net), 
            .CO(n28781));
    SB_LUT4 rem_4_add_1318_5_lut (.I0(GND_net), .I1(n1956), .I2(VCC_net), 
            .I3(n29033), .O(n2023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_18 (.CI(n28758), .I0(n3043), .I1(VCC_net), 
            .CO(n28759));
    SB_LUT4 rem_4_add_1988_12_lut (.I0(GND_net), .I1(n2949_adj_4435), .I2(VCC_net), 
            .I3(n28779), .O(n3016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_17_lut (.I0(GND_net), .I1(n3044), .I2(VCC_net), 
            .I3(n28757), .O(n3111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_17 (.CI(n28757), .I0(n3044), .I1(VCC_net), 
            .CO(n28758));
    SB_LUT4 rem_4_add_2055_16_lut (.I0(GND_net), .I1(n3045), .I2(VCC_net), 
            .I3(n28756), .O(n3112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_16 (.CI(n28756), .I0(n3045), .I1(VCC_net), 
            .CO(n28757));
    SB_CARRY rem_4_add_1318_5 (.CI(n29033), .I0(n1956), .I1(VCC_net), 
            .CO(n29034));
    SB_CARRY rem_4_add_1988_12 (.CI(n28779), .I0(n2949_adj_4435), .I1(VCC_net), 
            .CO(n28780));
    SB_LUT4 rem_4_add_1318_4_lut (.I0(GND_net), .I1(n1957), .I2(VCC_net), 
            .I3(n29032), .O(n2024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_15_lut (.I0(GND_net), .I1(n3046), .I2(VCC_net), 
            .I3(n28755), .O(n3113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_11_lut (.I0(GND_net), .I1(n2950_adj_4434), .I2(VCC_net), 
            .I3(n28778), .O(n3017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_4 (.CI(n29032), .I0(n1957), .I1(VCC_net), 
            .CO(n29033));
    SB_LUT4 div_46_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2055_15 (.CI(n28755), .I0(n3046), .I1(VCC_net), 
            .CO(n28756));
    SB_LUT4 rem_4_add_1318_3_lut (.I0(GND_net), .I1(n1958), .I2(GND_net), 
            .I3(n29031), .O(n2025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1600 (.I0(n90), .I1(n15517), .I2(GND_net), .I3(GND_net), 
            .O(n15564));
    defparam i1_2_lut_adj_1600.LUT_INIT = 16'hdddd;
    SB_CARRY rem_4_add_1988_11 (.CI(n28778), .I0(n2950_adj_4434), .I1(VCC_net), 
            .CO(n28779));
    SB_LUT4 rem_4_add_2055_14_lut (.I0(GND_net), .I1(n3047), .I2(VCC_net), 
            .I3(n28754), .O(n3114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_10_lut (.I0(GND_net), .I1(n2951_adj_4433), .I2(VCC_net), 
            .I3(n28777), .O(n3018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_14 (.CI(n28754), .I0(n3047), .I1(VCC_net), 
            .CO(n28755));
    SB_LUT4 div_46_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_1318_3 (.CI(n29031), .I0(n1958), .I1(GND_net), 
            .CO(n29032));
    SB_LUT4 rem_4_add_2055_13_lut (.I0(GND_net), .I1(n3048), .I2(VCC_net), 
            .I3(n28753), .O(n3115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2055_13 (.CI(n28753), .I0(n3048), .I1(VCC_net), 
            .CO(n28754));
    SB_LUT4 rem_4_add_2055_12_lut (.I0(GND_net), .I1(n3049), .I2(VCC_net), 
            .I3(n28752), .O(n3116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_12 (.CI(n28752), .I0(n3049), .I1(VCC_net), 
            .CO(n28753));
    SB_CARRY rem_4_add_1988_10 (.CI(n28777), .I0(n2951_adj_4433), .I1(VCC_net), 
            .CO(n28778));
    SB_LUT4 rem_4_add_2055_11_lut (.I0(GND_net), .I1(n3050), .I2(VCC_net), 
            .I3(n28751), .O(n3117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_2 (.CI(VCC_net), .I0(n2058), .I1(VCC_net), 
            .CO(n29031));
    SB_CARRY rem_4_add_2055_11 (.CI(n28751), .I0(n3050), .I1(VCC_net), 
            .CO(n28752));
    SB_LUT4 rem_4_add_1988_9_lut (.I0(GND_net), .I1(n2952_adj_4432), .I2(VCC_net), 
            .I3(n28776), .O(n3019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_19_lut (.I0(n2075_adj_4653), .I1(n2042), .I2(VCC_net), 
            .I3(n29030), .O(n2141)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1601 (.I0(n93), .I1(n15504), .I2(GND_net), .I3(GND_net), 
            .O(n15558));
    defparam i1_2_lut_adj_1601.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1602 (.I0(n96), .I1(n15498), .I2(GND_net), .I3(GND_net), 
            .O(n15494));
    defparam i1_2_lut_adj_1602.LUT_INIT = 16'hdddd;
    SB_LUT4 rem_4_add_2055_10_lut (.I0(GND_net), .I1(n3051), .I2(VCC_net), 
            .I3(n28750), .O(n3118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2055_10 (.CI(n28750), .I0(n3051), .I1(VCC_net), 
            .CO(n28751));
    SB_LUT4 div_46_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_add_2055_9_lut (.I0(GND_net), .I1(n3052), .I2(VCC_net), 
            .I3(n28749), .O(n3119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n15491), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_CARRY rem_4_add_2055_9 (.CI(n28749), .I0(n3052), .I1(VCC_net), 
            .CO(n28750));
    SB_LUT4 i36327_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n43089));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i36327_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2055_8_lut (.I0(GND_net), .I1(n3053), .I2(VCC_net), 
            .I3(n28748), .O(n3120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_mux_3_i1_3_lut (.I0(communication_counter[0]), .I1(n33_adj_4452), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3459));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i1_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2055_8 (.CI(n28748), .I0(n3053), .I1(VCC_net), 
            .CO(n28749));
    SB_LUT4 rem_4_add_1385_18_lut (.I0(GND_net), .I1(n2043), .I2(VCC_net), 
            .I3(n29029), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_7_lut (.I0(GND_net), .I1(n3054), .I2(GND_net), 
            .I3(n28747), .O(n3121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_7 (.CI(n28747), .I0(n3054), .I1(GND_net), 
            .CO(n28748));
    SB_LUT4 rem_4_add_2055_6_lut (.I0(GND_net), .I1(n3055), .I2(GND_net), 
            .I3(n28746), .O(n3122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_mux_3_i2_3_lut (.I0(communication_counter[1]), .I1(n32), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3458));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i2_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2055_6 (.CI(n28746), .I0(n3055), .I1(GND_net), 
            .CO(n28747));
    SB_LUT4 i36273_1_lut (.I0(n3457), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43037));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36273_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1385_18 (.CI(n29029), .I0(n2043), .I1(VCC_net), 
            .CO(n29030));
    SB_LUT4 rem_4_i2287_3_lut (.I0(n3358), .I1(n10087), .I2(n3362), .I3(GND_net), 
            .O(n3457));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2287_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i36270_1_lut (.I0(n3456), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43034));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36270_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2286_3_lut (.I0(n3357), .I1(n10086), .I2(n3362), .I3(GND_net), 
            .O(n3456));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2286_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i36267_1_lut (.I0(n3455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43031));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36267_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2285_3_lut (.I0(n3356), .I1(n10085), .I2(n3362), .I3(GND_net), 
            .O(n3455));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2285_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i36264_1_lut (.I0(n3454), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43028));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36264_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1988_9 (.CI(n28776), .I0(n2952_adj_4432), .I1(VCC_net), 
            .CO(n28777));
    SB_LUT4 rem_4_add_1385_17_lut (.I0(GND_net), .I1(n2044), .I2(VCC_net), 
            .I3(n29028), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_5_lut (.I0(GND_net), .I1(n3056), .I2(VCC_net), 
            .I3(n28745), .O(n3123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_17 (.CI(n29028), .I0(n2044), .I1(VCC_net), 
            .CO(n29029));
    SB_LUT4 rem_4_i2284_3_lut (.I0(n3355), .I1(n10084), .I2(n3362), .I3(GND_net), 
            .O(n3454));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2284_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_2055_5 (.CI(n28745), .I0(n3056), .I1(VCC_net), 
            .CO(n28746));
    SB_LUT4 i36261_1_lut (.I0(n3453), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43025));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36261_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2283_3_lut (.I0(n3354), .I1(n10083), .I2(n3362), .I3(GND_net), 
            .O(n3453));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2283_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i2215_3_lut (.I0(n3254), .I1(n3321), .I2(n3263), .I3(GND_net), 
            .O(n3353));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2217_3_lut (.I0(n3256), .I1(n3323), .I2(n3263), .I3(GND_net), 
            .O(n3355));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2216_3_lut (.I0(n3255), .I1(n3322), .I2(n3263), .I3(GND_net), 
            .O(n3354));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2055_4_lut (.I0(GND_net), .I1(n3057), .I2(VCC_net), 
            .I3(n28744), .O(n3124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_16_lut (.I0(GND_net), .I1(n2045), .I2(VCC_net), 
            .I3(n29027), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_mux_3_i3_3_lut (.I0(communication_counter[2]), .I1(n31_adj_4453), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3358));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2219_3_lut (.I0(n3258), .I1(n3325), .I2(n3263), .I3(GND_net), 
            .O(n3357));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY rem_4_add_2055_4 (.CI(n28744), .I0(n3057), .I1(VCC_net), 
            .CO(n28745));
    SB_LUT4 rem_4_add_1988_8_lut (.I0(GND_net), .I1(n2953_adj_4431), .I2(VCC_net), 
            .I3(n28775), .O(n3020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_3_lut (.I0(GND_net), .I1(n3058), .I2(GND_net), 
            .I3(n28743), .O(n3125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i2218_3_lut (.I0(n3257), .I1(n3324), .I2(n3263), .I3(GND_net), 
            .O(n3356));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2218_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_3 (.CI(n28743), .I0(n3058), .I1(GND_net), 
            .CO(n28744));
    SB_LUT4 rem_4_i2212_3_lut (.I0(n3251), .I1(n3318), .I2(n3263), .I3(GND_net), 
            .O(n3350));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2213_3_lut (.I0(n3252), .I1(n3319), .I2(n3263), .I3(GND_net), 
            .O(n3351));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2206_3_lut (.I0(n3245), .I1(n3312), .I2(n3263), .I3(GND_net), 
            .O(n3344));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12592_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n13195), .I3(GND_net), .O(n17274));   // verilog/coms.v(126[12] 289[6])
    defparam i12592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2208_3_lut (.I0(n3247), .I1(n3314), .I2(n3263), .I3(GND_net), 
            .O(n3346));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1603 (.I0(n3249), .I1(n3350), .I2(n3316), .I3(n3263), 
            .O(n37650));
    defparam i1_4_lut_adj_1603.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1604 (.I0(n3242), .I1(n3351), .I2(n3309), .I3(n3263), 
            .O(n37648));
    defparam i1_4_lut_adj_1604.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2201_3_lut (.I0(n3240), .I1(n3307), .I2(n3263), .I3(GND_net), 
            .O(n3339));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2200_3_lut (.I0(n3239), .I1(n3306), .I2(n3263), .I3(GND_net), 
            .O(n3338));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1605 (.I0(n3338), .I1(n3339), .I2(n37648), .I3(n37650), 
            .O(n37656));
    defparam i1_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2204_3_lut (.I0(n3243), .I1(n3310), .I2(n3263), .I3(GND_net), 
            .O(n3342));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2214_3_lut (.I0(n3253), .I1(n3320), .I2(n3263), .I3(GND_net), 
            .O(n3352));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1606 (.I0(n3244), .I1(n3344), .I2(n3311), .I3(n3263), 
            .O(n37576));
    defparam i1_4_lut_adj_1606.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2202_3_lut (.I0(n3241), .I1(n3308), .I2(n3263), .I3(GND_net), 
            .O(n3340));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1607 (.I0(n3246), .I1(n3342), .I2(n3313), .I3(n3263), 
            .O(n37578));
    defparam i1_4_lut_adj_1607.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_3_lut (.I0(n3356), .I1(n3357), .I2(n3358), .I3(GND_net), 
            .O(n35648));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1608 (.I0(n37578), .I1(n3340), .I2(n37576), .I3(n3352), 
            .O(n37584));
    defparam i1_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_2055_2 (.CI(VCC_net), .I0(n3158), .I1(VCC_net), 
            .CO(n28743));
    SB_CARRY rem_4_add_1988_8 (.CI(n28775), .I0(n2953_adj_4431), .I1(VCC_net), 
            .CO(n28776));
    SB_CARRY rem_4_add_1385_16 (.CI(n29027), .I0(n2045), .I1(VCC_net), 
            .CO(n29028));
    SB_LUT4 i12899_3_lut (.I0(setpoint[8]), .I1(n4300), .I2(n36839), .I3(GND_net), 
            .O(n17581));   // verilog/coms.v(126[12] 289[6])
    defparam i12899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24_3_lut (.I0(n40171), .I1(bit_ctr[8]), .I2(n4385), .I3(GND_net), 
            .O(n33323));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut (.I0(bit_ctr[7]), .I1(n40199), .I2(n4385), .I3(GND_net), 
            .O(n33385));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1609 (.I0(bit_ctr[6]), .I1(n40198), .I2(n4385), 
            .I3(GND_net), .O(n33383));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1609.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1610 (.I0(bit_ctr[5]), .I1(n40197), .I2(n4385), 
            .I3(GND_net), .O(n33381));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1610.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1385_15_lut (.I0(GND_net), .I1(n2046), .I2(VCC_net), 
            .I3(n29026), .O(n2113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1611 (.I0(n3354), .I1(n37584), .I2(n35648), .I3(n3355), 
            .O(n37586));
    defparam i1_4_lut_adj_1611.LUT_INIT = 16'heccc;
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_7_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b000001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_4_lut_adj_1612 (.I0(n3237), .I1(n37586), .I2(n3304), .I3(n3263), 
            .O(n37588));
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_add_1988_7_lut (.I0(GND_net), .I1(n2954_adj_4430), .I2(GND_net), 
            .I3(n28774), .O(n3021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_3 (.CI(n28770), .I0(n2958_adj_4426), .I1(GND_net), 
            .CO(n28771));
    SB_LUT4 i1_4_lut_adj_1613 (.I0(n3236), .I1(n37656), .I2(n3303), .I3(n3263), 
            .O(n37658));
    defparam i1_4_lut_adj_1613.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(n3353), .I1(n3250), .I2(n3317), .I3(n3263), 
            .O(n37690));
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'hfaee;
    SB_LUT4 rem_4_add_648_7_lut (.I0(n986), .I1(n953), .I2(VCC_net), .I3(n28229), 
            .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1385_15 (.CI(n29026), .I0(n2046), .I1(VCC_net), 
            .CO(n29027));
    SB_LUT4 i3_4_lut (.I0(n3248), .I1(n3346), .I2(n3315), .I3(n3263), 
            .O(n28_adj_5008));
    defparam i3_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1615 (.I0(n37658), .I1(n3235), .I2(n3302), .I3(n3263), 
            .O(n46_adj_5005));
    defparam i1_4_lut_adj_1615.LUT_INIT = 16'hfaee;
    SB_LUT4 rem_4_i1331_3_lut (.I0(n1954), .I1(n2021), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2053));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_14_lut (.I0(GND_net), .I1(n2047), .I2(VCC_net), 
            .I3(n29025), .O(n2114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1327_3_lut (.I0(n1950), .I1(n2017), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2049));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_648_6_lut (.I0(GND_net), .I1(n954), .I2(GND_net), 
            .I3(n28228), .O(n1021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1616 (.I0(n37588), .I1(n3233), .I2(n3300), .I3(n3263), 
            .O(n47_adj_5004));
    defparam i1_4_lut_adj_1616.LUT_INIT = 16'hfaee;
    SB_LUT4 rem_4_i2199_3_lut (.I0(n3238), .I1(n3305), .I2(n3263), .I3(GND_net), 
            .O(n3337));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1617 (.I0(n3234), .I1(n3337), .I2(n3301), .I3(n3263), 
            .O(n37460));
    defparam i1_4_lut_adj_1617.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2192_3_lut (.I0(n3231), .I1(n3298), .I2(n3263), .I3(GND_net), 
            .O(n3330));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1618 (.I0(n47_adj_5004), .I1(n46_adj_5005), .I2(n28_adj_5008), 
            .I3(n37690), .O(n37696));
    defparam i1_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1619 (.I0(n3232), .I1(n37460), .I2(n3299), .I3(n3263), 
            .O(n37462));
    defparam i1_4_lut_adj_1619.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1620 (.I0(n37992), .I1(n37462), .I2(n37696), 
            .I3(n3330), .O(n3362));
    defparam i1_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i36260_2_lut (.I0(n3362), .I1(n10082), .I2(GND_net), .I3(GND_net), 
            .O(n3452));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36260_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i32_1_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4965));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1328_3_lut (.I0(n1951), .I1(n2018), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2050));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[6]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_106[6]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_648_6 (.CI(n28228), .I0(n954), .I1(GND_net), .CO(n28229));
    SB_LUT4 rem_4_i1329_3_lut (.I0(n1952), .I1(n2019), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2051));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1329_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_14 (.CI(n29025), .I0(n2047), .I1(VCC_net), 
            .CO(n29026));
    SB_LUT4 rem_4_add_1385_13_lut (.I0(GND_net), .I1(n2048), .I2(VCC_net), 
            .I3(n29024), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_71_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[7]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY rem_4_add_1385_13 (.CI(n29024), .I0(n2048), .I1(VCC_net), 
            .CO(n29025));
    SB_LUT4 i22_3_lut_adj_1621 (.I0(bit_ctr[4]), .I1(n40196), .I2(n4385), 
            .I3(GND_net), .O(n33379));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1621.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1988_7 (.CI(n28774), .I0(n2954_adj_4430), .I1(GND_net), 
            .CO(n28775));
    SB_LUT4 rem_4_add_1385_12_lut (.I0(GND_net), .I1(n2049), .I2(VCC_net), 
            .I3(n29023), .O(n2116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1622 (.I0(bit_ctr[3]), .I1(n40195), .I2(n4385), 
            .I3(GND_net), .O(n33377));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1622.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_106[7]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1623 (.I0(bit_ctr[0]), .I1(n40177), .I2(n4385), 
            .I3(GND_net), .O(n33335));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1623.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1321_3_lut (.I0(n1944), .I1(n2011), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2043));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[8]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_106[8]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1330_3_lut (.I0(n1953), .I1(n2020), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2052));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1325_3_lut (.I0(n1948), .I1(n2015), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2047));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[9]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_106[9]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_12 (.CI(n29023), .I0(n2049), .I1(VCC_net), 
            .CO(n29024));
    SB_LUT4 rem_4_add_1385_11_lut (.I0(GND_net), .I1(n2050), .I2(VCC_net), 
            .I3(n29022), .O(n2117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1323_3_lut (.I0(n1946), .I1(n2013), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2045));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_11 (.CI(n29022), .I0(n2050), .I1(VCC_net), 
            .CO(n29023));
    SB_LUT4 rem_4_add_1385_10_lut (.I0(GND_net), .I1(n2051), .I2(VCC_net), 
            .I3(n29021), .O(n2118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_71_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[10]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY rem_4_add_1385_10 (.CI(n29021), .I0(n2051), .I1(VCC_net), 
            .CO(n29022));
    SB_LUT4 mux_70_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_106[10]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_9_lut (.I0(GND_net), .I1(n2052), .I2(VCC_net), 
            .I3(n29020), .O(n2119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_9 (.CI(n29020), .I0(n2052), .I1(VCC_net), 
            .CO(n29021));
    SB_LUT4 rem_4_add_1385_8_lut (.I0(GND_net), .I1(n2053), .I2(VCC_net), 
            .I3(n29019), .O(n2120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1324_3_lut (.I0(n1947), .I1(n2014), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2046));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_8 (.CI(n29019), .I0(n2053), .I1(VCC_net), 
            .CO(n29020));
    SB_LUT4 rem_4_add_1385_7_lut (.I0(GND_net), .I1(n2054), .I2(GND_net), 
            .I3(n29018), .O(n2121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1322_3_lut (.I0(n1945), .I1(n2012), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2044));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1333_3_lut (.I0(n1956), .I1(n2023), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2055));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1333_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_7 (.CI(n29018), .I0(n2054), .I1(GND_net), 
            .CO(n29019));
    SB_LUT4 rem_4_add_1385_6_lut (.I0(GND_net), .I1(n2055), .I2(GND_net), 
            .I3(n29017), .O(n2122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_6 (.CI(n29017), .I0(n2055), .I1(GND_net), 
            .CO(n29018));
    SB_LUT4 rem_4_add_1385_5_lut (.I0(GND_net), .I1(n2056), .I2(VCC_net), 
            .I3(n29016), .O(n2123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12615_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17297));   // verilog/coms.v(126[12] 289[6])
    defparam i12615_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12616_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17298));   // verilog/coms.v(126[12] 289[6])
    defparam i12616_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_71_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[11]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_106[11]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_5 (.CI(n29016), .I0(n2056), .I1(VCC_net), 
            .CO(n29017));
    SB_LUT4 rem_4_add_648_5_lut (.I0(GND_net), .I1(n955), .I2(GND_net), 
            .I3(n28227), .O(n1022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1326_3_lut (.I0(n1949), .I1(n2016), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2048));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[12]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_106[12]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_4_lut (.I0(GND_net), .I1(n2057), .I2(VCC_net), 
            .I3(n29015), .O(n2124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_71_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[13]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_106[13]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_4 (.CI(n29015), .I0(n2057), .I1(VCC_net), 
            .CO(n29016));
    SB_LUT4 i12617_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17299));   // verilog/coms.v(126[12] 289[6])
    defparam i12617_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12618_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17300));   // verilog/coms.v(126[12] 289[6])
    defparam i12618_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1332_3_lut (.I0(n1955), .I1(n2022), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2054));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_3_lut (.I0(GND_net), .I1(n2058), .I2(GND_net), 
            .I3(n29014), .O(n2125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_5 (.CI(n28227), .I0(n955), .I1(GND_net), .CO(n28228));
    SB_CARRY rem_4_add_1385_3 (.CI(n29014), .I0(n2058), .I1(GND_net), 
            .CO(n29015));
    SB_CARRY rem_4_add_1385_2 (.CI(VCC_net), .I0(n2158), .I1(VCC_net), 
            .CO(n29014));
    SB_LUT4 rem_4_add_1452_20_lut (.I0(n2174_adj_4638), .I1(n2141), .I2(VCC_net), 
            .I3(n29013), .O(n2240)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12619_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17301));   // verilog/coms.v(126[12] 289[6])
    defparam i12619_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_648_4_lut (.I0(GND_net), .I1(n956), .I2(VCC_net), 
            .I3(n28226), .O(n1023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_4_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i12620_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17302));   // verilog/coms.v(126[12] 289[6])
    defparam i12620_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12621_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17303));   // verilog/coms.v(126[12] 289[6])
    defparam i12621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1452_19_lut (.I0(GND_net), .I1(n2142), .I2(VCC_net), 
            .I3(n29012), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_4 (.CI(n28226), .I0(n956), .I1(VCC_net), .CO(n28227));
    SB_LUT4 rem_4_i1335_3_lut (.I0(n1958), .I1(n2025), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2057));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1335_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_19 (.CI(n29012), .I0(n2142), .I1(VCC_net), 
            .CO(n29013));
    SB_LUT4 rem_4_add_1452_18_lut (.I0(GND_net), .I1(n2143), .I2(VCC_net), 
            .I3(n29011), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF h1_55 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 rem_4_i1334_rep_44_3_lut (.I0(n1957), .I1(n2024), .I2(n1976_adj_4689), 
            .I3(GND_net), .O(n2056));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1334_rep_44_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1624 (.I0(n2056), .I1(n2057), .I2(n2058), .I3(GND_net), 
            .O(n35627));
    defparam i1_3_lut_adj_1624.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n2054), .I1(n2048), .I2(n35627), .I3(n2055), 
            .O(n17_adj_4363));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i27_3_lut (.I0(n1163), .I1(n35361), .I2(state[0]), .I3(GND_net), 
            .O(n19_adj_4920));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i22_3_lut_adj_1625 (.I0(bit_ctr[30]), .I1(n40191), .I2(n4385), 
            .I3(GND_net), .O(n33369));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1625.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1626 (.I0(bit_ctr[29]), .I1(n40190), .I2(n4385), 
            .I3(GND_net), .O(n33367));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1626.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i27_3_lut (.I0(communication_counter[26]), .I1(n7_adj_4510), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n958));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i655_3_lut (.I0(n958), .I1(n1025), .I2(n986), .I3(GND_net), 
            .O(n1057));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut (.I0(n2044), .I1(n2046), .I2(n2045), .I3(n2047), 
            .O(n21_adj_4361));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1452_18 (.CI(n29011), .I0(n2143), .I1(VCC_net), 
            .CO(n29012));
    SB_LUT4 rem_4_add_1452_17_lut (.I0(GND_net), .I1(n2144), .I2(VCC_net), 
            .I3(n29010), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_17 (.CI(n29010), .I0(n2144), .I1(VCC_net), 
            .CO(n29011));
    SB_LUT4 rem_4_add_1452_16_lut (.I0(GND_net), .I1(n2145), .I2(VCC_net), 
            .I3(n29009), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_3_lut (.I0(n2052), .I1(n2043), .I2(n2042), .I3(GND_net), 
            .O(n20_adj_4362));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n21_adj_4361), .I1(n17_adj_4363), .I2(n2049), 
            .I3(n2053), .O(n24_adj_4360));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1452_16 (.CI(n29009), .I0(n2145), .I1(VCC_net), 
            .CO(n29010));
    SB_LUT4 rem_4_add_1452_15_lut (.I0(GND_net), .I1(n2146), .I2(VCC_net), 
            .I3(n29008), .O(n2213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_15 (.CI(n29008), .I0(n2146), .I1(VCC_net), 
            .CO(n29009));
    SB_LUT4 rem_4_add_2122_30_lut (.I0(n3164), .I1(n3131), .I2(VCC_net), 
            .I3(n28719), .O(n3230)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_2122_29_lut (.I0(GND_net), .I1(n3132), .I2(VCC_net), 
            .I3(n28718), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_29 (.CI(n28718), .I0(n3132), .I1(VCC_net), 
            .CO(n28719));
    SB_LUT4 rem_4_add_2122_28_lut (.I0(GND_net), .I1(n3133), .I2(VCC_net), 
            .I3(n28717), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_14_lut (.I0(GND_net), .I1(n2147), .I2(VCC_net), 
            .I3(n29007), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i970_3_lut_3_lut (.I0(n1436), .I1(n5846), .I2(n1420), 
            .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i970_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_28 (.CI(n28717), .I0(n3133), .I1(VCC_net), 
            .CO(n28718));
    SB_LUT4 rem_4_add_2122_27_lut (.I0(GND_net), .I1(n3134), .I2(VCC_net), 
            .I3(n28716), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_27 (.CI(n28716), .I0(n3134), .I1(VCC_net), 
            .CO(n28717));
    SB_CARRY rem_4_add_1452_14 (.CI(n29007), .I0(n2147), .I1(VCC_net), 
            .CO(n29008));
    SB_LUT4 i12_4_lut (.I0(n2051), .I1(n24_adj_4360), .I2(n20_adj_4362), 
            .I3(n2050), .O(n2075_adj_4653));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i964_3_lut_3_lut (.I0(n1436), .I1(n5840), .I2(n1414), 
            .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i964_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1627 (.I0(bit_ctr[28]), .I1(n40189), .I2(n4385), 
            .I3(GND_net), .O(n33365));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1627.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1628 (.I0(bit_ctr[27]), .I1(n40188), .I2(n4385), 
            .I3(GND_net), .O(n33363));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1628.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2122_26_lut (.I0(GND_net), .I1(n3135), .I2(VCC_net), 
            .I3(n28715), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_13_lut (.I0(GND_net), .I1(n2148), .I2(VCC_net), 
            .I3(n29006), .O(n2215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_13 (.CI(n29006), .I0(n2148), .I1(VCC_net), 
            .CO(n29007));
    SB_LUT4 rem_4_add_1452_12_lut (.I0(GND_net), .I1(n2149), .I2(VCC_net), 
            .I3(n29005), .O(n2216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_26 (.CI(n28715), .I0(n3135), .I1(VCC_net), 
            .CO(n28716));
    SB_LUT4 rem_4_add_2122_25_lut (.I0(GND_net), .I1(n3136), .I2(VCC_net), 
            .I3(n28714), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_25 (.CI(n28714), .I0(n3136), .I1(VCC_net), 
            .CO(n28715));
    SB_CARRY rem_4_add_1452_12 (.CI(n29005), .I0(n2149), .I1(VCC_net), 
            .CO(n29006));
    SB_LUT4 rem_4_add_2122_24_lut (.I0(GND_net), .I1(n3137), .I2(VCC_net), 
            .I3(n28713), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i968_3_lut_3_lut (.I0(n1436), .I1(n5844), .I2(n1418), 
            .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i968_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1452_11_lut (.I0(GND_net), .I1(n2150), .I2(VCC_net), 
            .I3(n29004), .O(n2217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_24 (.CI(n28713), .I0(n3137), .I1(VCC_net), 
            .CO(n28714));
    SB_LUT4 rem_4_add_2122_23_lut (.I0(GND_net), .I1(n3138), .I2(VCC_net), 
            .I3(n28712), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i969_3_lut_3_lut (.I0(n1436), .I1(n5845), .I2(n1419), 
            .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i969_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i967_3_lut_3_lut (.I0(n1436), .I1(n5843), .I2(n1417), 
            .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i967_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_23 (.CI(n28712), .I0(n3138), .I1(VCC_net), 
            .CO(n28713));
    SB_CARRY rem_4_add_1452_11 (.CI(n29004), .I0(n2150), .I1(VCC_net), 
            .CO(n29005));
    SB_LUT4 rem_4_add_1452_10_lut (.I0(GND_net), .I1(n2151), .I2(VCC_net), 
            .I3(n29003), .O(n2218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_22_lut (.I0(GND_net), .I1(n3139), .I2(VCC_net), 
            .I3(n28711), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_22 (.CI(n28711), .I0(n3139), .I1(VCC_net), 
            .CO(n28712));
    SB_LUT4 rem_4_add_2122_21_lut (.I0(GND_net), .I1(n3140), .I2(VCC_net), 
            .I3(n28710), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_21 (.CI(n28710), .I0(n3140), .I1(VCC_net), 
            .CO(n28711));
    SB_LUT4 rem_4_add_2122_20_lut (.I0(GND_net), .I1(n3141), .I2(VCC_net), 
            .I3(n28709), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_20 (.CI(n28709), .I0(n3141), .I1(VCC_net), 
            .CO(n28710));
    SB_LUT4 rem_4_add_2122_19_lut (.I0(GND_net), .I1(n3142), .I2(VCC_net), 
            .I3(n28708), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_19 (.CI(n28708), .I0(n3142), .I1(VCC_net), 
            .CO(n28709));
    SB_CARRY rem_4_add_1452_10 (.CI(n29003), .I0(n2151), .I1(VCC_net), 
            .CO(n29004));
    SB_LUT4 rem_4_add_2122_18_lut (.I0(GND_net), .I1(n3143), .I2(VCC_net), 
            .I3(n28707), .O(n3210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_80[23]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_CARRY rem_4_add_2122_18 (.CI(n28707), .I0(n3143), .I1(VCC_net), 
            .CO(n28708));
    SB_LUT4 rem_4_add_2122_17_lut (.I0(GND_net), .I1(n3144), .I2(VCC_net), 
            .I3(n28706), .O(n3211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i963_3_lut_3_lut (.I0(n1436), .I1(n5839), .I2(n1413), 
            .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i963_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_17 (.CI(n28706), .I0(n3144), .I1(VCC_net), 
            .CO(n28707));
    SB_LUT4 rem_4_add_1452_9_lut (.I0(GND_net), .I1(n2152), .I2(VCC_net), 
            .I3(n29002), .O(n2219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_9 (.CI(n29002), .I0(n2152), .I1(VCC_net), 
            .CO(n29003));
    SB_LUT4 rem_4_add_1452_8_lut (.I0(GND_net), .I1(n2153), .I2(VCC_net), 
            .I3(n29001), .O(n2220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_16_lut (.I0(GND_net), .I1(n3145), .I2(VCC_net), 
            .I3(n28705), .O(n3212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_648_3_lut (.I0(GND_net), .I1(n957), .I2(VCC_net), 
            .I3(n28225), .O(n1024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_8 (.CI(n29001), .I0(n2153), .I1(VCC_net), 
            .CO(n29002));
    SB_LUT4 div_46_i971_3_lut_3_lut (.I0(n1436), .I1(n5847), .I2(n656), 
            .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i971_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1452_7_lut (.I0(GND_net), .I1(n2154), .I2(GND_net), 
            .I3(n29000), .O(n2221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_16 (.CI(n28705), .I0(n3145), .I1(VCC_net), 
            .CO(n28706));
    SB_CARRY rem_4_add_648_3 (.CI(n28225), .I0(n957), .I1(VCC_net), .CO(n28226));
    SB_CARRY rem_4_add_1452_7 (.CI(n29000), .I0(n2154), .I1(GND_net), 
            .CO(n29001));
    SB_LUT4 rem_4_add_648_2_lut (.I0(GND_net), .I1(n958), .I2(GND_net), 
            .I3(VCC_net), .O(n1025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i966_3_lut_3_lut (.I0(n1436), .I1(n5842), .I2(n1416), 
            .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i966_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_648_2 (.CI(VCC_net), .I0(n958), .I1(GND_net), .CO(n28225));
    SB_LUT4 div_46_i965_3_lut_3_lut (.I0(n1436), .I1(n5841), .I2(n1415), 
            .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i965_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1452_6_lut (.I0(GND_net), .I1(n2155), .I2(GND_net), 
            .I3(n28999), .O(n2222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_15_lut (.I0(GND_net), .I1(n3146), .I2(VCC_net), 
            .I3(n28704), .O(n3213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_6 (.CI(n28999), .I0(n2155), .I1(GND_net), 
            .CO(n29000));
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_229[23]), 
            .I2(n3_adj_4380), .I3(n28224), .O(displacement_23__N_80[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i962_3_lut_3_lut (.I0(n1436), .I1(n5838), .I2(n1412), 
            .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i962_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1452_5_lut (.I0(GND_net), .I1(n2156), .I2(VCC_net), 
            .I3(n28998), .O(n2223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_229[22]), 
            .I2(n3_adj_4380), .I3(n28223), .O(displacement_23__N_80[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_5 (.CI(n28998), .I0(n2156), .I1(VCC_net), 
            .CO(n28999));
    SB_LUT4 i33584_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n40346));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33584_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_mux_3_i16_3_lut (.I0(communication_counter[15]), .I1(n18_adj_4465), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2058));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_4_lut (.I0(GND_net), .I1(n2157), .I2(VCC_net), 
            .I3(n28997), .O(n2224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_4 (.CI(n28997), .I0(n2157), .I1(VCC_net), 
            .CO(n28998));
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n28223), .I0(displacement_23__N_229[22]), 
            .I1(n3_adj_4380), .CO(n28224));
    SB_LUT4 div_46_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4648));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1048_3_lut_3_lut (.I0(n1553), .I1(n5859), .I2(n1538), 
            .I3(GND_net), .O(n1652));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1048_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12593_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n13195), .I3(GND_net), .O(n17275));   // verilog/coms.v(126[12] 289[6])
    defparam i12593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_3_lut (.I0(GND_net), .I1(n2158), .I2(GND_net), 
            .I3(n28996), .O(n2225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_229[21]), 
            .I2(n3_adj_4380), .I3(n28222), .O(displacement_23__N_80[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1042_3_lut_3_lut (.I0(n1553), .I1(n5853), .I2(n1532), 
            .I3(GND_net), .O(n1646));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1042_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1452_3 (.CI(n28996), .I0(n2158), .I1(GND_net), 
            .CO(n28997));
    SB_LUT4 div_46_i1046_3_lut_3_lut (.I0(n1553), .I1(n5857), .I2(n1536), 
            .I3(GND_net), .O(n1650));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1046_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_15 (.CI(n28704), .I0(n3146), .I1(VCC_net), 
            .CO(n28705));
    SB_LUT4 rem_4_add_2122_14_lut (.I0(GND_net), .I1(n3147), .I2(VCC_net), 
            .I3(n28703), .O(n3214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_14 (.CI(n28703), .I0(n3147), .I1(VCC_net), 
            .CO(n28704));
    SB_LUT4 div_46_i1047_3_lut_3_lut (.I0(n1553), .I1(n5858), .I2(n1537), 
            .I3(GND_net), .O(n1651));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1047_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2122_13_lut (.I0(GND_net), .I1(n3148), .I2(VCC_net), 
            .I3(n28702), .O(n3215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_2 (.CI(VCC_net), .I0(n2258), .I1(VCC_net), 
            .CO(n28996));
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n28222), .I0(displacement_23__N_229[21]), 
            .I1(n3_adj_4380), .CO(n28223));
    SB_CARRY rem_4_add_2122_13 (.CI(n28702), .I0(n3148), .I1(VCC_net), 
            .CO(n28703));
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_229[20]), 
            .I2(n3_adj_4380), .I3(n28221), .O(displacement_23__N_80[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1045_3_lut_3_lut (.I0(n1553), .I1(n5856), .I2(n1535), 
            .I3(GND_net), .O(n1649));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1045_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1041_3_lut_3_lut (.I0(n1553), .I1(n5852), .I2(n1531), 
            .I3(GND_net), .O(n1645));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1041_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1049_3_lut_3_lut (.I0(n1553), .I1(n5860), .I2(n657), 
            .I3(GND_net), .O(n1653));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1049_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1044_3_lut_3_lut (.I0(n1553), .I1(n5855), .I2(n1534), 
            .I3(GND_net), .O(n1648));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1044_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1519_21_lut (.I0(n2273_adj_4629), .I1(n2240), .I2(VCC_net), 
            .I3(n28995), .O(n2339)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n28221), .I0(displacement_23__N_229[20]), 
            .I1(n3_adj_4380), .CO(n28222));
    SB_LUT4 rem_4_add_1519_20_lut (.I0(GND_net), .I1(n2241), .I2(VCC_net), 
            .I3(n28994), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_20 (.CI(n28994), .I0(n2241), .I1(VCC_net), 
            .CO(n28995));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_229[19]), 
            .I2(n6_adj_4371), .I3(n28220), .O(displacement_23__N_80[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_19_lut (.I0(GND_net), .I1(n2242), .I2(VCC_net), 
            .I3(n28993), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_12_lut (.I0(GND_net), .I1(n3149), .I2(VCC_net), 
            .I3(n28701), .O(n3216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_12 (.CI(n28701), .I0(n3149), .I1(VCC_net), 
            .CO(n28702));
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n28220), .I0(displacement_23__N_229[19]), 
            .I1(n6_adj_4371), .CO(n28221));
    SB_CARRY rem_4_add_1519_19 (.CI(n28993), .I0(n2242), .I1(VCC_net), 
            .CO(n28994));
    SB_LUT4 div_46_i1043_3_lut_3_lut (.I0(n1553), .I1(n5854), .I2(n1533), 
            .I3(GND_net), .O(n1647));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1043_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1040_3_lut_3_lut (.I0(n1553), .I1(n5851), .I2(n1530), 
            .I3(GND_net), .O(n1644));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1040_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1519_18_lut (.I0(GND_net), .I1(n2243), .I2(VCC_net), 
            .I3(n28992), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_229[18]), 
            .I2(n7_adj_4370), .I3(n28219), .O(displacement_23__N_80[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_18 (.CI(n28992), .I0(n2243), .I1(VCC_net), 
            .CO(n28993));
    SB_LUT4 rem_4_add_1519_17_lut (.I0(GND_net), .I1(n2244), .I2(VCC_net), 
            .I3(n28991), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1039_3_lut_3_lut (.I0(n1553), .I1(n5850), .I2(n1529), 
            .I3(GND_net), .O(n1643));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1039_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1124_3_lut_3_lut (.I0(n1667), .I1(n5873), .I2(n1653), 
            .I3(GND_net), .O(n1764));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1124_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1118_3_lut_3_lut (.I0(n1667), .I1(n5867), .I2(n1647), 
            .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1118_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n28219), .I0(displacement_23__N_229[18]), 
            .I1(n7_adj_4370), .CO(n28220));
    SB_CARRY rem_4_add_1519_17 (.CI(n28991), .I0(n2244), .I1(VCC_net), 
            .CO(n28992));
    SB_LUT4 rem_4_add_1519_16_lut (.I0(GND_net), .I1(n2245), .I2(VCC_net), 
            .I3(n28990), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_16 (.CI(n28990), .I0(n2245), .I1(VCC_net), 
            .CO(n28991));
    SB_LUT4 rem_4_add_2122_11_lut (.I0(GND_net), .I1(n3150), .I2(VCC_net), 
            .I3(n28700), .O(n3217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_229[17]), 
            .I2(n8_adj_4369), .I3(n28218), .O(displacement_23__N_80[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1123_3_lut_3_lut (.I0(n1667), .I1(n5872), .I2(n1652), 
            .I3(GND_net), .O(n1763));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1123_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1122_3_lut_3_lut (.I0(n1667), .I1(n5871), .I2(n1651), 
            .I3(GND_net), .O(n1762));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1122_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1519_15_lut (.I0(GND_net), .I1(n2246), .I2(VCC_net), 
            .I3(n28989), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_11 (.CI(n28700), .I0(n3150), .I1(VCC_net), 
            .CO(n28701));
    SB_LUT4 rem_4_add_2122_10_lut (.I0(GND_net), .I1(n3151), .I2(VCC_net), 
            .I3(n28699), .O(n3218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_10 (.CI(n28699), .I0(n3151), .I1(VCC_net), 
            .CO(n28700));
    SB_LUT4 div_46_i1121_3_lut_3_lut (.I0(n1667), .I1(n5870), .I2(n1650), 
            .I3(GND_net), .O(n1761));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1121_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1117_3_lut_3_lut (.I0(n1667), .I1(n5866), .I2(n1646), 
            .I3(GND_net), .O(n1757));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1117_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1125_3_lut_3_lut (.I0(n1667), .I1(n5874), .I2(n658), 
            .I3(GND_net), .O(n1765));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1125_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1519_15 (.CI(n28989), .I0(n2246), .I1(VCC_net), 
            .CO(n28990));
    SB_LUT4 rem_4_add_2122_9_lut (.I0(GND_net), .I1(n3152), .I2(VCC_net), 
            .I3(n28698), .O(n3219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_14_lut (.I0(GND_net), .I1(n2247), .I2(VCC_net), 
            .I3(n28988), .O(n2314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_9 (.CI(n28698), .I0(n3152), .I1(VCC_net), 
            .CO(n28699));
    SB_LUT4 rem_4_add_2122_8_lut (.I0(GND_net), .I1(n3153), .I2(VCC_net), 
            .I3(n28697), .O(n3220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23264_2_lut (.I0(n855), .I1(n884), .I2(GND_net), .I3(GND_net), 
            .O(n957));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i23264_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rem_4_i654_3_lut (.I0(n957), .I1(n1024), .I2(n986), .I3(GND_net), 
            .O(n1056));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[14]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_106[14]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1120_3_lut_3_lut (.I0(n1667), .I1(n5869), .I2(n1649), 
            .I3(GND_net), .O(n1760));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1120_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1519_14 (.CI(n28988), .I0(n2247), .I1(VCC_net), 
            .CO(n28989));
    SB_CARRY rem_4_add_2122_8 (.CI(n28697), .I0(n3153), .I1(VCC_net), 
            .CO(n28698));
    SB_LUT4 mux_71_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[15]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 rem_4_add_1519_13_lut (.I0(GND_net), .I1(n2248), .I2(VCC_net), 
            .I3(n28987), .O(n2315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1119_3_lut_3_lut (.I0(n1667), .I1(n5868), .I2(n1648), 
            .I3(GND_net), .O(n1759));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1119_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_70_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_106[15]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_7_lut (.I0(GND_net), .I1(n3154), .I2(GND_net), 
            .I3(n28696), .O(n3221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_13 (.CI(n28987), .I0(n2248), .I1(VCC_net), 
            .CO(n28988));
    SB_LUT4 rem_4_i586_3_lut (.I0(n749), .I1(n855), .I2(n884), .I3(GND_net), 
            .O(n956));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i586_3_lut.LUT_INIT = 16'h9a9a;
    SB_LUT4 rem_4_i653_3_lut (.I0(n956), .I1(n1023), .I2(n986), .I3(GND_net), 
            .O(n1055));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_12_lut (.I0(GND_net), .I1(n2249), .I2(VCC_net), 
            .I3(n28986), .O(n2316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_7 (.CI(n28696), .I0(n3154), .I1(GND_net), 
            .CO(n28697));
    SB_LUT4 rem_4_add_2122_6_lut (.I0(GND_net), .I1(n3155), .I2(GND_net), 
            .I3(n28695), .O(n3222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_6 (.CI(n28695), .I0(n3155), .I1(GND_net), 
            .CO(n28696));
    SB_LUT4 rem_4_add_2122_5_lut (.I0(GND_net), .I1(n3156), .I2(VCC_net), 
            .I3(n28694), .O(n3223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1115_3_lut_3_lut (.I0(n1667), .I1(n5864), .I2(n1644), 
            .I3(GND_net), .O(n1755));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1115_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_5 (.CI(n28694), .I0(n3156), .I1(VCC_net), 
            .CO(n28695));
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_105));   // verilog/TinyFPGA_B.v(207[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1116_3_lut_3_lut (.I0(n1667), .I1(n5865), .I2(n1645), 
            .I3(GND_net), .O(n1756));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1116_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1114_3_lut_3_lut (.I0(n1667), .I1(n5863), .I2(n1643), 
            .I3(GND_net), .O(n1754));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1114_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1519_12 (.CI(n28986), .I0(n2249), .I1(VCC_net), 
            .CO(n28987));
    SB_LUT4 rem_4_add_2122_4_lut (.I0(GND_net), .I1(n3157), .I2(VCC_net), 
            .I3(n28693), .O(n3224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_11_lut (.I0(GND_net), .I1(n2250), .I2(VCC_net), 
            .I3(n28985), .O(n2317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_11 (.CI(n28985), .I0(n2250), .I1(VCC_net), 
            .CO(n28986));
    SB_CARRY rem_4_add_2122_4 (.CI(n28693), .I0(n3157), .I1(VCC_net), 
            .CO(n28694));
    SB_LUT4 rem_4_add_2122_3_lut (.I0(GND_net), .I1(n3158), .I2(GND_net), 
            .I3(n28692), .O(n3225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1197_3_lut_3_lut (.I0(n1778), .I1(n5887), .I2(n1764), 
            .I3(GND_net), .O(n1872));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1197_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_3 (.CI(n28692), .I0(n3158), .I1(GND_net), 
            .CO(n28693));
    SB_CARRY rem_4_add_2122_2 (.CI(VCC_net), .I0(n3258), .I1(VCC_net), 
            .CO(n28692));
    SB_LUT4 div_46_i1187_3_lut_3_lut (.I0(n1778), .I1(n5877), .I2(n1754), 
            .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1187_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1195_3_lut_3_lut (.I0(n1778), .I1(n5885), .I2(n1762), 
            .I3(GND_net), .O(n1870));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1195_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1198_3_lut_3_lut (.I0(n1778), .I1(n5888), .I2(n1765), 
            .I3(GND_net), .O(n1873));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1198_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1192_3_lut_3_lut (.I0(n1778), .I1(n5882), .I2(n1759), 
            .I3(GND_net), .O(n1867));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1192_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1191_3_lut_3_lut (.I0(n1778), .I1(n5881), .I2(n1758), 
            .I3(GND_net), .O(n1866));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1191_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1194_3_lut_3_lut (.I0(n1778), .I1(n5884), .I2(n1761), 
            .I3(GND_net), .O(n1869));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1194_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1519_10_lut (.I0(GND_net), .I1(n2251), .I2(VCC_net), 
            .I3(n28984), .O(n2318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12594_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n13195), .I3(GND_net), .O(n17276));   // verilog/coms.v(126[12] 289[6])
    defparam i12594_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_10 (.CI(n28984), .I0(n2251), .I1(VCC_net), 
            .CO(n28985));
    SB_LUT4 rem_4_add_1519_9_lut (.I0(GND_net), .I1(n2252), .I2(VCC_net), 
            .I3(n28983), .O(n2319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_9 (.CI(n28983), .I0(n2252), .I1(VCC_net), 
            .CO(n28984));
    SB_LUT4 div_46_i1199_3_lut_3_lut (.I0(n1778), .I1(n5889), .I2(n659), 
            .I3(GND_net), .O(n1874));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1199_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1193_3_lut_3_lut (.I0(n1778), .I1(n5883), .I2(n1760), 
            .I3(GND_net), .O(n1868));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1193_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1189_3_lut_3_lut (.I0(n1778), .I1(n5879), .I2(n1756), 
            .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1189_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1519_8_lut (.I0(GND_net), .I1(n2253), .I2(VCC_net), 
            .I3(n28982), .O(n2320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_8 (.CI(n28982), .I0(n2253), .I1(VCC_net), 
            .CO(n28983));
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_add_1519_7_lut (.I0(GND_net), .I1(n2254), .I2(GND_net), 
            .I3(n28981), .O(n2321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1629 (.I0(bit_ctr[26]), .I1(n40187), .I2(n4385), 
            .I3(GND_net), .O(n33361));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1629.LUT_INIT = 16'hacac;
    SB_LUT4 i12229_4_lut (.I0(n26602), .I1(r_Clock_Count_adj_5054[1]), .I2(n320), 
            .I3(r_SM_Main_adj_5053[2]), .O(n16911));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12229_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_i1196_3_lut_3_lut (.I0(n1778), .I1(n5886), .I2(n1763), 
            .I3(GND_net), .O(n1871));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1196_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12233_4_lut (.I0(n16772), .I1(r_Bit_Index_adj_5055[2]), .I2(n4613), 
            .I3(n16641), .O(n16915));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12233_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_46_i1190_3_lut_3_lut (.I0(n1778), .I1(n5880), .I2(n1757), 
            .I3(GND_net), .O(n1865));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1190_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1188_3_lut_3_lut (.I0(n1778), .I1(n5878), .I2(n1755), 
            .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1188_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1519_7 (.CI(n28981), .I0(n2254), .I1(GND_net), 
            .CO(n28982));
    SB_LUT4 div_46_i1270_3_lut_3_lut (.I0(n1886), .I1(n5904), .I2(n1874), 
            .I3(GND_net), .O(n1979));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1270_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12595_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n13195), .I3(GND_net), .O(n17277));   // verilog/coms.v(126[12] 289[6])
    defparam i12595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1259_3_lut_3_lut (.I0(n1886), .I1(n5893), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_559_24_lut (.I0(duty[22]), .I1(n43079), .I2(n3), .I3(n28132), 
            .O(pwm_setpoint_22__N_57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_i1261_3_lut_3_lut (.I0(n1886), .I1(n5895), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1519_6_lut (.I0(GND_net), .I1(n2255), .I2(GND_net), 
            .I3(n28980), .O(n2322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_6 (.CI(n28980), .I0(n2255), .I1(GND_net), 
            .CO(n28981));
    SB_LUT4 rem_4_add_1519_5_lut (.I0(GND_net), .I1(n2256), .I2(VCC_net), 
            .I3(n28979), .O(n2323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_23_lut (.I0(duty[21]), .I1(n43079), .I2(n4_adj_4326), 
            .I3(n28131), .O(pwm_setpoint_22__N_57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1519_5 (.CI(n28979), .I0(n2256), .I1(VCC_net), 
            .CO(n28980));
    SB_CARRY add_559_23 (.CI(n28131), .I0(n43079), .I1(n4_adj_4326), .CO(n28132));
    SB_LUT4 rem_4_add_1519_4_lut (.I0(GND_net), .I1(n2257), .I2(VCC_net), 
            .I3(n28978), .O(n2324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_4 (.CI(n28978), .I0(n2257), .I1(VCC_net), 
            .CO(n28979));
    SB_LUT4 rem_4_add_1519_3_lut (.I0(GND_net), .I1(n2258), .I2(GND_net), 
            .I3(n28977), .O(n2325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_3 (.CI(n28977), .I0(n2258), .I1(GND_net), 
            .CO(n28978));
    SB_CARRY rem_4_add_1519_2 (.CI(VCC_net), .I0(n2358_adj_4622), .I1(VCC_net), 
            .CO(n28977));
    SB_LUT4 div_46_i1260_3_lut_3_lut (.I0(n1886), .I1(n5894), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1258_3_lut_3_lut (.I0(n1886), .I1(n5892), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1586_22_lut (.I0(n2372_adj_4620), .I1(n2339), .I2(VCC_net), 
            .I3(n28976), .O(n2438)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_559_22_lut (.I0(duty[20]), .I1(n43079), .I2(n5_adj_4327), 
            .I3(n28130), .O(pwm_setpoint_22__N_57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_i1269_3_lut_3_lut (.I0(n1886), .I1(n5903), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_559_22 (.CI(n28130), .I0(n43079), .I1(n5_adj_4327), .CO(n28131));
    SB_LUT4 rem_4_add_1586_21_lut (.I0(GND_net), .I1(n2340), .I2(VCC_net), 
            .I3(n28975), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_21_lut (.I0(duty[19]), .I1(n43079), .I2(n6_adj_4328), 
            .I3(n28129), .O(pwm_setpoint_22__N_57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_559_21 (.CI(n28129), .I0(n43079), .I1(n6_adj_4328), .CO(n28130));
    SB_CARRY rem_4_add_1586_21 (.CI(n28975), .I0(n2340), .I1(VCC_net), 
            .CO(n28976));
    SB_LUT4 rem_4_add_1586_20_lut (.I0(GND_net), .I1(n2341), .I2(VCC_net), 
            .I3(n28974), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_20 (.CI(n28974), .I0(n2341), .I1(VCC_net), 
            .CO(n28975));
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n28218), .I0(displacement_23__N_229[17]), 
            .I1(n8_adj_4369), .CO(n28219));
    SB_LUT4 rem_4_add_1586_19_lut (.I0(GND_net), .I1(n2342), .I2(VCC_net), 
            .I3(n28973), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_19 (.CI(n28973), .I0(n2342), .I1(VCC_net), 
            .CO(n28974));
    SB_LUT4 rem_4_add_1586_18_lut (.I0(GND_net), .I1(n2343), .I2(VCC_net), 
            .I3(n28972), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1268_3_lut_3_lut (.I0(n1886), .I1(n5902), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1267_3_lut_3_lut (.I0(n1886), .I1(n5901), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1586_18 (.CI(n28972), .I0(n2343), .I1(VCC_net), 
            .CO(n28973));
    SB_LUT4 rem_4_add_1586_17_lut (.I0(GND_net), .I1(n2344), .I2(VCC_net), 
            .I3(n28971), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_17 (.CI(n28971), .I0(n2344), .I1(VCC_net), 
            .CO(n28972));
    SB_LUT4 rem_4_add_1586_16_lut (.I0(GND_net), .I1(n2345), .I2(VCC_net), 
            .I3(n28970), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_16 (.CI(n28970), .I0(n2345), .I1(VCC_net), 
            .CO(n28971));
    SB_LUT4 rem_4_add_1586_15_lut (.I0(GND_net), .I1(n2346), .I2(VCC_net), 
            .I3(n28969), .O(n2413)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12236_4_lut (.I0(n16772), .I1(r_Bit_Index_adj_5055[1]), .I2(r_Bit_Index_adj_5055[0]), 
            .I3(n16641), .O(n16918));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12236_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_46_i1265_3_lut_3_lut (.I0(n1886), .I1(n5899), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1586_15 (.CI(n28969), .I0(n2346), .I1(VCC_net), 
            .CO(n28970));
    SB_LUT4 rem_4_add_1586_14_lut (.I0(GND_net), .I1(n2347), .I2(VCC_net), 
            .I3(n28968), .O(n2414)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_14 (.CI(n28968), .I0(n2347), .I1(VCC_net), 
            .CO(n28969));
    SB_LUT4 rem_4_add_1586_13_lut (.I0(GND_net), .I1(n2348), .I2(VCC_net), 
            .I3(n28967), .O(n2415)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_13 (.CI(n28967), .I0(n2348), .I1(VCC_net), 
            .CO(n28968));
    SB_LUT4 rem_4_add_1586_12_lut (.I0(GND_net), .I1(n2349), .I2(VCC_net), 
            .I3(n28966), .O(n2416)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_3_lut (.I0(GND_net), .I1(n2958_adj_4426), .I2(GND_net), 
            .I3(n28770), .O(n3025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_12 (.CI(n28966), .I0(n2349), .I1(VCC_net), 
            .CO(n28967));
    SB_CARRY rem_4_add_1988_4 (.CI(n28771), .I0(n2957_adj_4427), .I1(VCC_net), 
            .CO(n28772));
    SB_LUT4 rem_4_add_1988_4_lut (.I0(GND_net), .I1(n2957_adj_4427), .I2(VCC_net), 
            .I3(n28771), .O(n3024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_5 (.CI(n28772), .I0(n2956_adj_4428), .I1(VCC_net), 
            .CO(n28773));
    SB_LUT4 rem_4_add_1586_11_lut (.I0(GND_net), .I1(n2350), .I2(VCC_net), 
            .I3(n28965), .O(n2417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_11 (.CI(n28965), .I0(n2350), .I1(VCC_net), 
            .CO(n28966));
    SB_LUT4 rem_4_add_1988_5_lut (.I0(GND_net), .I1(n2956_adj_4428), .I2(VCC_net), 
            .I3(n28772), .O(n3023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_10_lut (.I0(GND_net), .I1(n2351), .I2(VCC_net), 
            .I3(n28964), .O(n2418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_10 (.CI(n28964), .I0(n2351), .I1(VCC_net), 
            .CO(n28965));
    SB_LUT4 rem_4_add_1586_9_lut (.I0(GND_net), .I1(n2352), .I2(VCC_net), 
            .I3(n28963), .O(n2419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_71_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[16]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_106[16]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1266_3_lut_3_lut (.I0(n1886), .I1(n5900), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1586_9 (.CI(n28963), .I0(n2352), .I1(VCC_net), 
            .CO(n28964));
    SB_LUT4 rem_4_add_1586_8_lut (.I0(GND_net), .I1(n2353), .I2(VCC_net), 
            .I3(n28962), .O(n2420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_20_lut (.I0(duty[18]), .I1(n43079), .I2(n7), .I3(n28128), 
            .O(pwm_setpoint_22__N_57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1988_6 (.CI(n28773), .I0(n2955_adj_4429), .I1(GND_net), 
            .CO(n28774));
    SB_LUT4 rem_4_add_1988_6_lut (.I0(GND_net), .I1(n2955_adj_4429), .I2(GND_net), 
            .I3(n28773), .O(n3022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_8 (.CI(n28962), .I0(n2353), .I1(VCC_net), 
            .CO(n28963));
    SB_LUT4 rem_4_add_1586_7_lut (.I0(GND_net), .I1(n2354), .I2(GND_net), 
            .I3(n28961), .O(n2421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12360_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n37092), .I3(GND_net), .O(n17042));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12360_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12804_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[6] [0]), 
            .I2(n36885), .I3(GND_net), .O(n17486));   // verilog/coms.v(126[12] 289[6])
    defparam i12804_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12803_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[7] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17485));   // verilog/coms.v(126[12] 289[6])
    defparam i12803_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12802_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[7] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17484));   // verilog/coms.v(126[12] 289[6])
    defparam i12802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12801_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[7] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17483));   // verilog/coms.v(126[12] 289[6])
    defparam i12801_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12800_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[7] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17482));   // verilog/coms.v(126[12] 289[6])
    defparam i12800_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12799_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[7] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17481));   // verilog/coms.v(126[12] 289[6])
    defparam i12799_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12798_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[7] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17480));   // verilog/coms.v(126[12] 289[6])
    defparam i12798_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12797_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[7] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17479));   // verilog/coms.v(126[12] 289[6])
    defparam i12797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12812_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[5] [0]), 
            .I2(n36885), .I3(GND_net), .O(n17494));   // verilog/coms.v(126[12] 289[6])
    defparam i12812_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12811_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[6] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17493));   // verilog/coms.v(126[12] 289[6])
    defparam i12811_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12822_3_lut (.I0(encoder0_position[3]), .I1(n2961), .I2(count_enable), 
            .I3(GND_net), .O(n17504));   // quad.v(35[10] 41[6])
    defparam i12822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12821_3_lut (.I0(encoder0_position[2]), .I1(n2962), .I2(count_enable), 
            .I3(GND_net), .O(n17503));   // quad.v(35[10] 41[6])
    defparam i12821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12820_3_lut (.I0(encoder0_position[1]), .I1(n2963), .I2(count_enable), 
            .I3(GND_net), .O(n17502));   // quad.v(35[10] 41[6])
    defparam i12820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1264_3_lut_3_lut (.I0(n1886), .I1(n5898), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12824_3_lut (.I0(encoder0_position[5]), .I1(n2959), .I2(count_enable), 
            .I3(GND_net), .O(n17506));   // quad.v(35[10] 41[6])
    defparam i12824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12361_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n37092), .I3(GND_net), .O(n17043));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12361_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12823_3_lut (.I0(encoder0_position[4]), .I1(n2960), .I2(count_enable), 
            .I3(GND_net), .O(n17505));   // quad.v(35[10] 41[6])
    defparam i12823_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1586_7 (.CI(n28961), .I0(n2354), .I1(GND_net), 
            .CO(n28962));
    SB_LUT4 rem_4_add_1586_6_lut (.I0(GND_net), .I1(n2355), .I2(GND_net), 
            .I3(n28960), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_6 (.CI(n28960), .I0(n2355), .I1(GND_net), 
            .CO(n28961));
    SB_LUT4 div_46_i1271_3_lut_3_lut (.I0(n1886), .I1(n5905), .I2(n660), 
            .I3(GND_net), .O(n1980));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1271_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12362_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n37092), .I3(GND_net), .O(n17044));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12362_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1263_3_lut_3_lut (.I0(n1886), .I1(n5897), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_229[16]), 
            .I2(n9_adj_4366), .I3(n28217), .O(displacement_23__N_80[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_20 (.CI(n28128), .I0(n43079), .I1(n7), .CO(n28129));
    SB_LUT4 rem_4_add_1586_5_lut (.I0(GND_net), .I1(n2356), .I2(VCC_net), 
            .I3(n28959), .O(n2423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_5 (.CI(n28959), .I0(n2356), .I1(VCC_net), 
            .CO(n28960));
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n28217), .I0(displacement_23__N_229[16]), 
            .I1(n9_adj_4366), .CO(n28218));
    SB_LUT4 rem_4_add_1586_4_lut (.I0(GND_net), .I1(n2357_adj_4623), .I2(VCC_net), 
            .I3(n28958), .O(n2424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_19_lut (.I0(duty[17]), .I1(n43079), .I2(n8_adj_4329), 
            .I3(n28127), .O(pwm_setpoint_22__N_57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12363_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n37092), .I3(GND_net), .O(n17045));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12826_3_lut (.I0(encoder0_position[7]), .I1(n2957), .I2(count_enable), 
            .I3(GND_net), .O(n17508));   // quad.v(35[10] 41[6])
    defparam i12826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12825_3_lut (.I0(encoder0_position[6]), .I1(n2958), .I2(count_enable), 
            .I3(GND_net), .O(n17507));   // quad.v(35[10] 41[6])
    defparam i12825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12364_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n37092), .I3(GND_net), .O(n17046));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12364_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12365_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n37092), .I3(GND_net), .O(n17047));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12828_3_lut (.I0(encoder0_position[9]), .I1(n2955), .I2(count_enable), 
            .I3(GND_net), .O(n17510));   // quad.v(35[10] 41[6])
    defparam i12828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12827_3_lut (.I0(encoder0_position[8]), .I1(n2956), .I2(count_enable), 
            .I3(GND_net), .O(n17509));   // quad.v(35[10] 41[6])
    defparam i12827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12366_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n37092), .I3(GND_net), .O(n17048));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12367_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n37092), .I3(GND_net), .O(n17049));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12367_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12830_3_lut (.I0(encoder0_position[11]), .I1(n2953), .I2(count_enable), 
            .I3(GND_net), .O(n17512));   // quad.v(35[10] 41[6])
    defparam i12830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1262_3_lut_3_lut (.I0(n1886), .I1(n5896), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12368_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n37092), .I3(GND_net), .O(n17050));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12368_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1586_4 (.CI(n28958), .I0(n2357_adj_4623), .I1(VCC_net), 
            .CO(n28959));
    SB_LUT4 i12829_3_lut (.I0(encoder0_position[10]), .I1(n2954), .I2(count_enable), 
            .I3(GND_net), .O(n17511));   // quad.v(35[10] 41[6])
    defparam i12829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12832_3_lut (.I0(encoder0_position[13]), .I1(n2951), .I2(count_enable), 
            .I3(GND_net), .O(n17514));   // quad.v(35[10] 41[6])
    defparam i12832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12831_3_lut (.I0(encoder0_position[12]), .I1(n2952), .I2(count_enable), 
            .I3(GND_net), .O(n17513));   // quad.v(35[10] 41[6])
    defparam i12831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_229[15]), 
            .I2(n10_adj_4365), .I3(n28216), .O(displacement_23__N_80[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_3_lut (.I0(GND_net), .I1(n2358_adj_4622), .I2(GND_net), 
            .I3(n28957), .O(n2425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12369_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n37092), .I3(GND_net), .O(n17051));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12370_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n37092), .I3(GND_net), .O(n17052));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12370_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n28216), .I0(displacement_23__N_229[15]), 
            .I1(n10_adj_4365), .CO(n28217));
    SB_CARRY rem_4_add_1586_3 (.CI(n28957), .I0(n2358_adj_4622), .I1(GND_net), 
            .CO(n28958));
    SB_CARRY rem_4_add_1586_2 (.CI(VCC_net), .I0(n2458_adj_4560), .I1(VCC_net), 
            .CO(n28957));
    SB_CARRY add_559_19 (.CI(n28127), .I0(n43079), .I1(n8_adj_4329), .CO(n28128));
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_80[22]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 i12371_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n37092), .I3(GND_net), .O(n17053));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12371_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1340_3_lut_3_lut (.I0(n1991), .I1(n5921), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1653_23_lut (.I0(n2438), .I1(n2438), .I2(n2471_adj_4558), 
            .I3(n28956), .O(n2537_adj_4557)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_229[14]), 
            .I2(n11_adj_4364), .I3(n28215), .O(displacement_23__N_80[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_18_lut (.I0(duty[16]), .I1(n43079), .I2(n9), .I3(n28126), 
            .O(pwm_setpoint_22__N_57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_559_18 (.CI(n28126), .I0(n43079), .I1(n9), .CO(n28127));
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n28215), .I0(displacement_23__N_229[14]), 
            .I1(n11_adj_4364), .CO(n28216));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_229[13]), 
            .I2(n12_adj_4395), .I3(n28214), .O(displacement_23__N_80[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_17_lut (.I0(duty[15]), .I1(n43079), .I2(n10_adj_4330), 
            .I3(n28125), .O(pwm_setpoint_22__N_57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_17_lut.LUT_INIT = 16'h8BB8;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_80[21]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_80[20]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_80[19]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_80[18]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_80[17]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_80[16]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n28214), .I0(displacement_23__N_229[13]), 
            .I1(n12_adj_4395), .CO(n28215));
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_80[15]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_80[14]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_80[13]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_80[12]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_80[11]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_80[10]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 mux_71_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[17]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_80[9]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_80[8]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_80[7]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_80[6]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_80[5]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_LUT4 mux_70_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_106[17]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_80[4]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_80[3]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_80[2]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_80[1]));   // verilog/TinyFPGA_B.v(249[10] 251[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[22]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[21]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[20]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 div_46_i1332_3_lut_3_lut (.I0(n1991), .I1(n5913), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[19]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[18]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 i12372_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n37092), .I3(GND_net), .O(n17054));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12372_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[17]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[16]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[15]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[14]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[13]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[12]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[11]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[10]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[9]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[8]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[7]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[6]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[5]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[4]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[3]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_CARRY add_559_17 (.CI(n28125), .I0(n43079), .I1(n10_adj_4330), 
            .CO(n28126));
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[2]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_LUT4 add_559_16_lut (.I0(duty[14]), .I1(n43079), .I2(n11), .I3(n28124), 
            .O(pwm_setpoint_22__N_57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_16_lut.LUT_INIT = 16'h8BB8;
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[1]));   // verilog/TinyFPGA_B.v(161[10] 174[6])
    SB_DFF communication_counter_1176__i0 (.Q(communication_counter[0]), .C(LED_c), 
           .D(n165));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_CARRY add_559_16 (.CI(n28124), .I0(n43079), .I1(n11), .CO(n28125));
    SB_LUT4 i22_3_lut_adj_1630 (.I0(bit_ctr[2]), .I1(n40194), .I2(n4385), 
            .I3(GND_net), .O(n33375));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1630.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1631 (.I0(bit_ctr[1]), .I1(n40193), .I2(n4385), 
            .I3(GND_net), .O(n33373));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1631.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_229[12]), 
            .I2(n13_adj_4396), .I3(n28213), .O(displacement_23__N_80[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n28213), .I0(displacement_23__N_229[12]), 
            .I1(n13_adj_4396), .CO(n28214));
    SB_LUT4 add_559_15_lut (.I0(duty[13]), .I1(n43079), .I2(n12), .I3(n28123), 
            .O(pwm_setpoint_22__N_57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_229[11]), 
            .I2(n14_adj_4397), .I3(n28212), .O(displacement_23__N_80[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n28212), .I0(displacement_23__N_229[11]), 
            .I1(n14_adj_4397), .CO(n28213));
    SB_LUT4 i12836_3_lut (.I0(encoder0_position[17]), .I1(n2947), .I2(count_enable), 
            .I3(GND_net), .O(n17518));   // quad.v(35[10] 41[6])
    defparam i12836_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_559_15 (.CI(n28123), .I0(n43079), .I1(n12), .CO(n28124));
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_229[10]), 
            .I2(n15_adj_4398), .I3(n28211), .O(displacement_23__N_80[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12835_3_lut (.I0(encoder0_position[16]), .I1(n2948), .I2(count_enable), 
            .I3(GND_net), .O(n17517));   // quad.v(35[10] 41[6])
    defparam i12835_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n28211), .I0(displacement_23__N_229[10]), 
            .I1(n15_adj_4398), .CO(n28212));
    SB_LUT4 div_46_i1331_3_lut_3_lut (.I0(n1991), .I1(n5912), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12834_3_lut (.I0(encoder0_position[15]), .I1(n2949), .I2(count_enable), 
            .I3(GND_net), .O(n17516));   // quad.v(35[10] 41[6])
    defparam i12834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12833_3_lut (.I0(encoder0_position[14]), .I1(n2950), .I2(count_enable), 
            .I3(GND_net), .O(n17515));   // quad.v(35[10] 41[6])
    defparam i12833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_22_lut (.I0(n2439), .I1(n2439), .I2(n2471_adj_4558), 
            .I3(n28955), .O(n2538_adj_4556)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_559_14_lut (.I0(duty[12]), .I1(n43079), .I2(n13_adj_4331), 
            .I3(n28122), .O(pwm_setpoint_22__N_57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_229[9]), 
            .I2(n16_adj_4399), .I3(n28210), .O(displacement_23__N_80[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n28210), .I0(displacement_23__N_229[9]), 
            .I1(n16_adj_4399), .CO(n28211));
    SB_LUT4 div_46_i1330_3_lut_3_lut (.I0(n1991), .I1(n5911), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_229[8]), 
            .I2(n17_adj_4400), .I3(n28209), .O(displacement_23__N_80[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n28209), .I0(displacement_23__N_229[8]), 
            .I1(n17_adj_4400), .CO(n28210));
    SB_CARRY add_559_14 (.CI(n28122), .I0(n43079), .I1(n13_adj_4331), 
            .CO(n28123));
    SB_LUT4 add_559_13_lut (.I0(duty[11]), .I1(n43079), .I2(n14), .I3(n28121), 
            .O(pwm_setpoint_22__N_57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_229[7]), 
            .I2(n18_adj_4401), .I3(n28208), .O(displacement_23__N_80[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1329_3_lut_3_lut (.I0(n1991), .I1(n5910), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1328_3_lut_3_lut (.I0(n1991), .I1(n5909), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1327_3_lut_3_lut (.I0(n1991), .I1(n5908), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12847_3_lut (.I0(encoder1_position[4]), .I1(n2910), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17529));   // quad.v(35[10] 41[6])
    defparam i12847_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_22 (.CI(n28955), .I0(n2439), .I1(n2471_adj_4558), 
            .CO(n28956));
    SB_CARRY add_559_13 (.CI(n28121), .I0(n43079), .I1(n14), .CO(n28122));
    SB_LUT4 i12846_3_lut (.I0(encoder1_position[3]), .I1(n2911), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17528));   // quad.v(35[10] 41[6])
    defparam i12846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12845_3_lut (.I0(encoder1_position[2]), .I1(n2912), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17527));   // quad.v(35[10] 41[6])
    defparam i12845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_21_lut (.I0(n2440), .I1(n2440), .I2(n2471_adj_4558), 
            .I3(n28954), .O(n2539_adj_4555)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_21_lut.LUT_INIT = 16'hCA3A;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_i1338_3_lut_3_lut (.I0(n1991), .I1(n5919), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12844_3_lut (.I0(encoder1_position[1]), .I1(n2913), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17526));   // quad.v(35[10] 41[6])
    defparam i12844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1339_3_lut_3_lut (.I0(n1991), .I1(n5920), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1176_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[31]), .I3(n28650), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_12_lut (.I0(duty[10]), .I1(n43079), .I2(n15_adj_4332), 
            .I3(n28120), .O(pwm_setpoint_22__N_57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1653_21 (.CI(n28954), .I0(n2440), .I1(n2471_adj_4558), 
            .CO(n28955));
    SB_LUT4 communication_counter_1176_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[30]), .I3(n28649), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_20_lut (.I0(n2441), .I1(n2441), .I2(n2471_adj_4558), 
            .I3(n28953), .O(n2540_adj_4554)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n28208), .I0(displacement_23__N_229[7]), 
            .I1(n18_adj_4401), .CO(n28209));
    SB_CARRY add_559_12 (.CI(n28120), .I0(n43079), .I1(n15_adj_4332), 
            .CO(n28121));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_229[6]), 
            .I2(n19_adj_4402), .I3(n28207), .O(displacement_23__N_80[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1337_3_lut_3_lut (.I0(n1991), .I1(n5918), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1176_add_4_32 (.CI(n28649), .I0(GND_net), 
            .I1(communication_counter[30]), .CO(n28650));
    SB_LUT4 add_559_11_lut (.I0(duty[9]), .I1(n43079), .I2(n16), .I3(n28119), 
            .O(pwm_setpoint_22__N_57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n28207), .I0(displacement_23__N_229[6]), 
            .I1(n19_adj_4402), .CO(n28208));
    SB_LUT4 communication_counter_1176_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[29]), .I3(n28648), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_31 (.CI(n28648), .I0(GND_net), 
            .I1(communication_counter[29]), .CO(n28649));
    SB_CARRY add_559_11 (.CI(n28119), .I0(n43079), .I1(n16), .CO(n28120));
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_229[5]), 
            .I2(n20_adj_4403), .I3(n28206), .O(displacement_23__N_80[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_10_lut (.I0(duty[8]), .I1(n43079), .I2(n17_adj_4333), 
            .I3(n28118), .O(pwm_setpoint_22__N_57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n28206), .I0(displacement_23__N_229[5]), 
            .I1(n20_adj_4403), .CO(n28207));
    SB_LUT4 communication_counter_1176_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[28]), .I3(n28647), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_30 (.CI(n28647), .I0(GND_net), 
            .I1(communication_counter[28]), .CO(n28648));
    SB_LUT4 communication_counter_1176_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[27]), .I3(n28646), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_29 (.CI(n28646), .I0(GND_net), 
            .I1(communication_counter[27]), .CO(n28647));
    SB_LUT4 div_46_i1335_3_lut_3_lut (.I0(n1991), .I1(n5916), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1176_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[26]), .I3(n28645), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_229[4]), 
            .I2(n21_adj_4404), .I3(n28205), .O(displacement_23__N_80[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1336_3_lut_3_lut (.I0(n1991), .I1(n5917), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n28205), .I0(displacement_23__N_229[4]), 
            .I1(n21_adj_4404), .CO(n28206));
    SB_CARRY add_559_10 (.CI(n28118), .I0(n43079), .I1(n17_adj_4333), 
            .CO(n28119));
    SB_LUT4 div_46_i1334_3_lut_3_lut (.I0(n1991), .I1(n5915), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1176_add_4_28 (.CI(n28645), .I0(GND_net), 
            .I1(communication_counter[26]), .CO(n28646));
    SB_LUT4 div_46_i1341_3_lut_3_lut (.I0(n1991), .I1(n5922), .I2(n661), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1176_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[25]), .I3(n28644), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1333_3_lut_3_lut (.I0(n1991), .I1(n5914), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_559_9_lut (.I0(duty[7]), .I1(n43079), .I2(n18_adj_4334), 
            .I3(n28117), .O(pwm_setpoint_22__N_57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i25_4_lut (.I0(n24867), .I1(n35361), .I2(state[0]), .I3(n15464), 
            .O(n11_adj_4921));   // verilog/neopixel.v(35[12] 117[6])
    defparam i25_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 div_46_i1407_3_lut_3_lut (.I0(n2093), .I1(n5938), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1991_3_lut (.I0(n2934), .I1(n3001), .I2(n2966), .I3(GND_net), 
            .O(n3033));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2010_3_lut (.I0(n2953_adj_4431), .I1(n3020), .I2(n2966), 
            .I3(GND_net), .O(n3052));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2005_3_lut (.I0(n2948_adj_4436), .I1(n3015), .I2(n2966), 
            .I3(GND_net), .O(n3047));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2009_3_lut (.I0(n2952_adj_4432), .I1(n3019), .I2(n2966), 
            .I3(GND_net), .O(n3051));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2003_3_lut (.I0(n2946_adj_4438), .I1(n3013), .I2(n2966), 
            .I3(GND_net), .O(n3045));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2008_3_lut (.I0(n2951_adj_4433), .I1(n3018), .I2(n2966), 
            .I3(GND_net), .O(n3050));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2006_3_lut (.I0(n2949_adj_4435), .I1(n3016), .I2(n2966), 
            .I3(GND_net), .O(n3048));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2004_3_lut (.I0(n2947_adj_4437), .I1(n3014), .I2(n2966), 
            .I3(GND_net), .O(n3046));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1403_3_lut_3_lut (.I0(n2093), .I1(n5934), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1402_3_lut_3_lut (.I0(n2093), .I1(n5933), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_229[3]), 
            .I2(n22_adj_4405), .I3(n28204), .O(displacement_23__N_80[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_27 (.CI(n28644), .I0(GND_net), 
            .I1(communication_counter[25]), .CO(n28645));
    SB_LUT4 communication_counter_1176_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[24]), .I3(n28643), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1397_3_lut_3_lut (.I0(n2093), .I1(n5928), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1396_3_lut_3_lut (.I0(n2093), .I1(n5927), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1176_add_4_26 (.CI(n28643), .I0(GND_net), 
            .I1(communication_counter[24]), .CO(n28644));
    SB_LUT4 div_46_i1395_3_lut_3_lut (.I0(n2093), .I1(n5926), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n28204), .I0(displacement_23__N_229[3]), 
            .I1(n22_adj_4405), .CO(n28205));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_229[2]), 
            .I2(n23_adj_4406), .I3(n28203), .O(displacement_23__N_80[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1398_3_lut_3_lut (.I0(n2093), .I1(n5929), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n28203), .I0(displacement_23__N_229[2]), 
            .I1(n23_adj_4406), .CO(n28204));
    SB_LUT4 div_46_i1394_3_lut_3_lut (.I0(n2093), .I1(n5925), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_559_9 (.CI(n28117), .I0(n43079), .I1(n18_adj_4334), .CO(n28118));
    SB_LUT4 communication_counter_1176_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[23]), .I3(n28642), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1405_3_lut_3_lut (.I0(n2093), .I1(n5936), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1176_add_4_25 (.CI(n28642), .I0(GND_net), 
            .I1(communication_counter[23]), .CO(n28643));
    SB_LUT4 communication_counter_1176_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[22]), .I3(n28641), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_71_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[18]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_106[18]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1406_3_lut_3_lut (.I0(n2093), .I1(n5937), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1176_add_4_24 (.CI(n28641), .I0(GND_net), 
            .I1(communication_counter[22]), .CO(n28642));
    SB_LUT4 div_46_i1404_3_lut_3_lut (.I0(n2093), .I1(n5935), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1176_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[21]), .I3(n28640), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1632 (.I0(\FRAME_MATCHER.state_31__N_2426 [2]), .I1(n7_adj_4477), 
            .I2(\FRAME_MATCHER.i_31__N_2390 ), .I3(n2855), .O(n6_adj_4389));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1632.LUT_INIT = 16'hfcec;
    SB_LUT4 i3_4_lut_adj_1633 (.I0(\FRAME_MATCHER.i_31__N_2386 ), .I1(n6_adj_4389), 
            .I2(n8849), .I3(n122), .O(n8_adj_4923));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_1633.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1634 (.I0(\FRAME_MATCHER.state_31__N_2426 [2]), .I1(n8_adj_4923), 
            .I2(n63), .I3(n4_adj_5006), .O(n43272));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1634.LUT_INIT = 16'hefcf;
    SB_CARRY rem_4_add_1653_20 (.CI(n28953), .I0(n2441), .I1(n2471_adj_4558), 
            .CO(n28954));
    SB_CARRY communication_counter_1176_add_4_23 (.CI(n28640), .I0(GND_net), 
            .I1(communication_counter[21]), .CO(n28641));
    SB_LUT4 i12842_3_lut (.I0(encoder0_position[23]), .I1(n2941), .I2(count_enable), 
            .I3(GND_net), .O(n17524));   // quad.v(35[10] 41[6])
    defparam i12842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12841_3_lut (.I0(encoder0_position[22]), .I1(n2942), .I2(count_enable), 
            .I3(GND_net), .O(n17523));   // quad.v(35[10] 41[6])
    defparam i12841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12840_3_lut (.I0(encoder0_position[21]), .I1(n2943), .I2(count_enable), 
            .I3(GND_net), .O(n17522));   // quad.v(35[10] 41[6])
    defparam i12840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12839_3_lut (.I0(encoder0_position[20]), .I1(n2944), .I2(count_enable), 
            .I3(GND_net), .O(n17521));   // quad.v(35[10] 41[6])
    defparam i12839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1408_3_lut_3_lut (.I0(n2093), .I1(n5939), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1176_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[20]), .I3(n28639), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12851_3_lut (.I0(encoder1_position[8]), .I1(n2906), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17533));   // quad.v(35[10] 41[6])
    defparam i12851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12850_3_lut (.I0(encoder1_position[7]), .I1(n2907), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17532));   // quad.v(35[10] 41[6])
    defparam i12850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12849_3_lut (.I0(encoder1_position[6]), .I1(n2908), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17531));   // quad.v(35[10] 41[6])
    defparam i12849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12848_3_lut (.I0(encoder1_position[5]), .I1(n2909), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17530));   // quad.v(35[10] 41[6])
    defparam i12848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1401_3_lut_3_lut (.I0(n2093), .I1(n5932), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1176_add_4_22 (.CI(n28639), .I0(GND_net), 
            .I1(communication_counter[20]), .CO(n28640));
    SB_LUT4 i12859_3_lut (.I0(encoder1_position[16]), .I1(n2898), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17541));   // quad.v(35[10] 41[6])
    defparam i12859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1176_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[19]), .I3(n28638), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12858_3_lut (.I0(encoder1_position[15]), .I1(n2899), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17540));   // quad.v(35[10] 41[6])
    defparam i12858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12869_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n37155), 
            .I3(GND_net), .O(n17551));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12869_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1399_3_lut_3_lut (.I0(n2093), .I1(n5930), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY communication_counter_1176_add_4_21 (.CI(n28638), .I0(GND_net), 
            .I1(communication_counter[19]), .CO(n28639));
    SB_LUT4 div_46_i1400_3_lut_3_lut (.I0(n2093), .I1(n5931), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1409_3_lut_3_lut (.I0(n2093), .I1(n5940), .I2(n662), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12868_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4379), 
            .I3(n15459), .O(n17550));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12868_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 communication_counter_1176_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[18]), .I3(n28637), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1468_3_lut_3_lut (.I0(n2192), .I1(n5952), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12871_3_lut (.I0(color[1]), .I1(n16695), .I2(n15_adj_4338), 
            .I3(GND_net), .O(n17553));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i12871_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_1176_add_4_20 (.CI(n28637), .I0(GND_net), 
            .I1(communication_counter[18]), .CO(n28638));
    SB_LUT4 div_46_i1459_3_lut_3_lut (.I0(n2192), .I1(n5943), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i24_3_lut_adj_1635 (.I0(n40170), .I1(bit_ctr[17]), .I2(n4385), 
            .I3(GND_net), .O(n33321));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1635.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut_adj_1636 (.I0(n40169), .I1(bit_ctr[16]), .I2(n4385), 
            .I3(GND_net), .O(n33319));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1636.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1469_3_lut_3_lut (.I0(n2192), .I1(n5953), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12879_3_lut (.I0(color[3]), .I1(n16695), .I2(n15_adj_4338), 
            .I3(GND_net), .O(n17561));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i12879_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 communication_counter_1176_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[17]), .I3(n28636), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1465_3_lut_3_lut (.I0(n2192), .I1(n5949), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12878_3_lut (.I0(color[2]), .I1(n16695), .I2(n15_adj_4338), 
            .I3(GND_net), .O(n17560));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i12878_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12810_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[6] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17492));   // verilog/coms.v(126[12] 289[6])
    defparam i12810_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12809_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[6] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17491));   // verilog/coms.v(126[12] 289[6])
    defparam i12809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12808_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[6] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17490));   // verilog/coms.v(126[12] 289[6])
    defparam i12808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1466_3_lut_3_lut (.I0(n2192), .I1(n5950), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1475_3_lut_3_lut (.I0(n2192), .I1(n5959), .I2(n663), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1463_3_lut_3_lut (.I0(n2192), .I1(n5947), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_559_8_lut (.I0(duty[6]), .I1(n43079), .I2(n19_adj_4335), 
            .I3(n28116), .O(pwm_setpoint_22__N_57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12807_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[6] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17489));   // verilog/coms.v(126[12] 289[6])
    defparam i12807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12806_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[6] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17488));   // verilog/coms.v(126[12] 289[6])
    defparam i12806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2011_3_lut (.I0(n2954_adj_4430), .I1(n3021), .I2(n2966), 
            .I3(GND_net), .O(n3053));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2007_3_lut (.I0(n2950_adj_4434), .I1(n3017), .I2(n2966), 
            .I3(GND_net), .O(n3049));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2001_3_lut (.I0(n2944_adj_4440), .I1(n3011), .I2(n2966), 
            .I3(GND_net), .O(n3043));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2000_3_lut (.I0(n2943_adj_4441), .I1(n3010), .I2(n2966), 
            .I3(GND_net), .O(n3042));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1995_3_lut (.I0(n2938), .I1(n3005), .I2(n2966), .I3(GND_net), 
            .O(n3037));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1993_3_lut (.I0(n2936), .I1(n3003), .I2(n2966), .I3(GND_net), 
            .O(n3035));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1994_3_lut (.I0(n2937), .I1(n3004), .I2(n2966), .I3(GND_net), 
            .O(n3036));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1992_3_lut (.I0(n2935), .I1(n3002), .I2(n2966), .I3(GND_net), 
            .O(n3034));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1999_3_lut (.I0(n2942_adj_4442), .I1(n3009), .I2(n2966), 
            .I3(GND_net), .O(n3041));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1997_3_lut (.I0(n2940), .I1(n3007), .I2(n2966), .I3(GND_net), 
            .O(n3039));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1998_3_lut (.I0(n2941_adj_4443), .I1(n3008), .I2(n2966), 
            .I3(GND_net), .O(n3040));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1996_3_lut (.I0(n2939), .I1(n3006), .I2(n2966), .I3(GND_net), 
            .O(n3038));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2013_3_lut (.I0(n2956_adj_4428), .I1(n3023), .I2(n2966), 
            .I3(GND_net), .O(n3055));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2012_3_lut (.I0(n2955_adj_4429), .I1(n3022), .I2(n2966), 
            .I3(GND_net), .O(n3054));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2002_3_lut (.I0(n2945_adj_4439), .I1(n3012), .I2(n2966), 
            .I3(GND_net), .O(n3044));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1462_3_lut_3_lut (.I0(n2192), .I1(n5946), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_559_8 (.CI(n28116), .I0(n43079), .I1(n19_adj_4335), .CO(n28117));
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_229[1]), 
            .I2(n24_adj_4407), .I3(n28202), .O(displacement_23__N_80[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12805_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[6] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17487));   // verilog/coms.v(126[12] 289[6])
    defparam i12805_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY communication_counter_1176_add_4_19 (.CI(n28636), .I0(GND_net), 
            .I1(communication_counter[17]), .CO(n28637));
    SB_LUT4 i12819_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[5] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17501));   // verilog/coms.v(126[12] 289[6])
    defparam i12819_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_559_7_lut (.I0(duty[5]), .I1(n43079), .I2(n20_adj_4336), 
            .I3(n28115), .O(pwm_setpoint_22__N_57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_559_7 (.CI(n28115), .I0(n43079), .I1(n20_adj_4336), .CO(n28116));
    SB_LUT4 rem_4_add_1653_19_lut (.I0(n2442), .I1(n2442), .I2(n2471_adj_4558), 
            .I3(n28952), .O(n2541_adj_4553)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12818_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[5] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17500));   // verilog/coms.v(126[12] 289[6])
    defparam i12818_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1461_3_lut_3_lut (.I0(n2192), .I1(n5945), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12817_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[5] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17499));   // verilog/coms.v(126[12] 289[6])
    defparam i12817_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1464_3_lut_3_lut (.I0(n2192), .I1(n5948), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n28202), .I0(displacement_23__N_229[1]), 
            .I1(n24_adj_4407), .CO(n28203));
    SB_CARRY rem_4_add_1653_19 (.CI(n28952), .I0(n2442), .I1(n2471_adj_4558), 
            .CO(n28953));
    SB_LUT4 rem_4_add_1653_18_lut (.I0(n2443), .I1(n2443), .I2(n2471_adj_4558), 
            .I3(n28951), .O(n2542_adj_4552)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1653_18 (.CI(n28951), .I0(n2443), .I1(n2471_adj_4558), 
            .CO(n28952));
    SB_LUT4 div_46_i1460_3_lut_3_lut (.I0(n2192), .I1(n5944), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12816_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[5] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17498));   // verilog/coms.v(126[12] 289[6])
    defparam i12816_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12815_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[5] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17497));   // verilog/coms.v(126[12] 289[6])
    defparam i12815_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12814_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[5] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17496));   // verilog/coms.v(126[12] 289[6])
    defparam i12814_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1653_17_lut (.I0(n2444), .I1(n2444), .I2(n2471_adj_4558), 
            .I3(n28950), .O(n2543_adj_4551)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_229[0]), 
            .I2(n25_adj_4408), .I3(VCC_net), .O(displacement_23__N_80[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_i1470_3_lut_3_lut (.I0(n2192), .I1(n5954), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2015_3_lut (.I0(n2958_adj_4426), .I1(n3025), .I2(n2966), 
            .I3(GND_net), .O(n3057));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2014_3_lut (.I0(n2957_adj_4427), .I1(n3024), .I2(n2966), 
            .I3(GND_net), .O(n3056));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1637 (.I0(n3056), .I1(n3057), .I2(n3058), .I3(GND_net), 
            .O(n35694));
    defparam i1_3_lut_adj_1637.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut (.I0(n3044), .I1(n3054), .I2(n35694), .I3(n3055), 
            .O(n30_adj_4932));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i14_4_lut (.I0(n3038), .I1(n3040), .I2(n3039), .I3(n3041), 
            .O(n37_adj_4930));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n3034), .I1(n3036), .I2(n3035), .I3(n3037), 
            .O(n36_adj_4931));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37_adj_4930), .I1(n3042), .I2(n30_adj_4932), 
            .I3(n3043), .O(n42_adj_4926));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n3049), .I1(n3053), .I2(n3046), .I3(n3048), 
            .O(n40_adj_4928));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n3052), .I1(n36_adj_4931), .I2(n3033), .I3(n3032), 
            .O(n41_adj_4927));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n3050), .I1(n3045), .I2(n3051), .I3(n3047), 
            .O(n39_adj_4929));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_4929), .I1(n41_adj_4927), .I2(n40_adj_4928), 
            .I3(n42_adj_4926), .O(n3065));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12813_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[5] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17495));   // verilog/coms.v(126[12] 289[6])
    defparam i12813_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12890_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1169), .I3(GND_net), .O(n17572));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i6_3_lut (.I0(communication_counter[5]), .I1(n28_adj_4456), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3058));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_559_6_lut (.I0(duty[4]), .I1(n43079), .I2(n21), .I3(n28114), 
            .O(pwm_setpoint_22__N_57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12888_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1169), .I3(GND_net), .O(n17570));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12887_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1169), .I3(GND_net), .O(n17569));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12886_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1169), .I3(GND_net), .O(n17568));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1471_3_lut_3_lut (.I0(n2192), .I1(n5955), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12885_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1169), .I3(GND_net), .O(n17567));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1473_3_lut_3_lut (.I0(n2192), .I1(n5957), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1472_3_lut_3_lut (.I0(n2192), .I1(n5956), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1474_3_lut_3_lut (.I0(n2192), .I1(n5958), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1467_3_lut_3_lut (.I0(n2192), .I1(n5951), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1528_3_lut_3_lut (.I0(n2288), .I1(n5968), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1522_3_lut_3_lut (.I0(n2288), .I1(n5962), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_3_lut_adj_1638 (.I0(n1956), .I1(n1957), .I2(n1958), .I3(GND_net), 
            .O(n35580));
    defparam i1_3_lut_adj_1638.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1639 (.I0(n1947), .I1(n1954), .I2(n35580), .I3(n1955), 
            .O(n15_adj_4936));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut_adj_1639.LUT_INIT = 16'heaaa;
    SB_LUT4 i7_4_lut_adj_1640 (.I0(n1944), .I1(n1945), .I2(n1943), .I3(n1946), 
            .O(n19_adj_4934));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1953), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4935));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n19_adj_4934), .I1(n15_adj_4936), .I2(n1948), 
            .I3(n1949), .O(n22_adj_4933));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1641 (.I0(n1952), .I1(n22_adj_4933), .I2(n18_adj_4935), 
            .I3(n1950), .O(n1976_adj_4689));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i17_3_lut (.I0(communication_counter[16]), .I1(n17_adj_4466), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1958));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut_adj_1642 (.I0(n40168), .I1(bit_ctr[15]), .I2(n4385), 
            .I3(GND_net), .O(n33317));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1642.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1525_3_lut_3_lut (.I0(n2288), .I1(n5965), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1523_3_lut_3_lut (.I0(n2288), .I1(n5963), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i18_3_lut (.I0(communication_counter[17]), .I1(n16_adj_4467), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i19_3_lut (.I0(communication_counter[18]), .I1(n15_adj_4468), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1758_adj_4498));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1199_3_lut (.I0(n1758_adj_4498), .I1(n1825), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1526_3_lut_3_lut (.I0(n2288), .I1(n5966), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1529_3_lut_3_lut (.I0(n2288), .I1(n5969), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i890_3_lut_3_lut (.I0(n1316), .I1(n5834), .I2(n1299), 
            .I3(GND_net), .O(n1419));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i890_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12898_3_lut (.I0(setpoint[7]), .I1(n4299), .I2(n36839), .I3(GND_net), 
            .O(n17580));   // verilog/coms.v(126[12] 289[6])
    defparam i12898_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_71_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[19]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_46_i1537_3_lut_3_lut (.I0(n2288), .I1(n5977), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_70_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_106[19]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1536_3_lut_3_lut (.I0(n2288), .I1(n5976), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1524_3_lut_3_lut (.I0(n2288), .I1(n5964), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i20_3_lut (.I0(communication_counter[19]), .I1(n14_adj_4469), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1658));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1131_3_lut (.I0(n1658), .I1(n1725), .I2(n1679), .I3(GND_net), 
            .O(n1757_adj_4497));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1198_3_lut (.I0(n1757_adj_4497), .I1(n1824), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[20]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_106[20]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1532_3_lut_3_lut (.I0(n2288), .I1(n5972), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1531_3_lut_3_lut (.I0(n2288), .I1(n5971), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2140_3_lut (.I0(n3147), .I1(n3214), .I2(n3164), .I3(GND_net), 
            .O(n3246));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2145_3_lut (.I0(n3152), .I1(n3219), .I2(n3164), .I3(GND_net), 
            .O(n3251));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2134_3_lut (.I0(n3141), .I1(n3208), .I2(n3164), .I3(GND_net), 
            .O(n3240));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1530_3_lut_3_lut (.I0(n2288), .I1(n5970), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2127_3_lut (.I0(n3134), .I1(n3201), .I2(n3164), .I3(GND_net), 
            .O(n3233));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2126_3_lut (.I0(n3133), .I1(n3200), .I2(n3164), .I3(GND_net), 
            .O(n3232));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2130_3_lut (.I0(n3137), .I1(n3204), .I2(n3164), .I3(GND_net), 
            .O(n3236));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2132_3_lut (.I0(n3139), .I1(n3206), .I2(n3164), .I3(GND_net), 
            .O(n3238));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2138_3_lut (.I0(n3145), .I1(n3212), .I2(n3164), .I3(GND_net), 
            .O(n3244));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2137_3_lut (.I0(n3144), .I1(n3211), .I2(n3164), .I3(GND_net), 
            .O(n3243));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2136_3_lut (.I0(n3143), .I1(n3210), .I2(n3164), .I3(GND_net), 
            .O(n3242));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1935_3_lut (.I0(n2846), .I1(n2913_adj_4445), .I2(n2867), 
            .I3(GND_net), .O(n2945_adj_4439));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1940_3_lut (.I0(n2851), .I1(n2918), .I2(n2867), .I3(GND_net), 
            .O(n2950_adj_4434));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1936_3_lut (.I0(n2847), .I1(n2914_adj_4444), .I2(n2867), 
            .I3(GND_net), .O(n2946_adj_4438));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1938_3_lut (.I0(n2849), .I1(n2916), .I2(n2867), .I3(GND_net), 
            .O(n2948_adj_4436));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1942_3_lut (.I0(n2853), .I1(n2920), .I2(n2867), .I3(GND_net), 
            .O(n2952_adj_4432));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1943_3_lut (.I0(n2854), .I1(n2921), .I2(n2867), .I3(GND_net), 
            .O(n2953_adj_4431));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1937_3_lut (.I0(n2848), .I1(n2915), .I2(n2867), .I3(GND_net), 
            .O(n2947_adj_4437));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1939_3_lut (.I0(n2850), .I1(n2917), .I2(n2867), .I3(GND_net), 
            .O(n2949_adj_4435));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1934_3_lut (.I0(n2845), .I1(n2912_adj_4446), .I2(n2867), 
            .I3(GND_net), .O(n2944_adj_4440));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1941_3_lut (.I0(n2852), .I1(n2919), .I2(n2867), .I3(GND_net), 
            .O(n2951_adj_4433));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1933_3_lut (.I0(n2844), .I1(n2911_adj_4447), .I2(n2867), 
            .I3(GND_net), .O(n2943_adj_4441));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1932_3_lut (.I0(n2843), .I1(n2910_adj_4448), .I2(n2867), 
            .I3(GND_net), .O(n2942_adj_4442));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1930_3_lut (.I0(n2841), .I1(n2908_adj_4450), .I2(n2867), 
            .I3(GND_net), .O(n2940));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1928_3_lut (.I0(n2839), .I1(n2906_adj_4319), .I2(n2867), 
            .I3(GND_net), .O(n2938));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1929_3_lut (.I0(n2840), .I1(n2907_adj_4451), .I2(n2867), 
            .I3(GND_net), .O(n2939));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1927_3_lut (.I0(n2838), .I1(n2905_adj_4470), .I2(n2867), 
            .I3(GND_net), .O(n2937));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2129_3_lut (.I0(n3136), .I1(n3203), .I2(n3164), .I3(GND_net), 
            .O(n3235));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12897_3_lut (.I0(setpoint[6]), .I1(n4298), .I2(n36839), .I3(GND_net), 
            .O(n17579));   // verilog/coms.v(126[12] 289[6])
    defparam i12897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2128_3_lut (.I0(n3135), .I1(n3202), .I2(n3164), .I3(GND_net), 
            .O(n3234));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2144_3_lut (.I0(n3151), .I1(n3218), .I2(n3164), .I3(GND_net), 
            .O(n3250));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1539_3_lut_3_lut (.I0(n2288), .I1(n5979), .I2(n664), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2147_3_lut (.I0(n3154), .I1(n3221), .I2(n3164), .I3(GND_net), 
            .O(n3253));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1945_3_lut (.I0(n2856), .I1(n2923), .I2(n2867), .I3(GND_net), 
            .O(n2955_adj_4429));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1944_3_lut (.I0(n2855_adj_4474), .I1(n2922), .I2(n2867), 
            .I3(GND_net), .O(n2954_adj_4430));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1931_3_lut (.I0(n2842), .I1(n2909_adj_4449), .I2(n2867), 
            .I3(GND_net), .O(n2941_adj_4443));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1947_3_lut (.I0(n2858), .I1(n2925), .I2(n2867), .I3(GND_net), 
            .O(n2957_adj_4427));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1946_3_lut (.I0(n2857), .I1(n2924), .I2(n2867), .I3(GND_net), 
            .O(n2956_adj_4428));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1865_3_lut (.I0(n2744), .I1(n2811), .I2(n2768), .I3(GND_net), 
            .O(n2843));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1863_3_lut (.I0(n2742), .I1(n2809), .I2(n2768), .I3(GND_net), 
            .O(n2841));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1864_3_lut (.I0(n2743), .I1(n2810), .I2(n2768), .I3(GND_net), 
            .O(n2842));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1862_3_lut (.I0(n2741), .I1(n2808), .I2(n2768), .I3(GND_net), 
            .O(n2840));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1867_3_lut (.I0(n2746), .I1(n2813), .I2(n2768), .I3(GND_net), 
            .O(n2845));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1866_3_lut (.I0(n2745), .I1(n2812), .I2(n2768), .I3(GND_net), 
            .O(n2844));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1873_3_lut (.I0(n2752), .I1(n2819), .I2(n2768), .I3(GND_net), 
            .O(n2851));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1874_3_lut (.I0(n2753), .I1(n2820), .I2(n2768), .I3(GND_net), 
            .O(n2852));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1872_3_lut (.I0(n2751), .I1(n2818), .I2(n2768), .I3(GND_net), 
            .O(n2850));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1872_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1875_3_lut (.I0(n2754), .I1(n2821), .I2(n2768), .I3(GND_net), 
            .O(n2853));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1868_3_lut (.I0(n2747), .I1(n2814), .I2(n2768), .I3(GND_net), 
            .O(n2846));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1868_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1869_3_lut (.I0(n2748), .I1(n2815), .I2(n2768), .I3(GND_net), 
            .O(n2847));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1870_3_lut (.I0(n2749), .I1(n2816), .I2(n2768), .I3(GND_net), 
            .O(n2848));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1877_3_lut (.I0(n2756), .I1(n2823), .I2(n2768), .I3(GND_net), 
            .O(n2855_adj_4474));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1871_3_lut (.I0(n2750), .I1(n2817), .I2(n2768), .I3(GND_net), 
            .O(n2849));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1876_3_lut (.I0(n2755), .I1(n2822), .I2(n2768), .I3(GND_net), 
            .O(n2854));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1861_3_lut (.I0(n2740), .I1(n2807), .I2(n2768), .I3(GND_net), 
            .O(n2839));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2142_3_lut (.I0(n3149), .I1(n3216), .I2(n3164), .I3(GND_net), 
            .O(n3248));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2143_3_lut (.I0(n3150), .I1(n3217), .I2(n3164), .I3(GND_net), 
            .O(n3249));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2125_3_lut (.I0(n3132), .I1(n3199), .I2(n3164), .I3(GND_net), 
            .O(n3231));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1527_3_lut_3_lut (.I0(n2288), .I1(n5967), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1860_3_lut (.I0(n2739), .I1(n2806), .I2(n2768), .I3(GND_net), 
            .O(n2838));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1858_3_lut (.I0(n2737), .I1(n2804), .I2(n2768), .I3(GND_net), 
            .O(n2836));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1857_3_lut (.I0(n2736), .I1(n2803), .I2(n2768), .I3(GND_net), 
            .O(n2835));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1798_3_lut (.I0(n2645), .I1(n2712), .I2(n2669), .I3(GND_net), 
            .O(n2744));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1804_3_lut (.I0(n2651), .I1(n2718), .I2(n2669), .I3(GND_net), 
            .O(n2750));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1799_3_lut (.I0(n2646), .I1(n2713_adj_4483), .I2(n2669), 
            .I3(GND_net), .O(n2745));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1803_3_lut (.I0(n2650), .I1(n2717_adj_4481), .I2(n2669), 
            .I3(GND_net), .O(n2749));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1807_3_lut (.I0(n2654), .I1(n2721), .I2(n2669), .I3(GND_net), 
            .O(n2753));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1802_3_lut (.I0(n2649), .I1(n2716), .I2(n2669), .I3(GND_net), 
            .O(n2748));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1735_3_lut (.I0(n2550_adj_4544), .I1(n2617), .I2(n2570), 
            .I3(GND_net), .O(n2649));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1737_3_lut (.I0(n2552_adj_4542), .I1(n2619_adj_4522), 
            .I2(n2570), .I3(GND_net), .O(n2651));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1792_3_lut (.I0(n2639), .I1(n2706_adj_4487), .I2(n2669), 
            .I3(GND_net), .O(n2738));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1791_3_lut (.I0(n2638_adj_4492), .I1(n2705_adj_4488), 
            .I2(n2669), .I3(GND_net), .O(n2737));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1790_3_lut (.I0(n2637_adj_4493), .I1(n2704_adj_4489), 
            .I2(n2669), .I3(GND_net), .O(n2736));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1796_3_lut (.I0(n2643_adj_4490), .I1(n2710), .I2(n2669), 
            .I3(GND_net), .O(n2742));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1794_3_lut (.I0(n2641), .I1(n2708), .I2(n2669), .I3(GND_net), 
            .O(n2740));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1795_3_lut (.I0(n2642_adj_4491), .I1(n2709_adj_4485), 
            .I2(n2669), .I3(GND_net), .O(n2741));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1793_3_lut (.I0(n2640), .I1(n2707_adj_4486), .I2(n2669), 
            .I3(GND_net), .O(n2739));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1809_3_lut (.I0(n2656), .I1(n2723_adj_4479), .I2(n2669), 
            .I3(GND_net), .O(n2755));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1797_3_lut (.I0(n2644), .I1(n2711_adj_4484), .I2(n2669), 
            .I3(GND_net), .O(n2743));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1808_3_lut (.I0(n2655), .I1(n2722), .I2(n2669), .I3(GND_net), 
            .O(n2754));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1738_3_lut (.I0(n2553_adj_4541), .I1(n2620_adj_4521), 
            .I2(n2570), .I3(GND_net), .O(n2652));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1734_3_lut (.I0(n2549_adj_4545), .I1(n2616), .I2(n2570), 
            .I3(GND_net), .O(n2648));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2141_3_lut (.I0(n3148), .I1(n3215), .I2(n3164), .I3(GND_net), 
            .O(n3247));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12908_3_lut (.I0(setpoint[17]), .I1(n4309), .I2(n36839), 
            .I3(GND_net), .O(n17590));   // verilog/coms.v(126[12] 289[6])
    defparam i12908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2149_3_lut (.I0(n3156), .I1(n3223), .I2(n3164), .I3(GND_net), 
            .O(n3255));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2148_3_lut (.I0(n3155), .I1(n3222), .I2(n3164), .I3(GND_net), 
            .O(n3254));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2131_3_lut (.I0(n3138), .I1(n3205), .I2(n3164), .I3(GND_net), 
            .O(n3237));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2135_3_lut (.I0(n3142), .I1(n3209), .I2(n3164), .I3(GND_net), 
            .O(n3241));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2133_3_lut (.I0(n3140), .I1(n3207), .I2(n3164), .I3(GND_net), 
            .O(n3239));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1801_3_lut (.I0(n2648), .I1(n2715_adj_4482), .I2(n2669), 
            .I3(GND_net), .O(n2747));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1806_3_lut (.I0(n2653), .I1(n2720), .I2(n2669), .I3(GND_net), 
            .O(n2752));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1800_3_lut (.I0(n2647), .I1(n2714), .I2(n2669), .I3(GND_net), 
            .O(n2746));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1805_3_lut (.I0(n2652), .I1(n2719_adj_4480), .I2(n2669), 
            .I3(GND_net), .O(n2751));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1723_3_lut (.I0(n2538_adj_4556), .I1(n2605), .I2(n2570), 
            .I3(GND_net), .O(n2637_adj_4493));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1739_3_lut (.I0(n2554), .I1(n2621_adj_4520), .I2(n2570), 
            .I3(GND_net), .O(n2653));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1731_3_lut (.I0(n2546_adj_4548), .I1(n2613), .I2(n2570), 
            .I3(GND_net), .O(n2645));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1729_3_lut (.I0(n2544_adj_4550), .I1(n2611), .I2(n2570), 
            .I3(GND_net), .O(n2643_adj_4490));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1730_3_lut (.I0(n2545_adj_4549), .I1(n2612), .I2(n2570), 
            .I3(GND_net), .O(n2644));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1728_3_lut (.I0(n2543_adj_4551), .I1(n2610), .I2(n2570), 
            .I3(GND_net), .O(n2642_adj_4491));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1736_3_lut (.I0(n2551_adj_4543), .I1(n2618_adj_4523), 
            .I2(n2570), .I3(GND_net), .O(n2650));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1733_3_lut (.I0(n2548_adj_4546), .I1(n2615), .I2(n2570), 
            .I3(GND_net), .O(n2647));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1732_3_lut (.I0(n2547_adj_4547), .I1(n2614), .I2(n2570), 
            .I3(GND_net), .O(n2646));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1743_3_lut (.I0(n2558_adj_4540), .I1(n2625_adj_4516), 
            .I2(n2570), .I3(GND_net), .O(n2657));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1741_3_lut (.I0(n2556), .I1(n2623_adj_4518), .I2(n2570), 
            .I3(GND_net), .O(n2655));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1740_3_lut (.I0(n2555), .I1(n2622_adj_4519), .I2(n2570), 
            .I3(GND_net), .O(n2654));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i11_3_lut (.I0(communication_counter[10]), .I1(n23_adj_4460), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2558_adj_4540));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1643 (.I0(n2556), .I1(n2557), .I2(n2558_adj_4540), 
            .I3(GND_net), .O(n35602));
    defparam i1_3_lut_adj_1643.LUT_INIT = 16'hfefe;
    SB_LUT4 i10_4_lut_adj_1644 (.I0(n2538_adj_4556), .I1(n2539_adj_4555), 
            .I2(n2537_adj_4557), .I3(n2540_adj_4554), .O(n28));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1645 (.I0(n2550_adj_4544), .I1(n2546_adj_4548), 
            .I2(n2553_adj_4541), .I3(n2549_adj_4545), .O(n31_adj_4339));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1646 (.I0(n2543_adj_4551), .I1(n2554), .I2(n35602), 
            .I3(n2555), .O(n22_adj_4340));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1646.LUT_INIT = 16'heaaa;
    SB_LUT4 i12_4_lut_adj_1647 (.I0(n2544_adj_4550), .I1(n2552_adj_4542), 
            .I2(n2547_adj_4547), .I3(n2545_adj_4549), .O(n30));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1648 (.I0(n31_adj_4339), .I1(n2551_adj_4543), 
            .I2(n28), .I3(n2548_adj_4546), .O(n34));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut (.I0(n2541_adj_4553), .I1(n2542_adj_4552), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4341));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_i2139_3_lut (.I0(n3146), .I1(n3213), .I2(n3164), .I3(GND_net), 
            .O(n3245));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2146_3_lut (.I0(n3153), .I1(n3220), .I2(n3164), .I3(GND_net), 
            .O(n3252));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2151_3_lut (.I0(n3158), .I1(n3225), .I2(n3164), .I3(GND_net), 
            .O(n3257));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2150_3_lut (.I0(n3157), .I1(n3224), .I2(n3164), .I3(GND_net), 
            .O(n3256));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1649 (.I0(n3256), .I1(n3257), .I2(n3258), .I3(GND_net), 
            .O(n35699));
    defparam i1_3_lut_adj_1649.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_i1534_3_lut_3_lut (.I0(n2288), .I1(n5974), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i17_4_lut_adj_1650 (.I0(n3252), .I1(n3245), .I2(n3239), .I3(n3241), 
            .O(n42));
    defparam i17_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n3237), .I1(n3254), .I2(n35699), .I3(n3255), 
            .O(n31));
    defparam i6_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 div_46_i1535_3_lut_3_lut (.I0(n2288), .I1(n5975), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13_3_lut (.I0(n3247), .I1(n3231), .I2(n3230), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_i1533_3_lut_3_lut (.I0(n2288), .I1(n5973), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i18_4_lut_adj_1651 (.I0(n3249), .I1(n3248), .I2(n3253), .I3(n3250), 
            .O(n43));
    defparam i18_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1652 (.I0(n21_adj_4341), .I1(n34), .I2(n30), 
            .I3(n22_adj_4340), .O(n2570));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1727_3_lut (.I0(n2542_adj_4552), .I1(n2609), .I2(n2570), 
            .I3(GND_net), .O(n2641));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1725_3_lut (.I0(n2540_adj_4554), .I1(n2607), .I2(n2570), 
            .I3(GND_net), .O(n2639));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1726_3_lut (.I0(n2541_adj_4553), .I1(n2608), .I2(n2570), 
            .I3(GND_net), .O(n2640));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1724_3_lut (.I0(n2539_adj_4555), .I1(n2606), .I2(n2570), 
            .I3(GND_net), .O(n2638_adj_4492));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1742_3_lut (.I0(n2557), .I1(n2624_adj_4517), .I2(n2570), 
            .I3(GND_net), .O(n2656));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1653 (.I0(n2638_adj_4492), .I1(n2640), .I2(n2639), 
            .I3(n2641), .O(n30_adj_5001));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1654 (.I0(n2656), .I1(n2658), .I2(GND_net), .I3(GND_net), 
            .O(n37954));
    defparam i1_2_lut_adj_1654.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(n2654), .I1(n37954), .I2(n2655), .I3(n2657), 
            .O(n35678));
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'ha080;
    SB_LUT4 i15_4_lut (.I0(n2653), .I1(n30_adj_5001), .I2(n2637_adj_4493), 
            .I3(n2636_adj_4502), .O(n34_adj_4997));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1656 (.I0(n2646), .I1(n2647), .I2(n35678), .I3(n2650), 
            .O(n32_adj_4999));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1657 (.I0(n2648), .I1(n2651), .I2(n2652), .I3(n2649), 
            .O(n33_adj_4998));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1658 (.I0(n2642_adj_4491), .I1(n2644), .I2(n2643_adj_4490), 
            .I3(n2645), .O(n31_adj_5000));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1659 (.I0(n31_adj_5000), .I1(n33_adj_4998), .I2(n32_adj_4999), 
            .I3(n34_adj_4997), .O(n2669));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i10_3_lut (.I0(communication_counter[9]), .I1(n24_adj_4459), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2658));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1811_3_lut (.I0(n2658), .I1(n2725), .I2(n2669), .I3(GND_net), 
            .O(n2757));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1810_3_lut (.I0(n2657), .I1(n2724_adj_4478), .I2(n2669), 
            .I3(GND_net), .O(n2756));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1660 (.I0(n2756), .I1(n2757), .I2(n2758), .I3(GND_net), 
            .O(n35615));
    defparam i1_3_lut_adj_1660.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_4_lut_adj_1661 (.I0(n2751), .I1(n2746), .I2(n2752), .I3(n2747), 
            .O(n34_adj_4958));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut_adj_1661.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(n2754), .I1(n2743), .I2(n35615), .I3(n2755), 
            .O(n25_adj_4962));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i12_4_lut_adj_1662 (.I0(n2739), .I1(n2741), .I2(n2740), .I3(n2742), 
            .O(n32_adj_4959));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1663 (.I0(n2736), .I1(n2737), .I2(n2735), .I3(n2738), 
            .O(n31_adj_4960));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1664 (.I0(n2748), .I1(n2753), .I2(n2749), .I3(n2745), 
            .O(n35_adj_4957));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1665 (.I0(n25_adj_4962), .I1(n34_adj_4958), .I2(n2750), 
            .I3(n2744), .O(n37_adj_4955));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1666 (.I0(n37_adj_4955), .I1(n35_adj_4957), .I2(n31_adj_4960), 
            .I3(n32_adj_4959), .O(n2768));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i19_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1667 (.I0(n3234), .I1(n3235), .I2(n3242), .I3(n3243), 
            .O(n40));
    defparam i15_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n31), .I1(n42), .I2(n3244), .I3(n3238), .O(n46));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1668 (.I0(n3236), .I1(n3232), .I2(n3233), .I3(n3240), 
            .O(n39));
    defparam i14_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1669 (.I0(n43), .I1(n3251), .I2(n38), .I3(n3246), 
            .O(n47));
    defparam i22_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i9_3_lut (.I0(communication_counter[8]), .I1(n25_adj_4458), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2758));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1879_3_lut (.I0(n2758), .I1(n2825), .I2(n2768), .I3(GND_net), 
            .O(n2857));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1878_3_lut (.I0(n2757), .I1(n2824), .I2(n2768), .I3(GND_net), 
            .O(n2856));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1670 (.I0(n2856), .I1(n2857), .I2(n2858), .I3(GND_net), 
            .O(n35686));
    defparam i1_3_lut_adj_1670.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1671 (.I0(n2835), .I1(n2834), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4417));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1671.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1672 (.I0(n2854), .I1(n2849), .I2(n35686), .I3(n2855_adj_4474), 
            .O(n28_adj_4416));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1672.LUT_INIT = 16'heccc;
    SB_LUT4 i15_4_lut_adj_1673 (.I0(n2848), .I1(n2847), .I2(n2846), .I3(n2853), 
            .O(n36));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1674 (.I0(n2840), .I1(n2842), .I2(n2841), .I3(n2843), 
            .O(n34_adj_4415));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1675 (.I0(n2836), .I1(n2838), .I2(n2837), .I3(n2839), 
            .O(n33));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1676 (.I0(n2850), .I1(n2852), .I2(n2851), .I3(n22_adj_4417), 
            .O(n37));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1676.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1677 (.I0(n2844), .I1(n36), .I2(n28_adj_4416), 
            .I3(n2845), .O(n39_adj_4414));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n39_adj_4414), .I1(n37), .I2(n33), .I3(n34_adj_4415), 
            .O(n2867));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1859_3_lut (.I0(n2738), .I1(n2805), .I2(n2768), .I3(GND_net), 
            .O(n2837));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1926_3_lut (.I0(n2837), .I1(n2904_adj_4471), .I2(n2867), 
            .I3(GND_net), .O(n2936));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1925_3_lut (.I0(n2836), .I1(n2903_adj_4472), .I2(n2867), 
            .I3(GND_net), .O(n2935));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1924_3_lut (.I0(n2835), .I1(n2902_adj_4473), .I2(n2867), 
            .I3(GND_net), .O(n2934));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1678 (.I0(n2956_adj_4428), .I1(n2957_adj_4427), 
            .I2(n2958_adj_4426), .I3(GND_net), .O(n35632));
    defparam i1_3_lut_adj_1678.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_1679 (.I0(n2941_adj_4443), .I1(n2954_adj_4430), 
            .I2(n35632), .I3(n2955_adj_4429), .O(n27_adj_4942));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut_adj_1679.LUT_INIT = 16'heaaa;
    SB_LUT4 i13_4_lut_adj_1680 (.I0(n2937), .I1(n2939), .I2(n2938), .I3(n2940), 
            .O(n35_adj_4940));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1680.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1681 (.I0(n2934), .I1(n2935), .I2(n2933), .I3(n2936), 
            .O(n34_adj_4941));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1681.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1682 (.I0(n35_adj_4940), .I1(n27_adj_4942), .I2(n2942_adj_4442), 
            .I3(n2943_adj_4441), .O(n40_adj_4922));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1683 (.I0(n2949_adj_4435), .I1(n2947_adj_4437), 
            .I2(n2953_adj_4431), .I3(n2952_adj_4432), .O(n38_adj_4938));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2951_adj_4433), .I1(n34_adj_4941), .I2(n2944_adj_4440), 
            .I3(GND_net), .O(n39_adj_4937));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1684 (.I0(n2948_adj_4436), .I1(n2946_adj_4438), 
            .I2(n2950_adj_4434), .I3(n2945_adj_4439), .O(n37_adj_4939));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1685 (.I0(n37_adj_4939), .I1(n39_adj_4937), .I2(n38_adj_4938), 
            .I3(n40_adj_4922), .O(n2966));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i21_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1538_3_lut_3_lut (.I0(n2288), .I1(n5978), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1589_3_lut_3_lut (.I0(n2381), .I1(n5988), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39), .I2(n46), .I3(n40), .O(n3263));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1583_3_lut_3_lut (.I0(n2381), .I1(n5982), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i7_3_lut (.I0(communication_counter[6]), .I1(n27_adj_4457), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2958_adj_4426));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(one_wire_N_513[5]), .I1(one_wire_N_513[9]), .I2(start), 
            .I3(GND_net), .O(n14_adj_4355));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1686 (.I0(one_wire_N_513[6]), .I1(one_wire_N_513[10]), 
            .I2(one_wire_N_513[8]), .I3(one_wire_N_513[11]), .O(n15_adj_4354));
    defparam i6_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1687 (.I0(n15_adj_4354), .I1(state[1]), .I2(n14_adj_4355), 
            .I3(one_wire_N_513[7]), .O(n35481));
    defparam i8_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1584_3_lut_3_lut (.I0(n2381), .I1(n5983), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1587_3_lut_3_lut (.I0(n2381), .I1(n5986), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1588_3_lut_3_lut (.I0(n2381), .I1(n5987), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1585_3_lut_3_lut (.I0(n2381), .I1(n5984), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i21_3_lut (.I0(communication_counter[20]), .I1(n13_adj_4504), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1558));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1063_3_lut (.I0(n1558), .I1(n1625), .I2(n1580), .I3(GND_net), 
            .O(n1657));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1130_3_lut (.I0(n1657), .I1(n1724), .I2(n1679), .I3(GND_net), 
            .O(n1756_adj_4496));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1197_3_lut (.I0(n1756_adj_4496), .I1(n1823), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i8_3_lut (.I0(communication_counter[7]), .I1(n26), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2858));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1586_3_lut_3_lut (.I0(n2381), .I1(n5985), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1653_17 (.CI(n28950), .I0(n2444), .I1(n2471_adj_4558), 
            .CO(n28951));
    SB_LUT4 communication_counter_1176_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[16]), .I3(n28635), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_559_6 (.CI(n28114), .I0(n43079), .I1(n21), .CO(n28115));
    SB_LUT4 rem_4_add_1653_16_lut (.I0(n2445), .I1(n2445), .I2(n2471_adj_4558), 
            .I3(n28949), .O(n2544_adj_4550)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_559_5_lut (.I0(duty[3]), .I1(n43079), .I2(n22), .I3(n28113), 
            .O(pwm_setpoint_22__N_57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1653_16 (.CI(n28949), .I0(n2445), .I1(n2471_adj_4558), 
            .CO(n28950));
    SB_LUT4 rem_4_add_1653_15_lut (.I0(n2446), .I1(n2446), .I2(n2471_adj_4558), 
            .I3(n28948), .O(n2545_adj_4549)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_559_5 (.CI(n28113), .I0(n43079), .I1(n22), .CO(n28114));
    SB_CARRY rem_4_add_1653_15 (.CI(n28948), .I0(n2446), .I1(n2471_adj_4558), 
            .CO(n28949));
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_229[0]), 
            .I1(n25_adj_4408), .CO(n28202));
    SB_LUT4 rem_4_add_1653_14_lut (.I0(n2447_adj_4571), .I1(n2447_adj_4571), 
            .I2(n2471_adj_4558), .I3(n28947), .O(n2546_adj_4548)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1653_14 (.CI(n28947), .I0(n2447_adj_4571), .I1(n2471_adj_4558), 
            .CO(n28948));
    SB_LUT4 div_46_i1594_3_lut_3_lut (.I0(n2381), .I1(n5993), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[21]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_106[21]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1595_3_lut_3_lut (.I0(n2381), .I1(n5994), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36321_1_lut (.I0(n2471_adj_4558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n43083));
    defparam i36321_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_559_4_lut (.I0(duty[2]), .I1(n43079), .I2(n23), .I3(n28112), 
            .O(pwm_setpoint_22__N_57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1653_13_lut (.I0(n2448_adj_4570), .I1(n2448_adj_4570), 
            .I2(n2471_adj_4558), .I3(n28946), .O(n2547_adj_4547)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY communication_counter_1176_add_4_18 (.CI(n28635), .I0(GND_net), 
            .I1(communication_counter[16]), .CO(n28636));
    SB_LUT4 i12907_3_lut (.I0(setpoint[16]), .I1(n4308), .I2(n36839), 
            .I3(GND_net), .O(n17589));   // verilog/coms.v(126[12] 289[6])
    defparam i12907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1600_3_lut_3_lut (.I0(n2381), .I1(n5999), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i584_3_lut (.I0(n852), .I1(n6_adj_4410), .I2(n884), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i584_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_3_lut_adj_1688 (.I0(n1056), .I1(n1057), .I2(n1058), .I3(GND_net), 
            .O(n35534));
    defparam i1_3_lut_adj_1688.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1689 (.I0(n1054), .I1(n1055), .I2(GND_net), .I3(GND_net), 
            .O(n37550));
    defparam i1_2_lut_adj_1689.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n1052), .I1(n37550), .I2(n1053), .I3(n35534), 
            .O(n1085));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'hfefa;
    SB_LUT4 unary_minus_28_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_4337));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1653_13 (.CI(n28946), .I0(n2448_adj_4570), .I1(n2471_adj_4558), 
            .CO(n28947));
    SB_LUT4 communication_counter_1176_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[15]), .I3(n28634), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_12_lut (.I0(n2449_adj_4569), .I1(n2449_adj_4569), 
            .I2(n2471_adj_4558), .I3(n28945), .O(n2548_adj_4546)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY communication_counter_1176_add_4_17 (.CI(n28634), .I0(GND_net), 
            .I1(communication_counter[15]), .CO(n28635));
    SB_LUT4 communication_counter_1176_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[14]), .I3(n28633), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_16 (.CI(n28633), .I0(GND_net), 
            .I1(communication_counter[14]), .CO(n28634));
    SB_LUT4 communication_counter_1176_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[13]), .I3(n28632), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_12 (.CI(n28945), .I0(n2449_adj_4569), .I1(n2471_adj_4558), 
            .CO(n28946));
    SB_CARRY communication_counter_1176_add_4_15 (.CI(n28632), .I0(GND_net), 
            .I1(communication_counter[13]), .CO(n28633));
    SB_LUT4 div_46_i1599_3_lut_3_lut (.I0(n2381), .I1(n5998), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1176_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[12]), .I3(n28631), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_14 (.CI(n28631), .I0(GND_net), 
            .I1(communication_counter[12]), .CO(n28632));
    SB_LUT4 rem_4_add_1653_11_lut (.I0(n2450_adj_4568), .I1(n2450_adj_4568), 
            .I2(n2471_adj_4558), .I3(n28944), .O(n2549_adj_4545)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1653_11 (.CI(n28944), .I0(n2450_adj_4568), .I1(n2471_adj_4558), 
            .CO(n28945));
    SB_CARRY add_559_4 (.CI(n28112), .I0(n43079), .I1(n23), .CO(n28113));
    SB_LUT4 communication_counter_1176_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[11]), .I3(n28630), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_13 (.CI(n28630), .I0(GND_net), 
            .I1(communication_counter[11]), .CO(n28631));
    SB_LUT4 div_46_i1598_3_lut_3_lut (.I0(n2381), .I1(n5997), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 communication_counter_1176_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[10]), .I3(n28629), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_559_3_lut (.I0(duty[1]), .I1(n43079), .I2(n24_adj_4337), 
            .I3(n28111), .O(pwm_setpoint_22__N_57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1653_10_lut (.I0(n2451_adj_4567), .I1(n2451_adj_4567), 
            .I2(n2471_adj_4558), .I3(n28943), .O(n2550_adj_4544)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1653_10 (.CI(n28943), .I0(n2451_adj_4567), .I1(n2471_adj_4558), 
            .CO(n28944));
    SB_LUT4 rem_4_add_1653_9_lut (.I0(n2452_adj_4566), .I1(n2452_adj_4566), 
            .I2(n2471_adj_4558), .I3(n28942), .O(n2551_adj_4543)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_559_3 (.CI(n28111), .I0(n43079), .I1(n24_adj_4337), .CO(n28112));
    SB_CARRY rem_4_add_1653_9 (.CI(n28942), .I0(n2452_adj_4566), .I1(n2471_adj_4558), 
            .CO(n28943));
    SB_LUT4 rem_4_add_1653_8_lut (.I0(n2453_adj_4565), .I1(n2453_adj_4565), 
            .I2(n2471_adj_4558), .I3(n28941), .O(n2552_adj_4542)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY communication_counter_1176_add_4_12 (.CI(n28629), .I0(GND_net), 
            .I1(communication_counter[10]), .CO(n28630));
    SB_LUT4 communication_counter_1176_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[9]), .I3(n28628), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_8 (.CI(n28941), .I0(n2453_adj_4565), .I1(n2471_adj_4558), 
            .CO(n28942));
    SB_CARRY communication_counter_1176_add_4_11 (.CI(n28628), .I0(GND_net), 
            .I1(communication_counter[9]), .CO(n28629));
    SB_LUT4 rem_4_add_1653_7_lut (.I0(n2454_adj_4564), .I1(n2454_adj_4564), 
            .I2(n43083), .I3(n28940), .O(n2553_adj_4541)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1653_7 (.CI(n28940), .I0(n2454_adj_4564), .I1(n43083), 
            .CO(n28941));
    SB_LUT4 rem_4_add_1653_6_lut (.I0(n2455_adj_4563), .I1(n2455_adj_4563), 
            .I2(n43083), .I3(n28939), .O(n2554)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1653_6 (.CI(n28939), .I0(n2455_adj_4563), .I1(n43083), 
            .CO(n28940));
    SB_LUT4 rem_4_add_1653_5_lut (.I0(n2456_adj_4562), .I1(n2456_adj_4562), 
            .I2(n2471_adj_4558), .I3(n28938), .O(n2555)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1653_5 (.CI(n28938), .I0(n2456_adj_4562), .I1(n2471_adj_4558), 
            .CO(n28939));
    SB_LUT4 add_559_2_lut (.I0(duty[0]), .I1(n43079), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_559_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_559_2 (.CI(VCC_net), .I0(n43079), .I1(n25), .CO(n28111));
    SB_LUT4 communication_counter_1176_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[8]), .I3(n28627), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_4_lut (.I0(n2457_adj_4561), .I1(n2457_adj_4561), 
            .I2(n2471_adj_4558), .I3(n28937), .O(n2556)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1653_4 (.CI(n28937), .I0(n2457_adj_4561), .I1(n2471_adj_4558), 
            .CO(n28938));
    SB_LUT4 rem_4_add_1653_3_lut (.I0(n2458_adj_4560), .I1(n2458_adj_4560), 
            .I2(n43083), .I3(n28936), .O(n2557)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY rem_4_add_1653_3 (.CI(n28936), .I0(n2458_adj_4560), .I1(n43083), 
            .CO(n28937));
    SB_CARRY communication_counter_1176_add_4_10 (.CI(n28627), .I0(GND_net), 
            .I1(communication_counter[8]), .CO(n28628));
    SB_CARRY rem_4_add_1653_2 (.CI(VCC_net), .I0(n2558_adj_4540), .I1(VCC_net), 
            .CO(n28936));
    SB_LUT4 communication_counter_1176_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[7]), .I3(n28626), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_9 (.CI(n28626), .I0(GND_net), 
            .I1(communication_counter[7]), .CO(n28627));
    SB_LUT4 rem_4_add_1720_24_lut (.I0(n2570), .I1(n2537_adj_4557), .I2(VCC_net), 
            .I3(n28935), .O(n2636_adj_4502)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_1176_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[6]), .I3(n28625), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_8 (.CI(n28625), .I0(GND_net), 
            .I1(communication_counter[6]), .CO(n28626));
    SB_LUT4 communication_counter_1176_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[5]), .I3(n28624), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_23_lut (.I0(GND_net), .I1(n2538_adj_4556), .I2(VCC_net), 
            .I3(n28934), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_7 (.CI(n28624), .I0(GND_net), 
            .I1(communication_counter[5]), .CO(n28625));
    SB_CARRY rem_4_add_1720_23 (.CI(n28934), .I0(n2538_adj_4556), .I1(VCC_net), 
            .CO(n28935));
    SB_LUT4 rem_4_add_1720_22_lut (.I0(GND_net), .I1(n2539_adj_4555), .I2(VCC_net), 
            .I3(n28933), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_22 (.CI(n28933), .I0(n2539_adj_4555), .I1(VCC_net), 
            .CO(n28934));
    SB_LUT4 communication_counter_1176_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[4]), .I3(n28623), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_6 (.CI(n28623), .I0(GND_net), 
            .I1(communication_counter[4]), .CO(n28624));
    SB_LUT4 communication_counter_1176_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[3]), .I3(n28622), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_21_lut (.I0(GND_net), .I1(n2540_adj_4554), .I2(VCC_net), 
            .I3(n28932), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_5 (.CI(n28622), .I0(GND_net), 
            .I1(communication_counter[3]), .CO(n28623));
    SB_LUT4 communication_counter_1176_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[2]), .I3(n28621), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_4 (.CI(n28621), .I0(GND_net), 
            .I1(communication_counter[2]), .CO(n28622));
    SB_LUT4 communication_counter_1176_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[1]), .I3(n28620), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_3 (.CI(n28620), .I0(GND_net), 
            .I1(communication_counter[1]), .CO(n28621));
    SB_LUT4 communication_counter_1176_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1176_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1176_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(communication_counter[0]), .CO(n28620));
    SB_LUT4 rem_4_add_2189_30_lut (.I0(n3263), .I1(n3230), .I2(VCC_net), 
            .I3(n28619), .O(n37992)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1720_21 (.CI(n28932), .I0(n2540_adj_4554), .I1(VCC_net), 
            .CO(n28933));
    SB_LUT4 rem_4_add_2189_29_lut (.I0(GND_net), .I1(n3231), .I2(VCC_net), 
            .I3(n28618), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_20_lut (.I0(GND_net), .I1(n2541_adj_4553), .I2(VCC_net), 
            .I3(n28931), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_29 (.CI(n28618), .I0(n3231), .I1(VCC_net), 
            .CO(n28619));
    SB_CARRY rem_4_add_1720_20 (.CI(n28931), .I0(n2541_adj_4553), .I1(VCC_net), 
            .CO(n28932));
    SB_LUT4 rem_4_add_2189_28_lut (.I0(GND_net), .I1(n3232), .I2(VCC_net), 
            .I3(n28617), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_28 (.CI(n28617), .I0(n3232), .I1(VCC_net), 
            .CO(n28618));
    SB_LUT4 rem_4_add_2189_27_lut (.I0(GND_net), .I1(n3233), .I2(VCC_net), 
            .I3(n28616), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_27 (.CI(n28616), .I0(n3233), .I1(VCC_net), 
            .CO(n28617));
    SB_LUT4 rem_4_add_2189_26_lut (.I0(GND_net), .I1(n3234), .I2(VCC_net), 
            .I3(n28615), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1601_3_lut_3_lut (.I0(n2381), .I1(n6000), .I2(n665), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2189_26 (.CI(n28615), .I0(n3234), .I1(VCC_net), 
            .CO(n28616));
    SB_LUT4 rem_4_add_2189_25_lut (.I0(GND_net), .I1(n3235), .I2(VCC_net), 
            .I3(n28614), .O(n3302)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_25 (.CI(n28614), .I0(n3235), .I1(VCC_net), 
            .CO(n28615));
    SB_LUT4 rem_4_add_2189_24_lut (.I0(GND_net), .I1(n3236), .I2(VCC_net), 
            .I3(n28613), .O(n3303)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_24 (.CI(n28613), .I0(n3236), .I1(VCC_net), 
            .CO(n28614));
    SB_LUT4 rem_4_add_2189_23_lut (.I0(GND_net), .I1(n3237), .I2(VCC_net), 
            .I3(n28612), .O(n3304)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_23 (.CI(n28612), .I0(n3237), .I1(VCC_net), 
            .CO(n28613));
    SB_LUT4 rem_4_add_2189_22_lut (.I0(GND_net), .I1(n3238), .I2(VCC_net), 
            .I3(n28611), .O(n3305)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_22 (.CI(n28611), .I0(n3238), .I1(VCC_net), 
            .CO(n28612));
    SB_LUT4 rem_4_add_2189_21_lut (.I0(GND_net), .I1(n3239), .I2(VCC_net), 
            .I3(n28610), .O(n3306)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1593_3_lut_3_lut (.I0(n2381), .I1(n5992), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1720_19_lut (.I0(GND_net), .I1(n2542_adj_4552), .I2(VCC_net), 
            .I3(n28930), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_21 (.CI(n28610), .I0(n3239), .I1(VCC_net), 
            .CO(n28611));
    SB_LUT4 div_46_i1592_3_lut_3_lut (.I0(n2381), .I1(n5991), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1720_19 (.CI(n28930), .I0(n2542_adj_4552), .I1(VCC_net), 
            .CO(n28931));
    SB_LUT4 rem_4_add_1720_18_lut (.I0(GND_net), .I1(n2543_adj_4551), .I2(VCC_net), 
            .I3(n28929), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_18 (.CI(n28929), .I0(n2543_adj_4551), .I1(VCC_net), 
            .CO(n28930));
    SB_LUT4 rem_4_add_1720_17_lut (.I0(GND_net), .I1(n2544_adj_4550), .I2(VCC_net), 
            .I3(n28928), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_20_lut (.I0(GND_net), .I1(n3240), .I2(VCC_net), 
            .I3(n28609), .O(n3307)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_17 (.CI(n28928), .I0(n2544_adj_4550), .I1(VCC_net), 
            .CO(n28929));
    SB_LUT4 rem_4_add_1720_16_lut (.I0(GND_net), .I1(n2545_adj_4549), .I2(VCC_net), 
            .I3(n28927), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_20 (.CI(n28609), .I0(n3240), .I1(VCC_net), 
            .CO(n28610));
    SB_CARRY rem_4_add_1720_16 (.CI(n28927), .I0(n2545_adj_4549), .I1(VCC_net), 
            .CO(n28928));
    SB_LUT4 unary_minus_28_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_71_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[22]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_106[22]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1597_3_lut_3_lut (.I0(n2381), .I1(n5996), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12906_3_lut (.I0(setpoint[15]), .I1(n4307), .I2(n36839), 
            .I3(GND_net), .O(n17588));   // verilog/coms.v(126[12] 289[6])
    defparam i12906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1691 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4951));   // verilog/TinyFPGA_B.v(229[5:22])
    defparam i4_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1692 (.I0(control_mode[6]), .I1(n10_adj_4951), 
            .I2(control_mode[2]), .I3(GND_net), .O(n15508));   // verilog/TinyFPGA_B.v(229[5:22])
    defparam i5_3_lut_adj_1692.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_mux_3_i26_3_lut (.I0(communication_counter[25]), .I1(n8_adj_4509), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1058));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n15508), 
            .I3(GND_net), .O(n15_adj_4322));   // verilog/TinyFPGA_B.v(229[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_71_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[23]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_106[23]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1596_3_lut_3_lut (.I0(n2381), .I1(n5995), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1591_3_lut_3_lut (.I0(n2381), .I1(n5990), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4408));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12373_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n37092), .I3(GND_net), .O(n17055));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12374_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n37092), .I3(GND_net), .O(n17056));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12375_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n37092), .I3(GND_net), .O(n17057));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12376_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n37092), .I3(GND_net), .O(n17058));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12377_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n37092), .I3(GND_net), .O(n17059));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12378_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n37092), .I3(GND_net), .O(n17060));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1590_3_lut_3_lut (.I0(n2381), .I1(n5989), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12379_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n37092), .I3(GND_net), .O(n17061));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12380_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n37092), .I3(GND_net), .O(n17062));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i22_3_lut (.I0(communication_counter[21]), .I1(n12_adj_4505), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i995_3_lut (.I0(n1458), .I1(n1525), .I2(n1481), .I3(GND_net), 
            .O(n1557));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1062_3_lut (.I0(n1557), .I1(n1624), .I2(n1580), .I3(GND_net), 
            .O(n1656));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1129_3_lut (.I0(n1656), .I1(n1723), .I2(n1679), .I3(GND_net), 
            .O(n1755_adj_4495));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12381_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n37092), .I3(GND_net), .O(n17063));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36309_1_lut (.I0(n1877), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43071));
    defparam i36309_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12382_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n37092), .I3(GND_net), .O(n17064));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12383_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n37092), .I3(GND_net), .O(n17065));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12384_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n37092), .I3(GND_net), .O(n17066));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12385_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n37092), .I3(GND_net), .O(n17067));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12386_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n37092), .I3(GND_net), .O(n17068));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12387_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n37092), .I3(GND_net), .O(n17069));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12388_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n37092), .I3(GND_net), .O(n17070));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12389_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n37092), .I3(GND_net), .O(n17071));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1649_3_lut_3_lut (.I0(n2471), .I1(n6010), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12390_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n37092), .I3(GND_net), .O(n17072));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12390_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1642_3_lut_3_lut (.I0(n2471), .I1(n6003), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_19_lut (.I0(GND_net), .I1(n3241), .I2(VCC_net), 
            .I3(n28608), .O(n3308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1644_3_lut_3_lut (.I0(n2471), .I1(n6005), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i24_3_lut_adj_1693 (.I0(n40172), .I1(bit_ctr[9]), .I2(n4385), 
            .I3(GND_net), .O(n33325));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1693.LUT_INIT = 16'hcaca;
    SB_LUT4 i12838_3_lut (.I0(encoder0_position[19]), .I1(n2945), .I2(count_enable), 
            .I3(GND_net), .O(n17520));   // quad.v(35[10] 41[6])
    defparam i12838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12392_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17074));   // verilog/coms.v(126[12] 289[6])
    defparam i12392_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12393_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17075));   // verilog/coms.v(126[12] 289[6])
    defparam i12393_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12394_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17076));   // verilog/coms.v(126[12] 289[6])
    defparam i12394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12395_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17077));   // verilog/coms.v(126[12] 289[6])
    defparam i12395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12396_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17078));   // verilog/coms.v(126[12] 289[6])
    defparam i12396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12397_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17079));   // verilog/coms.v(126[12] 289[6])
    defparam i12397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1643_3_lut_3_lut (.I0(n2471), .I1(n6004), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12398_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17080));   // verilog/coms.v(126[12] 289[6])
    defparam i12398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12399_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n36885), .I3(GND_net), .O(n17081));   // verilog/coms.v(126[12] 289[6])
    defparam i12399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12400_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17082));   // verilog/coms.v(126[12] 289[6])
    defparam i12400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12401_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17083));   // verilog/coms.v(126[12] 289[6])
    defparam i12401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4336));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12402_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17084));   // verilog/coms.v(126[12] 289[6])
    defparam i12402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12403_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17085));   // verilog/coms.v(126[12] 289[6])
    defparam i12403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1647_3_lut_3_lut (.I0(n2471), .I1(n6008), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12404_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17086));   // verilog/coms.v(126[12] 289[6])
    defparam i12404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12405_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17087));   // verilog/coms.v(126[12] 289[6])
    defparam i12405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12837_3_lut (.I0(encoder0_position[18]), .I1(n2946), .I2(count_enable), 
            .I3(GND_net), .O(n17519));   // quad.v(35[10] 41[6])
    defparam i12837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12406_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17088));   // verilog/coms.v(126[12] 289[6])
    defparam i12406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1645_3_lut_3_lut (.I0(n2471), .I1(n6006), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12910_3_lut (.I0(setpoint[19]), .I1(n4311), .I2(n36839), 
            .I3(GND_net), .O(n17592));   // verilog/coms.v(126[12] 289[6])
    defparam i12910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12407_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n36885), .I3(GND_net), .O(n17089));   // verilog/coms.v(126[12] 289[6])
    defparam i12407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12408_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17090));   // verilog/coms.v(126[12] 289[6])
    defparam i12408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12409_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17091));   // verilog/coms.v(126[12] 289[6])
    defparam i12409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12410_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17092));   // verilog/coms.v(126[12] 289[6])
    defparam i12410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4407));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_2189_19 (.CI(n28608), .I0(n3241), .I1(VCC_net), 
            .CO(n28609));
    SB_LUT4 i12411_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17093));   // verilog/coms.v(126[12] 289[6])
    defparam i12411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1648_3_lut_3_lut (.I0(n2471), .I1(n6009), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1720_15_lut (.I0(GND_net), .I1(n2546_adj_4548), .I2(VCC_net), 
            .I3(n28926), .O(n2613)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12412_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17094));   // verilog/coms.v(126[12] 289[6])
    defparam i12412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1661_3_lut_3_lut (.I0(n2471), .I1(n6022), .I2(n666), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1720_15 (.CI(n28926), .I0(n2546_adj_4548), .I1(VCC_net), 
            .CO(n28927));
    SB_LUT4 i12413_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17095));   // verilog/coms.v(126[12] 289[6])
    defparam i12413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2189_18_lut (.I0(GND_net), .I1(n3242), .I2(VCC_net), 
            .I3(n28607), .O(n3309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_14_lut (.I0(GND_net), .I1(n2547_adj_4547), .I2(VCC_net), 
            .I3(n28925), .O(n2614)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1646_3_lut_3_lut (.I0(n2471), .I1(n6007), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12414_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17096));   // verilog/coms.v(126[12] 289[6])
    defparam i12414_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2189_18 (.CI(n28607), .I0(n3242), .I1(VCC_net), 
            .CO(n28608));
    SB_LUT4 i12415_3_lut (.I0(gearBoxRatio[1]), .I1(\data_in_frame[19] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17097));   // verilog/coms.v(126[12] 289[6])
    defparam i12415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1650_3_lut_3_lut (.I0(n2471), .I1(n6011), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12416_3_lut (.I0(gearBoxRatio[2]), .I1(\data_in_frame[19] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17098));   // verilog/coms.v(126[12] 289[6])
    defparam i12416_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12417_3_lut (.I0(gearBoxRatio[3]), .I1(\data_in_frame[19] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17099));   // verilog/coms.v(126[12] 289[6])
    defparam i12417_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1651_3_lut_3_lut (.I0(n2471), .I1(n6012), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12418_3_lut (.I0(gearBoxRatio[4]), .I1(\data_in_frame[19] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17100));   // verilog/coms.v(126[12] 289[6])
    defparam i12418_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_28_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4335));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2189_17_lut (.I0(GND_net), .I1(n3243), .I2(VCC_net), 
            .I3(n28606), .O(n3310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_14 (.CI(n28925), .I0(n2547_adj_4547), .I1(VCC_net), 
            .CO(n28926));
    SB_LUT4 rem_4_add_1720_13_lut (.I0(GND_net), .I1(n2548_adj_4546), .I2(VCC_net), 
            .I3(n28924), .O(n2615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_13 (.CI(n28924), .I0(n2548_adj_4546), .I1(VCC_net), 
            .CO(n28925));
    SB_LUT4 rem_4_add_1720_12_lut (.I0(GND_net), .I1(n2549_adj_4545), .I2(VCC_net), 
            .I3(n28923), .O(n2616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_17 (.CI(n28606), .I0(n3243), .I1(VCC_net), 
            .CO(n28607));
    SB_LUT4 i12419_3_lut (.I0(gearBoxRatio[5]), .I1(\data_in_frame[19] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17101));   // verilog/coms.v(126[12] 289[6])
    defparam i12419_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_2189_16_lut (.I0(GND_net), .I1(n3244), .I2(VCC_net), 
            .I3(n28605), .O(n3311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_16 (.CI(n28605), .I0(n3244), .I1(VCC_net), 
            .CO(n28606));
    SB_LUT4 rem_4_add_2189_15_lut (.I0(GND_net), .I1(n3245), .I2(VCC_net), 
            .I3(n28604), .O(n3312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_15 (.CI(n28604), .I0(n3245), .I1(VCC_net), 
            .CO(n28605));
    SB_LUT4 rem_4_add_2189_14_lut (.I0(GND_net), .I1(n3246), .I2(VCC_net), 
            .I3(n28603), .O(n3313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_12 (.CI(n28923), .I0(n2549_adj_4545), .I1(VCC_net), 
            .CO(n28924));
    SB_LUT4 rem_4_add_1720_11_lut (.I0(GND_net), .I1(n2550_adj_4544), .I2(VCC_net), 
            .I3(n28922), .O(n2617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12420_3_lut (.I0(gearBoxRatio[6]), .I1(\data_in_frame[19] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17102));   // verilog/coms.v(126[12] 289[6])
    defparam i12420_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2189_14 (.CI(n28603), .I0(n3246), .I1(VCC_net), 
            .CO(n28604));
    SB_LUT4 rem_4_add_2189_13_lut (.I0(GND_net), .I1(n3247), .I2(VCC_net), 
            .I3(n28602), .O(n3314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_13 (.CI(n28602), .I0(n3247), .I1(VCC_net), 
            .CO(n28603));
    SB_LUT4 rem_4_add_2189_12_lut (.I0(GND_net), .I1(n3248), .I2(VCC_net), 
            .I3(n28601), .O(n3315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12421_3_lut (.I0(gearBoxRatio[7]), .I1(\data_in_frame[19] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17103));   // verilog/coms.v(126[12] 289[6])
    defparam i12421_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_2189_12 (.CI(n28601), .I0(n3248), .I1(VCC_net), 
            .CO(n28602));
    SB_CARRY rem_4_add_1720_11 (.CI(n28922), .I0(n2550_adj_4544), .I1(VCC_net), 
            .CO(n28923));
    SB_LUT4 rem_4_add_2189_11_lut (.I0(GND_net), .I1(n3249), .I2(VCC_net), 
            .I3(n28600), .O(n3316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12909_3_lut (.I0(setpoint[18]), .I1(n4310), .I2(n36839), 
            .I3(GND_net), .O(n17591));   // verilog/coms.v(126[12] 289[6])
    defparam i12909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1656_3_lut_3_lut (.I0(n2471), .I1(n6017), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1653_3_lut_3_lut (.I0(n2471), .I1(n6014), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12422_3_lut (.I0(gearBoxRatio[8]), .I1(\data_in_frame[18] [0]), 
            .I2(n36885), .I3(GND_net), .O(n17104));   // verilog/coms.v(126[12] 289[6])
    defparam i12422_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12423_3_lut (.I0(gearBoxRatio[9]), .I1(\data_in_frame[18] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17105));   // verilog/coms.v(126[12] 289[6])
    defparam i12423_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1652_3_lut_3_lut (.I0(n2471), .I1(n6013), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1720_10_lut (.I0(GND_net), .I1(n2551_adj_4543), .I2(VCC_net), 
            .I3(n28921), .O(n2618_adj_4523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_10 (.CI(n28921), .I0(n2551_adj_4543), .I1(VCC_net), 
            .CO(n28922));
    SB_LUT4 rem_4_add_1720_9_lut (.I0(GND_net), .I1(n2552_adj_4542), .I2(VCC_net), 
            .I3(n28920), .O(n2619_adj_4522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_11 (.CI(n28600), .I0(n3249), .I1(VCC_net), 
            .CO(n28601));
    SB_CARRY rem_4_add_1720_9 (.CI(n28920), .I0(n2552_adj_4542), .I1(VCC_net), 
            .CO(n28921));
    SB_LUT4 rem_4_add_1720_8_lut (.I0(GND_net), .I1(n2553_adj_4541), .I2(VCC_net), 
            .I3(n28919), .O(n2620_adj_4521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_10_lut (.I0(GND_net), .I1(n3250), .I2(VCC_net), 
            .I3(n28599), .O(n3317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_8 (.CI(n28919), .I0(n2553_adj_4541), .I1(VCC_net), 
            .CO(n28920));
    SB_CARRY rem_4_add_2189_10 (.CI(n28599), .I0(n3250), .I1(VCC_net), 
            .CO(n28600));
    SB_LUT4 rem_4_add_1720_7_lut (.I0(GND_net), .I1(n2554), .I2(GND_net), 
            .I3(n28918), .O(n2621_adj_4520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_7 (.CI(n28918), .I0(n2554), .I1(GND_net), 
            .CO(n28919));
    SB_LUT4 rem_4_add_1720_6_lut (.I0(GND_net), .I1(n2555), .I2(GND_net), 
            .I3(n28917), .O(n2622_adj_4519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_6 (.CI(n28917), .I0(n2555), .I1(GND_net), 
            .CO(n28918));
    SB_LUT4 rem_4_add_1720_5_lut (.I0(GND_net), .I1(n2556), .I2(VCC_net), 
            .I3(n28916), .O(n2623_adj_4518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12424_3_lut (.I0(gearBoxRatio[10]), .I1(\data_in_frame[18] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17106));   // verilog/coms.v(126[12] 289[6])
    defparam i12424_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1720_5 (.CI(n28916), .I0(n2556), .I1(VCC_net), 
            .CO(n28917));
    SB_LUT4 rem_4_add_1720_4_lut (.I0(GND_net), .I1(n2557), .I2(VCC_net), 
            .I3(n28915), .O(n2624_adj_4517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_11_lut (.I0(n1382), .I1(n1349), .I2(VCC_net), 
            .I3(n27989), .O(n1448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1720_4 (.CI(n28915), .I0(n2557), .I1(VCC_net), 
            .CO(n28916));
    SB_LUT4 div_46_i1660_3_lut_3_lut (.I0(n2471), .I1(n6021), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_9_lut (.I0(GND_net), .I1(n3251), .I2(VCC_net), 
            .I3(n28598), .O(n3318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_10_lut (.I0(GND_net), .I1(n1350), .I2(VCC_net), 
            .I3(n27988), .O(n1417_adj_4536)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12425_3_lut (.I0(gearBoxRatio[11]), .I1(\data_in_frame[18] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17107));   // verilog/coms.v(126[12] 289[6])
    defparam i12425_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1720_3_lut (.I0(GND_net), .I1(n2558_adj_4540), .I2(GND_net), 
            .I3(n28914), .O(n2625_adj_4516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_9 (.CI(n28598), .I0(n3251), .I1(VCC_net), 
            .CO(n28599));
    SB_CARRY rem_4_add_1720_3 (.CI(n28914), .I0(n2558_adj_4540), .I1(GND_net), 
            .CO(n28915));
    SB_LUT4 rem_4_add_2189_8_lut (.I0(GND_net), .I1(n3252), .I2(VCC_net), 
            .I3(n28597), .O(n3319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1659_3_lut_3_lut (.I0(n2471), .I1(n6020), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2189_8 (.CI(n28597), .I0(n3252), .I1(VCC_net), 
            .CO(n28598));
    SB_LUT4 rem_4_add_2189_7_lut (.I0(GND_net), .I1(n3253), .I2(VCC_net), 
            .I3(n28596), .O(n3320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_7 (.CI(n28596), .I0(n3253), .I1(VCC_net), 
            .CO(n28597));
    SB_CARRY rem_4_add_1720_2 (.CI(VCC_net), .I0(n2658), .I1(VCC_net), 
            .CO(n28914));
    SB_LUT4 rem_4_add_1787_25_lut (.I0(n2669), .I1(n2636_adj_4502), .I2(VCC_net), 
            .I3(n28913), .O(n2735)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1787_24_lut (.I0(GND_net), .I1(n2637_adj_4493), .I2(VCC_net), 
            .I3(n28912), .O(n2704_adj_4489)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_24 (.CI(n28912), .I0(n2637_adj_4493), .I1(VCC_net), 
            .CO(n28913));
    SB_CARRY rem_4_add_916_10 (.CI(n27988), .I0(n1350), .I1(VCC_net), 
            .CO(n27989));
    SB_LUT4 rem_4_add_2189_6_lut (.I0(GND_net), .I1(n3254), .I2(GND_net), 
            .I3(n28595), .O(n3321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_6 (.CI(n28595), .I0(n3254), .I1(GND_net), 
            .CO(n28596));
    SB_LUT4 rem_4_add_2189_5_lut (.I0(GND_net), .I1(n3255), .I2(GND_net), 
            .I3(n28594), .O(n3322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_23_lut (.I0(GND_net), .I1(n2638_adj_4492), .I2(VCC_net), 
            .I3(n28911), .O(n2705_adj_4488)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_5 (.CI(n28594), .I0(n3255), .I1(GND_net), 
            .CO(n28595));
    SB_CARRY rem_4_add_1787_23 (.CI(n28911), .I0(n2638_adj_4492), .I1(VCC_net), 
            .CO(n28912));
    SB_LUT4 rem_4_add_1787_22_lut (.I0(GND_net), .I1(n2639), .I2(VCC_net), 
            .I3(n28910), .O(n2706_adj_4487)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_22 (.CI(n28910), .I0(n2639), .I1(VCC_net), 
            .CO(n28911));
    SB_LUT4 rem_4_add_1787_21_lut (.I0(GND_net), .I1(n2640), .I2(VCC_net), 
            .I3(n28909), .O(n2707_adj_4486)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_21 (.CI(n28909), .I0(n2640), .I1(VCC_net), 
            .CO(n28910));
    SB_LUT4 rem_4_add_1787_20_lut (.I0(GND_net), .I1(n2641), .I2(VCC_net), 
            .I3(n28908), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_20 (.CI(n28908), .I0(n2641), .I1(VCC_net), 
            .CO(n28909));
    SB_LUT4 rem_4_add_1787_19_lut (.I0(GND_net), .I1(n2642_adj_4491), .I2(VCC_net), 
            .I3(n28907), .O(n2709_adj_4485)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_4_lut (.I0(GND_net), .I1(n3256), .I2(VCC_net), 
            .I3(n28593), .O(n3323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_4 (.CI(n28593), .I0(n3256), .I1(VCC_net), 
            .CO(n28594));
    SB_LUT4 rem_4_add_2189_3_lut (.I0(GND_net), .I1(n3257), .I2(VCC_net), 
            .I3(n28592), .O(n3324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_3 (.CI(n28592), .I0(n3257), .I1(VCC_net), 
            .CO(n28593));
    SB_LUT4 rem_4_add_2189_2_lut (.I0(GND_net), .I1(n3258), .I2(GND_net), 
            .I3(VCC_net), .O(n3325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_2 (.CI(VCC_net), .I0(n3258), .I1(GND_net), 
            .CO(n28592));
    SB_LUT4 rem_4_add_2298_9_lut (.I0(n43021), .I1(n2_adj_4965), .I2(n3452), 
            .I3(n28591), .O(color_23__N_164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_2298_8_lut (.I0(n43025), .I1(n2_adj_4965), .I2(n3453), 
            .I3(n28590), .O(color_23__N_164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_8 (.CI(n28590), .I0(n2_adj_4965), .I1(n3453), 
            .CO(n28591));
    SB_LUT4 rem_4_add_2298_7_lut (.I0(n43028), .I1(n2_adj_4965), .I2(n3454), 
            .I3(n28589), .O(color_23__N_164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_7 (.CI(n28589), .I0(n2_adj_4965), .I1(n3454), 
            .CO(n28590));
    SB_LUT4 rem_4_add_2298_6_lut (.I0(n43031), .I1(n2_adj_4965), .I2(n3455), 
            .I3(n28588), .O(color_23__N_164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_6 (.CI(n28588), .I0(n2_adj_4965), .I1(n3455), 
            .CO(n28589));
    SB_LUT4 rem_4_add_2298_5_lut (.I0(n43034), .I1(n2_adj_4965), .I2(n3456), 
            .I3(n28587), .O(color_23__N_164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_5 (.CI(n28587), .I0(n2_adj_4965), .I1(n3456), 
            .CO(n28588));
    SB_LUT4 rem_4_add_2298_4_lut (.I0(n43037), .I1(n2_adj_4965), .I2(n3457), 
            .I3(n28586), .O(color_23__N_164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_4 (.CI(n28586), .I0(n2_adj_4965), .I1(n3457), 
            .CO(n28587));
    SB_LUT4 rem_4_add_2298_3_lut (.I0(communication_counter[1]), .I1(n2_adj_4965), 
            .I2(n3458), .I3(n28585), .O(color_23__N_164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_3 (.CI(n28585), .I0(n2_adj_4965), .I1(n3458), 
            .CO(n28586));
    SB_LUT4 rem_4_add_2298_2_lut (.I0(communication_counter[0]), .I1(n2_adj_4965), 
            .I2(n3459), .I3(VCC_net), .O(color_23__N_164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_2 (.CI(VCC_net), .I0(n2_adj_4965), .I1(n3459), 
            .CO(n28585));
    SB_LUT4 add_5468_7_lut (.I0(GND_net), .I1(n3353), .I2(VCC_net), .I3(n28584), 
            .O(n10082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5468_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5468_6_lut (.I0(GND_net), .I1(n3354), .I2(GND_net), .I3(n28583), 
            .O(n10083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5468_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5468_6 (.CI(n28583), .I0(n3354), .I1(GND_net), .CO(n28584));
    SB_LUT4 add_5468_5_lut (.I0(GND_net), .I1(n3355), .I2(GND_net), .I3(n28582), 
            .O(n10084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5468_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5468_5 (.CI(n28582), .I0(n3355), .I1(GND_net), .CO(n28583));
    SB_LUT4 add_5468_4_lut (.I0(GND_net), .I1(n3356), .I2(VCC_net), .I3(n28581), 
            .O(n10085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5468_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5468_4 (.CI(n28581), .I0(n3356), .I1(VCC_net), .CO(n28582));
    SB_LUT4 add_5468_3_lut (.I0(GND_net), .I1(n3357), .I2(VCC_net), .I3(n28580), 
            .O(n10086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5468_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5468_3 (.CI(n28580), .I0(n3357), .I1(VCC_net), .CO(n28581));
    SB_LUT4 add_5468_2_lut (.I0(GND_net), .I1(n3358), .I2(GND_net), .I3(VCC_net), 
            .O(n10087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5468_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5468_2 (.CI(VCC_net), .I0(n3358), .I1(GND_net), .CO(n28580));
    SB_CARRY rem_4_add_1787_19 (.CI(n28907), .I0(n2642_adj_4491), .I1(VCC_net), 
            .CO(n28908));
    SB_LUT4 add_2273_25_lut (.I0(n249), .I1(n43089), .I2(n248), .I3(n28579), 
            .O(displacement_23__N_229[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2273_24_lut (.I0(n393), .I1(n43089), .I2(n392), .I3(n28578), 
            .O(displacement_23__N_229[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1787_18_lut (.I0(GND_net), .I1(n2643_adj_4490), .I2(VCC_net), 
            .I3(n28906), .O(n2710)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2273_24 (.CI(n28578), .I0(n43089), .I1(n392), .CO(n28579));
    SB_LUT4 add_2273_23_lut (.I0(n534), .I1(n43089), .I2(n533), .I3(n28577), 
            .O(displacement_23__N_229[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1787_18 (.CI(n28906), .I0(n2643_adj_4490), .I1(VCC_net), 
            .CO(n28907));
    SB_CARRY add_2273_23 (.CI(n28577), .I0(n43089), .I1(n533), .CO(n28578));
    SB_LUT4 add_2273_22_lut (.I0(n672), .I1(n43089), .I2(n671), .I3(n28576), 
            .O(displacement_23__N_229[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_22 (.CI(n28576), .I0(n43089), .I1(n671), .CO(n28577));
    SB_LUT4 rem_4_add_1787_17_lut (.I0(GND_net), .I1(n2644), .I2(VCC_net), 
            .I3(n28905), .O(n2711_adj_4484)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2273_21_lut (.I0(n807), .I1(n43089), .I2(n806), .I3(n28575), 
            .O(displacement_23__N_229[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1787_17 (.CI(n28905), .I0(n2644), .I1(VCC_net), 
            .CO(n28906));
    SB_CARRY add_2273_21 (.CI(n28575), .I0(n43089), .I1(n806), .CO(n28576));
    SB_LUT4 add_2273_20_lut (.I0(n939), .I1(n43089), .I2(n938), .I3(n28574), 
            .O(displacement_23__N_229[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12426_3_lut (.I0(gearBoxRatio[12]), .I1(\data_in_frame[18] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17108));   // verilog/coms.v(126[12] 289[6])
    defparam i12426_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12427_3_lut (.I0(gearBoxRatio[13]), .I1(\data_in_frame[18] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17109));   // verilog/coms.v(126[12] 289[6])
    defparam i12427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1658_3_lut_3_lut (.I0(n2471), .I1(n6019), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12428_3_lut (.I0(gearBoxRatio[14]), .I1(\data_in_frame[18] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17110));   // verilog/coms.v(126[12] 289[6])
    defparam i12428_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_916_9_lut (.I0(GND_net), .I1(n1351), .I2(VCC_net), 
            .I3(n27987), .O(n1418_adj_4537)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_16_lut (.I0(GND_net), .I1(n2645), .I2(VCC_net), 
            .I3(n28904), .O(n2712)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_16 (.CI(n28904), .I0(n2645), .I1(VCC_net), 
            .CO(n28905));
    SB_CARRY add_2273_20 (.CI(n28574), .I0(n43089), .I1(n938), .CO(n28575));
    SB_LUT4 add_2273_19_lut (.I0(n1068), .I1(n43089), .I2(n1067), .I3(n28573), 
            .O(displacement_23__N_229[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_19 (.CI(n28573), .I0(n43089), .I1(n1067), .CO(n28574));
    SB_LUT4 i12912_3_lut (.I0(setpoint[21]), .I1(n4313), .I2(n36839), 
            .I3(GND_net), .O(n17594));   // verilog/coms.v(126[12] 289[6])
    defparam i12912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12429_3_lut (.I0(gearBoxRatio[15]), .I1(\data_in_frame[18] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17111));   // verilog/coms.v(126[12] 289[6])
    defparam i12429_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1657_3_lut_3_lut (.I0(n2471), .I1(n6018), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12430_3_lut (.I0(gearBoxRatio[16]), .I1(\data_in_frame[17] [0]), 
            .I2(n36885), .I3(GND_net), .O(n17112));   // verilog/coms.v(126[12] 289[6])
    defparam i12430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1655_3_lut_3_lut (.I0(n2471), .I1(n6016), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12431_3_lut (.I0(gearBoxRatio[17]), .I1(\data_in_frame[17] [1]), 
            .I2(n36885), .I3(GND_net), .O(n17113));   // verilog/coms.v(126[12] 289[6])
    defparam i12431_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2273_18_lut (.I0(n1194), .I1(n43089), .I2(n1193), .I3(n28572), 
            .O(displacement_23__N_229[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_18 (.CI(n28572), .I0(n43089), .I1(n1193), .CO(n28573));
    SB_LUT4 rem_4_add_1787_15_lut (.I0(GND_net), .I1(n2646), .I2(VCC_net), 
            .I3(n28903), .O(n2713_adj_4483)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_15 (.CI(n28903), .I0(n2646), .I1(VCC_net), 
            .CO(n28904));
    SB_LUT4 rem_4_add_1787_14_lut (.I0(GND_net), .I1(n2647), .I2(VCC_net), 
            .I3(n28902), .O(n2714)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2273_17_lut (.I0(n1317), .I1(n43089), .I2(n1316), .I3(n28571), 
            .O(displacement_23__N_229[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i12432_3_lut (.I0(gearBoxRatio[18]), .I1(\data_in_frame[17] [2]), 
            .I2(n36885), .I3(GND_net), .O(n17114));   // verilog/coms.v(126[12] 289[6])
    defparam i12432_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12911_3_lut (.I0(setpoint[20]), .I1(n4312), .I2(n36839), 
            .I3(GND_net), .O(n17593));   // verilog/coms.v(126[12] 289[6])
    defparam i12911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1654_3_lut_3_lut (.I0(n2471), .I1(n6015), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1787_14 (.CI(n28902), .I0(n2647), .I1(VCC_net), 
            .CO(n28903));
    SB_LUT4 rem_4_add_1787_13_lut (.I0(GND_net), .I1(n2648), .I2(VCC_net), 
            .I3(n28901), .O(n2715_adj_4482)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_13 (.CI(n28901), .I0(n2648), .I1(VCC_net), 
            .CO(n28902));
    SB_CARRY add_2273_17 (.CI(n28571), .I0(n43089), .I1(n1316), .CO(n28572));
    SB_LUT4 add_2273_16_lut (.I0(n1437), .I1(n43089), .I2(n1436), .I3(n28570), 
            .O(displacement_23__N_229[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1787_12_lut (.I0(GND_net), .I1(n2649), .I2(VCC_net), 
            .I3(n28900), .O(n2716)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12433_3_lut (.I0(gearBoxRatio[19]), .I1(\data_in_frame[17] [3]), 
            .I2(n36885), .I3(GND_net), .O(n17115));   // verilog/coms.v(126[12] 289[6])
    defparam i12433_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12434_3_lut (.I0(gearBoxRatio[20]), .I1(\data_in_frame[17] [4]), 
            .I2(n36885), .I3(GND_net), .O(n17116));   // verilog/coms.v(126[12] 289[6])
    defparam i12434_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2273_16 (.CI(n28570), .I0(n43089), .I1(n1436), .CO(n28571));
    SB_LUT4 i12435_3_lut (.I0(gearBoxRatio[21]), .I1(\data_in_frame[17] [5]), 
            .I2(n36885), .I3(GND_net), .O(n17117));   // verilog/coms.v(126[12] 289[6])
    defparam i12435_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1787_12 (.CI(n28900), .I0(n2649), .I1(VCC_net), 
            .CO(n28901));
    SB_LUT4 add_2273_15_lut (.I0(n1554), .I1(n43089), .I2(n1553), .I3(n28569), 
            .O(displacement_23__N_229[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_15 (.CI(n28569), .I0(n43089), .I1(n1553), .CO(n28570));
    SB_LUT4 rem_4_add_1787_11_lut (.I0(GND_net), .I1(n2650), .I2(VCC_net), 
            .I3(n28899), .O(n2717_adj_4481)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2273_14_lut (.I0(n1668), .I1(n43089), .I2(n1667), .I3(n28568), 
            .O(displacement_23__N_229[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_14 (.CI(n28568), .I0(n43089), .I1(n1667), .CO(n28569));
    SB_LUT4 add_2273_13_lut (.I0(n1779), .I1(n43089), .I2(n1778), .I3(n28567), 
            .O(displacement_23__N_229[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_13 (.CI(n28567), .I0(n43089), .I1(n1778), .CO(n28568));
    SB_LUT4 add_2273_12_lut (.I0(n1887), .I1(n43089), .I2(n1886), .I3(n28566), 
            .O(displacement_23__N_229[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_12 (.CI(n28566), .I0(n43089), .I1(n1886), .CO(n28567));
    SB_LUT4 add_2273_11_lut (.I0(n1992), .I1(n43089), .I2(n1991), .I3(n28565), 
            .O(displacement_23__N_229[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_11 (.CI(n28565), .I0(n43089), .I1(n1991), .CO(n28566));
    SB_LUT4 add_2273_10_lut (.I0(n2094), .I1(n43089), .I2(n2093), .I3(n28564), 
            .O(displacement_23__N_229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_10 (.CI(n28564), .I0(n43089), .I1(n2093), .CO(n28565));
    SB_LUT4 add_2273_9_lut (.I0(n2193), .I1(n43089), .I2(n2192), .I3(n28563), 
            .O(displacement_23__N_229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_9 (.CI(n28563), .I0(n43089), .I1(n2192), .CO(n28564));
    SB_LUT4 add_2273_8_lut (.I0(n2289), .I1(n43089), .I2(n2288), .I3(n28562), 
            .O(displacement_23__N_229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_8 (.CI(n28562), .I0(n43089), .I1(n2288), .CO(n28563));
    SB_LUT4 add_2273_7_lut (.I0(n2382), .I1(n43089), .I2(n2381), .I3(n28561), 
            .O(displacement_23__N_229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_7 (.CI(n28561), .I0(n43089), .I1(n2381), .CO(n28562));
    SB_LUT4 add_2273_6_lut (.I0(n2472), .I1(n43089), .I2(n2471), .I3(n28560), 
            .O(displacement_23__N_229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_6 (.CI(n28560), .I0(n43089), .I1(n2471), .CO(n28561));
    SB_LUT4 add_2273_5_lut (.I0(n2559), .I1(n43089), .I2(n2558), .I3(n28559), 
            .O(displacement_23__N_229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_5 (.CI(n28559), .I0(n43089), .I1(n2558), .CO(n28560));
    SB_LUT4 add_2273_4_lut (.I0(n2643), .I1(n43089), .I2(n2642), .I3(n28558), 
            .O(displacement_23__N_229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_4 (.CI(n28558), .I0(n43089), .I1(n2642), .CO(n28559));
    SB_LUT4 add_2273_3_lut (.I0(n2724), .I1(n43089), .I2(n2723), .I3(n28557), 
            .O(displacement_23__N_229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2273_3 (.CI(n28557), .I0(n43089), .I1(n2723), .CO(n28558));
    SB_LUT4 add_2273_2_lut (.I0(n2802), .I1(n43089), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2273_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_916_9 (.CI(n27987), .I0(n1351), .I1(VCC_net), .CO(n27988));
    SB_LUT4 rem_4_add_916_8_lut (.I0(GND_net), .I1(n1352), .I2(VCC_net), 
            .I3(n27986), .O(n1419_adj_4538)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2273_2 (.CI(VCC_net), .I0(n43089), .I1(n2801), .CO(n28557));
    SB_CARRY rem_4_add_916_8 (.CI(n27986), .I0(n1352), .I1(VCC_net), .CO(n27987));
    SB_LUT4 rem_4_add_916_7_lut (.I0(GND_net), .I1(n1353), .I2(VCC_net), 
            .I3(n27985), .O(n1420_adj_4539)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_11 (.CI(n28899), .I0(n2650), .I1(VCC_net), 
            .CO(n28900));
    SB_CARRY rem_4_add_916_7 (.CI(n27985), .I0(n1353), .I1(VCC_net), .CO(n27986));
    SB_LUT4 rem_4_add_916_6_lut (.I0(GND_net), .I1(n1354), .I2(GND_net), 
            .I3(n27984), .O(n1421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12436_3_lut (.I0(gearBoxRatio[22]), .I1(\data_in_frame[17] [6]), 
            .I2(n36885), .I3(GND_net), .O(n17118));   // verilog/coms.v(126[12] 289[6])
    defparam i12436_3_lut.LUT_INIT = 16'hacac;
    SB_DFF communication_counter_1176__i1 (.Q(communication_counter[1]), .C(LED_c), 
           .D(n164));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_CARRY rem_4_add_916_6 (.CI(n27984), .I0(n1354), .I1(GND_net), .CO(n27985));
    SB_LUT4 i12437_3_lut (.I0(gearBoxRatio[23]), .I1(\data_in_frame[17] [7]), 
            .I2(n36885), .I3(GND_net), .O(n17119));   // verilog/coms.v(126[12] 289[6])
    defparam i12437_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12438_3_lut (.I0(Kp[1]), .I1(\data_in_frame[2] [1]), .I2(n36885), 
            .I3(GND_net), .O(n17120));   // verilog/coms.v(126[12] 289[6])
    defparam i12438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1787_10_lut (.I0(GND_net), .I1(n2651), .I2(VCC_net), 
            .I3(n28898), .O(n2718)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12439_3_lut (.I0(Kp[2]), .I1(\data_in_frame[2] [2]), .I2(n36885), 
            .I3(GND_net), .O(n17121));   // verilog/coms.v(126[12] 289[6])
    defparam i12439_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1787_10 (.CI(n28898), .I0(n2651), .I1(VCC_net), 
            .CO(n28899));
    SB_LUT4 i12440_3_lut (.I0(Kp[3]), .I1(\data_in_frame[2] [3]), .I2(n36885), 
            .I3(GND_net), .O(n17122));   // verilog/coms.v(126[12] 289[6])
    defparam i12440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2272_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n28556), 
            .O(n6072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12441_3_lut (.I0(Kp[4]), .I1(\data_in_frame[2] [4]), .I2(n36885), 
            .I3(GND_net), .O(n17123));   // verilog/coms.v(126[12] 289[6])
    defparam i12441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1712_3_lut_3_lut (.I0(n2558), .I1(n6038), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12442_3_lut (.I0(Kp[5]), .I1(\data_in_frame[2] [5]), .I2(n36885), 
            .I3(GND_net), .O(n17124));   // verilog/coms.v(126[12] 289[6])
    defparam i12442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12443_3_lut (.I0(Kp[6]), .I1(\data_in_frame[2] [6]), .I2(n36885), 
            .I3(GND_net), .O(n17125));   // verilog/coms.v(126[12] 289[6])
    defparam i12443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1699_3_lut_3_lut (.I0(n2558), .I1(n6025), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12444_3_lut (.I0(Kp[7]), .I1(\data_in_frame[2] [7]), .I2(n36885), 
            .I3(GND_net), .O(n17126));   // verilog/coms.v(126[12] 289[6])
    defparam i12444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12445_3_lut (.I0(Ki[1]), .I1(\data_in_frame[3] [1]), .I2(n36885), 
            .I3(GND_net), .O(n17127));   // verilog/coms.v(126[12] 289[6])
    defparam i12445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2272_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n28555), 
            .O(n6073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_5_lut (.I0(GND_net), .I1(n1355), .I2(GND_net), 
            .I3(n27983), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_24 (.CI(n28555), .I0(n2700), .I1(n79), .CO(n28556));
    SB_LUT4 i12446_3_lut (.I0(Ki[2]), .I1(\data_in_frame[3] [2]), .I2(n36885), 
            .I3(GND_net), .O(n17128));   // verilog/coms.v(126[12] 289[6])
    defparam i12446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2272_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n28554), 
            .O(n6074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4406));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2272_23 (.CI(n28554), .I0(n2701), .I1(n80), .CO(n28555));
    SB_LUT4 add_2272_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n28553), 
            .O(n6075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_22 (.CI(n28553), .I0(n2702), .I1(n81), .CO(n28554));
    SB_LUT4 add_2272_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n28552), 
            .O(n6076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_21 (.CI(n28552), .I0(n2703), .I1(n82), .CO(n28553));
    SB_LUT4 add_2272_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n28551), 
            .O(n6077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_20 (.CI(n28551), .I0(n2704), .I1(n83), .CO(n28552));
    SB_LUT4 add_2272_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n28550), 
            .O(n6078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_19 (.CI(n28550), .I0(n2705), .I1(n84), .CO(n28551));
    SB_LUT4 add_2272_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n28549), 
            .O(n6079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_18 (.CI(n28549), .I0(n2706), .I1(n85), .CO(n28550));
    SB_LUT4 add_2272_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n28548), 
            .O(n6080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_17 (.CI(n28548), .I0(n2707), .I1(n86), .CO(n28549));
    SB_LUT4 add_2272_16_lut (.I0(GND_net), .I1(n2708_adj_4418), .I2(n87), 
            .I3(n28547), .O(n6081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_16 (.CI(n28547), .I0(n2708_adj_4418), .I1(n87), 
            .CO(n28548));
    SB_LUT4 add_2272_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n28546), 
            .O(n6082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_15 (.CI(n28546), .I0(n2709), .I1(n88), .CO(n28547));
    SB_LUT4 add_2272_14_lut (.I0(GND_net), .I1(n2710_adj_4419), .I2(n89), 
            .I3(n28545), .O(n6083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_14 (.CI(n28545), .I0(n2710_adj_4419), .I1(n89), 
            .CO(n28546));
    SB_LUT4 add_2272_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n28544), 
            .O(n6084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_13 (.CI(n28544), .I0(n2711), .I1(n90), .CO(n28545));
    SB_LUT4 add_2272_12_lut (.I0(GND_net), .I1(n2712_adj_4420), .I2(n91), 
            .I3(n28543), .O(n6085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_12 (.CI(n28543), .I0(n2712_adj_4420), .I1(n91), 
            .CO(n28544));
    SB_LUT4 add_2272_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n28542), 
            .O(n6086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_11 (.CI(n28542), .I0(n2713), .I1(n92), .CO(n28543));
    SB_LUT4 add_2272_10_lut (.I0(GND_net), .I1(n2714_adj_4421), .I2(n93), 
            .I3(n28541), .O(n6087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_10 (.CI(n28541), .I0(n2714_adj_4421), .I1(n93), 
            .CO(n28542));
    SB_LUT4 add_2272_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n28540), 
            .O(n6088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_9 (.CI(n28540), .I0(n2715), .I1(n94), .CO(n28541));
    SB_LUT4 add_2272_8_lut (.I0(GND_net), .I1(n2716_adj_4422), .I2(n95), 
            .I3(n28539), .O(n6089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_8 (.CI(n28539), .I0(n2716_adj_4422), .I1(n95), .CO(n28540));
    SB_LUT4 add_2272_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n28538), 
            .O(n6090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_7 (.CI(n28538), .I0(n2717), .I1(n96), .CO(n28539));
    SB_LUT4 add_2272_6_lut (.I0(GND_net), .I1(n2718_adj_4423), .I2(n97), 
            .I3(n28537), .O(n6091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_6 (.CI(n28537), .I0(n2718_adj_4423), .I1(n97), .CO(n28538));
    SB_LUT4 add_2272_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n28536), 
            .O(n6092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_5 (.CI(n28536), .I0(n2719), .I1(n98), .CO(n28537));
    SB_LUT4 add_2272_4_lut (.I0(GND_net), .I1(n2720_adj_4424), .I2(n99), 
            .I3(n28535), .O(n6093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_4 (.CI(n28535), .I0(n2720_adj_4424), .I1(n99), .CO(n28536));
    SB_LUT4 add_2272_3_lut (.I0(GND_net), .I1(n669), .I2(n558), .I3(n28534), 
            .O(n6094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2272_3 (.CI(n28534), .I0(n669), .I1(n558), .CO(n28535));
    SB_CARRY add_2272_2 (.CI(VCC_net), .I0(n670), .I1(VCC_net), .CO(n28534));
    SB_LUT4 add_2271_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n28533), 
            .O(n6048)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2271_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n28532), 
            .O(n6049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_22 (.CI(n28532), .I0(n2619), .I1(n80), .CO(n28533));
    SB_LUT4 add_2271_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n28531), 
            .O(n6050)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_21 (.CI(n28531), .I0(n2620), .I1(n81), .CO(n28532));
    SB_LUT4 add_2271_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n28530), 
            .O(n6051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_20 (.CI(n28530), .I0(n2621), .I1(n82), .CO(n28531));
    SB_LUT4 add_2271_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n28529), 
            .O(n6052)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_19 (.CI(n28529), .I0(n2622), .I1(n83), .CO(n28530));
    SB_LUT4 add_2271_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n28528), 
            .O(n6053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_18 (.CI(n28528), .I0(n2623), .I1(n84), .CO(n28529));
    SB_LUT4 add_2271_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n28527), 
            .O(n6054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_17 (.CI(n28527), .I0(n2624), .I1(n85), .CO(n28528));
    SB_LUT4 add_2271_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n28526), 
            .O(n6055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_16 (.CI(n28526), .I0(n2625), .I1(n86), .CO(n28527));
    SB_LUT4 add_2271_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n28525), 
            .O(n6056)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_15 (.CI(n28525), .I0(n2626), .I1(n87), .CO(n28526));
    SB_LUT4 add_2271_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n28524), 
            .O(n6057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_14 (.CI(n28524), .I0(n2627), .I1(n88), .CO(n28525));
    SB_LUT4 add_2271_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n28523), 
            .O(n6058)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_13 (.CI(n28523), .I0(n2628), .I1(n89), .CO(n28524));
    SB_LUT4 add_2271_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n28522), 
            .O(n6059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_12 (.CI(n28522), .I0(n2629), .I1(n90), .CO(n28523));
    SB_LUT4 add_2271_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n28521), 
            .O(n6060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_11 (.CI(n28521), .I0(n2630), .I1(n91), .CO(n28522));
    SB_LUT4 add_2271_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n28520), 
            .O(n6061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_10 (.CI(n28520), .I0(n2631), .I1(n92), .CO(n28521));
    SB_LUT4 add_2271_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n28519), 
            .O(n6062)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_9 (.CI(n28519), .I0(n2632), .I1(n93), .CO(n28520));
    SB_LUT4 add_2271_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n28518), 
            .O(n6063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_8 (.CI(n28518), .I0(n2633), .I1(n94), .CO(n28519));
    SB_LUT4 add_2271_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n28517), 
            .O(n6064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_7 (.CI(n28517), .I0(n2634), .I1(n95), .CO(n28518));
    SB_LUT4 add_2271_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n28516), 
            .O(n6065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_6 (.CI(n28516), .I0(n2635), .I1(n96), .CO(n28517));
    SB_LUT4 add_2271_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n28515), 
            .O(n6066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_5 (.CI(n28515), .I0(n2636), .I1(n97), .CO(n28516));
    SB_LUT4 add_2271_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n28514), 
            .O(n6067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_4 (.CI(n28514), .I0(n2637), .I1(n98), .CO(n28515));
    SB_LUT4 add_2271_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n28513), 
            .O(n6068)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_3 (.CI(n28513), .I0(n2638), .I1(n99), .CO(n28514));
    SB_LUT4 add_2271_2_lut (.I0(GND_net), .I1(n668), .I2(n558), .I3(VCC_net), 
            .O(n6069)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2271_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2271_2 (.CI(VCC_net), .I0(n668), .I1(n558), .CO(n28513));
    SB_LUT4 add_2270_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n28512), 
            .O(n6025)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2270_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n28511), 
            .O(n6026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_21 (.CI(n28511), .I0(n2535), .I1(n81), .CO(n28512));
    SB_LUT4 add_2270_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n28510), 
            .O(n6027)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_20 (.CI(n28510), .I0(n2536), .I1(n82), .CO(n28511));
    SB_LUT4 add_2270_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n28509), 
            .O(n6028)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_19 (.CI(n28509), .I0(n2537), .I1(n83), .CO(n28510));
    SB_LUT4 add_2270_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n28508), 
            .O(n6029)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_18 (.CI(n28508), .I0(n2538), .I1(n84), .CO(n28509));
    SB_LUT4 rem_4_add_1787_9_lut (.I0(GND_net), .I1(n2652), .I2(VCC_net), 
            .I3(n28897), .O(n2719_adj_4480)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2270_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n28507), 
            .O(n6030)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_17 (.CI(n28507), .I0(n2539), .I1(n85), .CO(n28508));
    SB_LUT4 add_2270_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n28506), 
            .O(n6031)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_16 (.CI(n28506), .I0(n2540), .I1(n86), .CO(n28507));
    SB_LUT4 add_2270_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n28505), 
            .O(n6032)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_15 (.CI(n28505), .I0(n2541), .I1(n87), .CO(n28506));
    SB_CARRY rem_4_add_1787_9 (.CI(n28897), .I0(n2652), .I1(VCC_net), 
            .CO(n28898));
    SB_LUT4 add_2270_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n28504), 
            .O(n6033)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_14 (.CI(n28504), .I0(n2542), .I1(n88), .CO(n28505));
    SB_LUT4 add_2270_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n28503), 
            .O(n6034)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_5 (.CI(n27983), .I0(n1355), .I1(GND_net), .CO(n27984));
    SB_CARRY add_2270_13 (.CI(n28503), .I0(n2543), .I1(n89), .CO(n28504));
    SB_LUT4 rem_4_add_1787_8_lut (.I0(GND_net), .I1(n2653), .I2(VCC_net), 
            .I3(n28896), .O(n2720)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2270_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n28502), 
            .O(n6035)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_12 (.CI(n28502), .I0(n2544), .I1(n90), .CO(n28503));
    SB_LUT4 add_2270_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n28501), 
            .O(n6036)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_11 (.CI(n28501), .I0(n2545), .I1(n91), .CO(n28502));
    SB_LUT4 div_46_i1700_3_lut_3_lut (.I0(n2558), .I1(n6026), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2270_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n28500), 
            .O(n6037)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1702_3_lut_3_lut (.I0(n2558), .I1(n6028), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1787_8 (.CI(n28896), .I0(n2653), .I1(VCC_net), 
            .CO(n28897));
    SB_CARRY add_2270_10 (.CI(n28500), .I0(n2546), .I1(n92), .CO(n28501));
    SB_LUT4 add_2270_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n28499), 
            .O(n6038)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_9 (.CI(n28499), .I0(n2547), .I1(n93), .CO(n28500));
    SB_LUT4 rem_4_add_1787_7_lut (.I0(GND_net), .I1(n2654), .I2(GND_net), 
            .I3(n28895), .O(n2721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2270_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n28498), 
            .O(n6039)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1701_3_lut_3_lut (.I0(n2558), .I1(n6027), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2270_8 (.CI(n28498), .I0(n2548), .I1(n94), .CO(n28499));
    SB_CARRY rem_4_add_1787_7 (.CI(n28895), .I0(n2654), .I1(GND_net), 
            .CO(n28896));
    SB_LUT4 add_2270_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n28497), 
            .O(n6040)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_6_lut (.I0(GND_net), .I1(n2655), .I2(GND_net), 
            .I3(n28894), .O(n2722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_7 (.CI(n28497), .I0(n2549), .I1(n95), .CO(n28498));
    SB_LUT4 add_2270_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n28496), 
            .O(n6041)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_4_lut (.I0(GND_net), .I1(n1356), .I2(VCC_net), 
            .I3(n27982), .O(n1423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_6 (.CI(n28894), .I0(n2655), .I1(GND_net), 
            .CO(n28895));
    SB_CARRY add_2270_6 (.CI(n28496), .I0(n2550), .I1(n96), .CO(n28497));
    SB_LUT4 add_2270_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n28495), 
            .O(n6042)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_5 (.CI(n28495), .I0(n2551), .I1(n97), .CO(n28496));
    SB_LUT4 add_2270_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n28494), 
            .O(n6043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_5_lut (.I0(GND_net), .I1(n2656), .I2(VCC_net), 
            .I3(n28893), .O(n2723_adj_4479)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_4 (.CI(n28494), .I0(n2552), .I1(n98), .CO(n28495));
    SB_CARRY rem_4_add_1787_5 (.CI(n28893), .I0(n2656), .I1(VCC_net), 
            .CO(n28894));
    SB_LUT4 add_2270_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n28493), 
            .O(n6044)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12447_3_lut (.I0(Ki[3]), .I1(\data_in_frame[3] [3]), .I2(n36885), 
            .I3(GND_net), .O(n17129));   // verilog/coms.v(126[12] 289[6])
    defparam i12447_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_916_4 (.CI(n27982), .I0(n1356), .I1(VCC_net), .CO(n27983));
    SB_LUT4 rem_4_add_1787_4_lut (.I0(GND_net), .I1(n2657), .I2(VCC_net), 
            .I3(n28892), .O(n2724_adj_4478)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2270_3 (.CI(n28493), .I0(n2553), .I1(n99), .CO(n28494));
    SB_LUT4 rem_4_add_916_3_lut (.I0(GND_net), .I1(n1357), .I2(VCC_net), 
            .I3(n27981), .O(n1424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_4 (.CI(n28892), .I0(n2657), .I1(VCC_net), 
            .CO(n28893));
    SB_LUT4 add_2270_2_lut (.I0(GND_net), .I1(n667), .I2(n558), .I3(VCC_net), 
            .O(n6045)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2270_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_3 (.CI(n27981), .I0(n1357), .I1(VCC_net), .CO(n27982));
    SB_LUT4 rem_4_add_1787_3_lut (.I0(GND_net), .I1(n2658), .I2(GND_net), 
            .I3(n28891), .O(n2725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_3 (.CI(n28891), .I0(n2658), .I1(GND_net), 
            .CO(n28892));
    SB_CARRY add_2270_2 (.CI(VCC_net), .I0(n667), .I1(n558), .CO(n28493));
    SB_LUT4 add_2269_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n28492), 
            .O(n6003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1719_3_lut_3_lut (.I0(n2558), .I1(n6045), .I2(n667), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_916_2_lut (.I0(GND_net), .I1(n1358), .I2(GND_net), 
            .I3(VCC_net), .O(n1425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_2 (.CI(VCC_net), .I0(n2758), .I1(VCC_net), 
            .CO(n28891));
    SB_LUT4 rem_4_add_1854_26_lut (.I0(n2768), .I1(n2735), .I2(VCC_net), 
            .I3(n28890), .O(n2834)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2269_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n28491), 
            .O(n6004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_20 (.CI(n28491), .I0(n2448), .I1(n82), .CO(n28492));
    SB_LUT4 add_2269_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n28490), 
            .O(n6005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_19 (.CI(n28490), .I0(n2449), .I1(n83), .CO(n28491));
    SB_LUT4 add_2269_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n28489), 
            .O(n6006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_18 (.CI(n28489), .I0(n2450), .I1(n84), .CO(n28490));
    SB_LUT4 add_2269_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n28488), 
            .O(n6007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_17 (.CI(n28488), .I0(n2451), .I1(n85), .CO(n28489));
    SB_LUT4 add_2269_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n28487), 
            .O(n6008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_16 (.CI(n28487), .I0(n2452), .I1(n86), .CO(n28488));
    SB_LUT4 add_2269_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n28486), 
            .O(n6009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_15 (.CI(n28486), .I0(n2453), .I1(n87), .CO(n28487));
    SB_LUT4 add_2269_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n28485), 
            .O(n6010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_14 (.CI(n28485), .I0(n2454), .I1(n88), .CO(n28486));
    SB_LUT4 add_2269_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n28484), 
            .O(n6011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_13 (.CI(n28484), .I0(n2455), .I1(n89), .CO(n28485));
    SB_LUT4 add_2269_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n28483), 
            .O(n6012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_12 (.CI(n28483), .I0(n2456), .I1(n90), .CO(n28484));
    SB_LUT4 add_2269_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n28482), 
            .O(n6013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_11 (.CI(n28482), .I0(n2457), .I1(n91), .CO(n28483));
    SB_LUT4 add_2269_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n28481), 
            .O(n6014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_10 (.CI(n28481), .I0(n2458), .I1(n92), .CO(n28482));
    SB_LUT4 add_2269_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n28480), 
            .O(n6015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_9 (.CI(n28480), .I0(n2459), .I1(n93), .CO(n28481));
    SB_LUT4 add_2269_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n28479), 
            .O(n6016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_8 (.CI(n28479), .I0(n2460), .I1(n94), .CO(n28480));
    SB_LUT4 add_2269_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n28478), 
            .O(n6017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_7 (.CI(n28478), .I0(n2461), .I1(n95), .CO(n28479));
    SB_LUT4 add_2269_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n28477), 
            .O(n6018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_6 (.CI(n28477), .I0(n2462), .I1(n96), .CO(n28478));
    SB_LUT4 add_2269_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n28476), 
            .O(n6019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_5 (.CI(n28476), .I0(n2463), .I1(n97), .CO(n28477));
    SB_LUT4 add_2269_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n28475), 
            .O(n6020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_4 (.CI(n28475), .I0(n2464), .I1(n98), .CO(n28476));
    SB_LUT4 add_2269_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n28474), 
            .O(n6021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_3 (.CI(n28474), .I0(n2465), .I1(n99), .CO(n28475));
    SB_LUT4 add_2269_2_lut (.I0(GND_net), .I1(n666), .I2(n558), .I3(VCC_net), 
            .O(n6022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2269_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2269_2 (.CI(VCC_net), .I0(n666), .I1(n558), .CO(n28474));
    SB_LUT4 add_2268_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n28473), 
            .O(n5982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2268_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n28472), 
            .O(n5983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_19 (.CI(n28472), .I0(n2358), .I1(n83), .CO(n28473));
    SB_LUT4 add_2268_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n28471), 
            .O(n5984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_18 (.CI(n28471), .I0(n2359), .I1(n84), .CO(n28472));
    SB_LUT4 add_2268_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n28470), 
            .O(n5985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_17 (.CI(n28470), .I0(n2360), .I1(n85), .CO(n28471));
    SB_LUT4 add_2268_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n28469), 
            .O(n5986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_16 (.CI(n28469), .I0(n2361), .I1(n86), .CO(n28470));
    SB_LUT4 add_2268_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n28468), 
            .O(n5987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_15 (.CI(n28468), .I0(n2362), .I1(n87), .CO(n28469));
    SB_LUT4 add_2268_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n28467), 
            .O(n5988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_14 (.CI(n28467), .I0(n2363), .I1(n88), .CO(n28468));
    SB_LUT4 add_2268_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n28466), 
            .O(n5989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_13 (.CI(n28466), .I0(n2364), .I1(n89), .CO(n28467));
    SB_LUT4 add_2268_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n28465), 
            .O(n5990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_12 (.CI(n28465), .I0(n2365), .I1(n90), .CO(n28466));
    SB_LUT4 add_2268_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n28464), 
            .O(n5991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_11 (.CI(n28464), .I0(n2366), .I1(n91), .CO(n28465));
    SB_LUT4 add_2268_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n28463), 
            .O(n5992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_10 (.CI(n28463), .I0(n2367), .I1(n92), .CO(n28464));
    SB_LUT4 add_2268_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n28462), 
            .O(n5993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_9 (.CI(n28462), .I0(n2368), .I1(n93), .CO(n28463));
    SB_LUT4 add_2268_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n28461), 
            .O(n5994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_8 (.CI(n28461), .I0(n2369), .I1(n94), .CO(n28462));
    SB_LUT4 add_2268_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n28460), 
            .O(n5995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_7 (.CI(n28460), .I0(n2370), .I1(n95), .CO(n28461));
    SB_LUT4 add_2268_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n28459), 
            .O(n5996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_6 (.CI(n28459), .I0(n2371), .I1(n96), .CO(n28460));
    SB_LUT4 add_2268_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n28458), 
            .O(n5997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_5 (.CI(n28458), .I0(n2372), .I1(n97), .CO(n28459));
    SB_LUT4 add_2268_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n28457), 
            .O(n5998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_4 (.CI(n28457), .I0(n2373), .I1(n98), .CO(n28458));
    SB_LUT4 add_2268_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n28456), 
            .O(n5999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_3 (.CI(n28456), .I0(n2374), .I1(n99), .CO(n28457));
    SB_LUT4 add_2268_2_lut (.I0(GND_net), .I1(n665), .I2(n558), .I3(VCC_net), 
            .O(n6000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2268_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2268_2 (.CI(VCC_net), .I0(n665), .I1(n558), .CO(n28456));
    SB_LUT4 add_2267_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n28455), 
            .O(n5962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2267_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n28454), 
            .O(n5963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_18 (.CI(n28454), .I0(n2265), .I1(n84), .CO(n28455));
    SB_LUT4 add_2267_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n28453), 
            .O(n5964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_17 (.CI(n28453), .I0(n2266), .I1(n85), .CO(n28454));
    SB_LUT4 add_2267_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n28452), 
            .O(n5965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_16 (.CI(n28452), .I0(n2267), .I1(n86), .CO(n28453));
    SB_LUT4 add_2267_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n28451), 
            .O(n5966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_15 (.CI(n28451), .I0(n2268), .I1(n87), .CO(n28452));
    SB_LUT4 add_2267_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n28450), 
            .O(n5967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_14 (.CI(n28450), .I0(n2269), .I1(n88), .CO(n28451));
    SB_LUT4 add_2267_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n28449), 
            .O(n5968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_13 (.CI(n28449), .I0(n2270), .I1(n89), .CO(n28450));
    SB_LUT4 add_2267_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n28448), 
            .O(n5969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_12 (.CI(n28448), .I0(n2271), .I1(n90), .CO(n28449));
    SB_LUT4 add_2267_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n28447), 
            .O(n5970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_11 (.CI(n28447), .I0(n2272), .I1(n91), .CO(n28448));
    SB_LUT4 add_2267_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n28446), 
            .O(n5971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_10 (.CI(n28446), .I0(n2273), .I1(n92), .CO(n28447));
    SB_LUT4 add_2267_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n28445), 
            .O(n5972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_9 (.CI(n28445), .I0(n2274), .I1(n93), .CO(n28446));
    SB_LUT4 add_2267_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n28444), 
            .O(n5973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_8 (.CI(n28444), .I0(n2275), .I1(n94), .CO(n28445));
    SB_LUT4 add_2267_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n28443), 
            .O(n5974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_7 (.CI(n28443), .I0(n2276), .I1(n95), .CO(n28444));
    SB_LUT4 add_2267_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n28442), 
            .O(n5975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_6 (.CI(n28442), .I0(n2277), .I1(n96), .CO(n28443));
    SB_LUT4 add_2267_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n28441), 
            .O(n5976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_5 (.CI(n28441), .I0(n2278), .I1(n97), .CO(n28442));
    SB_LUT4 add_2267_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n28440), 
            .O(n5977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_4 (.CI(n28440), .I0(n2279), .I1(n98), .CO(n28441));
    SB_LUT4 rem_4_i651_3_lut (.I0(n954), .I1(n1021), .I2(n986), .I3(GND_net), 
            .O(n1053));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2267_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n28439), 
            .O(n5978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_3 (.CI(n28439), .I0(n2280), .I1(n99), .CO(n28440));
    SB_LUT4 add_2267_2_lut (.I0(GND_net), .I1(n664), .I2(n558), .I3(VCC_net), 
            .O(n5979)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2267_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2267_2 (.CI(VCC_net), .I0(n664), .I1(n558), .CO(n28439));
    SB_LUT4 add_2266_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n28438), 
            .O(n5943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2266_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n28437), 
            .O(n5944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_17 (.CI(n28437), .I0(n2169), .I1(n85), .CO(n28438));
    SB_LUT4 add_2266_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n28436), 
            .O(n5945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_16 (.CI(n28436), .I0(n2170), .I1(n86), .CO(n28437));
    SB_LUT4 add_2266_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n28435), 
            .O(n5946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_15 (.CI(n28435), .I0(n2171), .I1(n87), .CO(n28436));
    SB_LUT4 add_2266_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n28434), 
            .O(n5947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_14 (.CI(n28434), .I0(n2172), .I1(n88), .CO(n28435));
    SB_LUT4 add_2266_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n28433), 
            .O(n5948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_13 (.CI(n28433), .I0(n2173), .I1(n89), .CO(n28434));
    SB_LUT4 add_2266_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n28432), 
            .O(n5949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_12 (.CI(n28432), .I0(n2174), .I1(n90), .CO(n28433));
    SB_LUT4 add_2266_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n28431), 
            .O(n5950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_11 (.CI(n28431), .I0(n2175), .I1(n91), .CO(n28432));
    SB_LUT4 add_2266_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n28430), 
            .O(n5951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_10 (.CI(n28430), .I0(n2176), .I1(n92), .CO(n28431));
    SB_LUT4 add_2266_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n28429), 
            .O(n5952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_9 (.CI(n28429), .I0(n2177), .I1(n93), .CO(n28430));
    SB_LUT4 add_2266_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n28428), 
            .O(n5953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_8 (.CI(n28428), .I0(n2178), .I1(n94), .CO(n28429));
    SB_LUT4 add_2266_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n28427), 
            .O(n5954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_7 (.CI(n28427), .I0(n2179), .I1(n95), .CO(n28428));
    SB_LUT4 div_46_i1705_3_lut_3_lut (.I0(n2558), .I1(n6031), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12448_3_lut (.I0(Ki[4]), .I1(\data_in_frame[3] [4]), .I2(n36885), 
            .I3(GND_net), .O(n17130));   // verilog/coms.v(126[12] 289[6])
    defparam i12448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1706_3_lut_3_lut (.I0(n2558), .I1(n6032), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1708_3_lut_3_lut (.I0(n2558), .I1(n6034), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1709_3_lut_3_lut (.I0(n2558), .I1(n6035), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12914_3_lut (.I0(setpoint[23]), .I1(n4315), .I2(n36839), 
            .I3(GND_net), .O(n17596));   // verilog/coms.v(126[12] 289[6])
    defparam i12914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12449_3_lut (.I0(Ki[5]), .I1(\data_in_frame[3] [5]), .I2(n36885), 
            .I3(GND_net), .O(n17131));   // verilog/coms.v(126[12] 289[6])
    defparam i12449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12450_3_lut (.I0(Ki[6]), .I1(\data_in_frame[3] [6]), .I2(n36885), 
            .I3(GND_net), .O(n17132));   // verilog/coms.v(126[12] 289[6])
    defparam i12450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1710_3_lut_3_lut (.I0(n2558), .I1(n6036), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1854_25_lut (.I0(GND_net), .I1(n2736), .I2(VCC_net), 
            .I3(n28889), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_2 (.CI(VCC_net), .I0(n1358), .I1(GND_net), 
            .CO(n27981));
    SB_LUT4 i12451_3_lut (.I0(Ki[7]), .I1(\data_in_frame[3] [7]), .I2(n36885), 
            .I3(GND_net), .O(n17133));   // verilog/coms.v(126[12] 289[6])
    defparam i12451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12452_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17134));   // verilog/coms.v(126[12] 289[6])
    defparam i12452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4405));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2266_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n28426), 
            .O(n5955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_25 (.CI(n28889), .I0(n2736), .I1(VCC_net), 
            .CO(n28890));
    SB_LUT4 unary_minus_28_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4334));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1711_3_lut_3_lut (.I0(n2558), .I1(n6037), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12453_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17135));   // verilog/coms.v(126[12] 289[6])
    defparam i12453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12454_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17136));   // verilog/coms.v(126[12] 289[6])
    defparam i12454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12455_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17137));   // verilog/coms.v(126[12] 289[6])
    defparam i12455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1703_3_lut_3_lut (.I0(n2558), .I1(n6029), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2266_6 (.CI(n28426), .I0(n2180), .I1(n96), .CO(n28427));
    SB_LUT4 div_46_i1717_3_lut_3_lut (.I0(n2558), .I1(n6043), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4404));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12456_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17138));   // verilog/coms.v(126[12] 289[6])
    defparam i12456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12457_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17139));   // verilog/coms.v(126[12] 289[6])
    defparam i12457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12459_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17141));   // verilog/coms.v(126[12] 289[6])
    defparam i12459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12460_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17142));   // verilog/coms.v(126[12] 289[6])
    defparam i12460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12461_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17143));   // verilog/coms.v(126[12] 289[6])
    defparam i12461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12462_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17144));   // verilog/coms.v(126[12] 289[6])
    defparam i12462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1716_3_lut_3_lut (.I0(n2558), .I1(n6042), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12463_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17145));   // verilog/coms.v(126[12] 289[6])
    defparam i12463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4333));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4403));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1715_3_lut_3_lut (.I0(n2558), .I1(n6041), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4402));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4332));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12464_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17146));   // verilog/coms.v(126[12] 289[6])
    defparam i12464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1713_3_lut_3_lut (.I0(n2558), .I1(n6039), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1854_24_lut (.I0(GND_net), .I1(n2737), .I2(VCC_net), 
            .I3(n28888), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12465_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17147));   // verilog/coms.v(126[12] 289[6])
    defparam i12465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1707_3_lut_3_lut (.I0(n2558), .I1(n6033), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12467_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17149));   // verilog/coms.v(126[12] 289[6])
    defparam i12467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12469_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17151));   // verilog/coms.v(126[12] 289[6])
    defparam i12469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4401));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1718_3_lut_3_lut (.I0(n2558), .I1(n6044), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12471_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17153));   // verilog/coms.v(126[12] 289[6])
    defparam i12471_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_24 (.CI(n28888), .I0(n2737), .I1(VCC_net), 
            .CO(n28889));
    SB_LUT4 i12472_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17154));   // verilog/coms.v(126[12] 289[6])
    defparam i12472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12473_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17155));   // verilog/coms.v(126[12] 289[6])
    defparam i12473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12475_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17157));   // verilog/coms.v(126[12] 289[6])
    defparam i12475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2266_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n28425), 
            .O(n5956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12476_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17158));   // verilog/coms.v(126[12] 289[6])
    defparam i12476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1704_3_lut_3_lut (.I0(n2558), .I1(n6030), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2266_5 (.CI(n28425), .I0(n2181), .I1(n97), .CO(n28426));
    SB_LUT4 rem_4_add_782_9_lut (.I0(n1184), .I1(n1151), .I2(VCC_net), 
            .I3(n27980), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1694 (.I0(n1156), .I1(n1158), .I2(GND_net), .I3(GND_net), 
            .O(n37554));
    defparam i1_2_lut_adj_1694.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n1154), .I1(n37554), .I2(n1155), .I3(n1157), 
            .O(n35530));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'ha080;
    SB_LUT4 i3_4_lut_adj_1696 (.I0(n35530), .I1(n1152), .I2(n1151), .I3(n1153), 
            .O(n1184));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i718_3_lut (.I0(n1053), .I1(n1120), .I2(n1085), .I3(GND_net), 
            .O(n1152));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1697 (.I0(n1256), .I1(n1257), .I2(n1258), .I3(GND_net), 
            .O(n35528));
    defparam i1_3_lut_adj_1697.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_i1714_3_lut_3_lut (.I0(n2558), .I1(n6040), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1854_23_lut (.I0(GND_net), .I1(n2738), .I2(VCC_net), 
            .I3(n28887), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n1254), .I1(n1250), .I2(n35528), .I3(n1255), 
            .O(n6_adj_4368));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1699 (.I0(n1251), .I1(n1253), .I2(n1252), .I3(n6_adj_4368), 
            .O(n1283));
    defparam i4_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i785_3_lut (.I0(n1152), .I1(n1219), .I2(n1184), .I3(GND_net), 
            .O(n1251));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1700 (.I0(n1356), .I1(n1357), .I2(n1358), .I3(GND_net), 
            .O(n35524));
    defparam i1_3_lut_adj_1700.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1701 (.I0(n1351), .I1(n1354), .I2(n35524), .I3(n1355), 
            .O(n8_adj_5002));
    defparam i2_4_lut_adj_1701.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1702 (.I0(n1350), .I1(n1349), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_5003));
    defparam i1_2_lut_adj_1702.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1703 (.I0(n1352), .I1(n7_adj_5003), .I2(n1353), 
            .I3(n8_adj_5002), .O(n1382));
    defparam i5_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i852_3_lut (.I0(n1251), .I1(n1318), .I2(n1283), .I3(GND_net), 
            .O(n1350));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1704 (.I0(n1456), .I1(n1458), .I2(GND_net), .I3(GND_net), 
            .O(n37686));
    defparam i1_2_lut_adj_1704.LUT_INIT = 16'heeee;
    SB_LUT4 i12913_3_lut (.I0(setpoint[22]), .I1(n4314), .I2(n36839), 
            .I3(GND_net), .O(n17595));   // verilog/coms.v(126[12] 289[6])
    defparam i12913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n1454), .I1(n37686), .I2(n1455), .I3(n1457), 
            .O(n35558));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'ha080;
    SB_LUT4 i5_4_lut_adj_1706 (.I0(n35558), .I1(n1451), .I2(n1450), .I3(n1452), 
            .O(n12_adj_4924));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1707 (.I0(n1453), .I1(n12_adj_4924), .I2(n1449), 
            .I3(n1448), .O(n1481));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i6_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i919_3_lut (.I0(n1350), .I1(n1417_adj_4536), .I2(n1382), 
            .I3(GND_net), .O(n1449));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1708 (.I0(n1556), .I1(n1557), .I2(n1558), .I3(GND_net), 
            .O(n35555));
    defparam i1_3_lut_adj_1708.LUT_INIT = 16'hfefe;
    SB_LUT4 i22_3_lut_adj_1709 (.I0(bit_ctr[18]), .I1(n40173), .I2(n4385), 
            .I3(GND_net), .O(n33327));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1709.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1710 (.I0(n1554_adj_4534), .I1(n1551), .I2(n35555), 
            .I3(n1555), .O(n11_adj_4919));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut_adj_1710.LUT_INIT = 16'heccc;
    SB_CARRY rem_4_add_1854_23 (.CI(n28887), .I0(n2738), .I1(VCC_net), 
            .CO(n28888));
    SB_LUT4 i5_4_lut_adj_1711 (.I0(n1548), .I1(n1549), .I2(n1547), .I3(n1550), 
            .O(n13_adj_4918));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i5_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1712 (.I0(n13_adj_4918), .I1(n11_adj_4919), .I2(n1553_adj_4533), 
            .I3(n1552), .O(n1580));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i986_3_lut (.I0(n1449), .I1(n1516), .I2(n1481), .I3(GND_net), 
            .O(n1548));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1713 (.I0(n1647_adj_4526), .I1(n1646_adj_4525), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4503));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1713.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1714 (.I0(n1656), .I1(n1657), .I2(n1658), .I3(GND_net), 
            .O(n35572));
    defparam i1_3_lut_adj_1714.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1715 (.I0(n1653_adj_4532), .I1(n1652_adj_4531), 
            .I2(n1651_adj_4530), .I3(n10_adj_4503), .O(n16_adj_4499));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i7_4_lut_adj_1715.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1716 (.I0(n1648_adj_4527), .I1(n1654), .I2(n35572), 
            .I3(n1655), .O(n11_adj_4501));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i2_4_lut_adj_1716.LUT_INIT = 16'heaaa;
    SB_LUT4 add_2266_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n28424), 
            .O(n5957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_4 (.CI(n28424), .I0(n2182), .I1(n98), .CO(n28425));
    SB_LUT4 add_2266_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n28423), 
            .O(n5958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_3 (.CI(n28423), .I0(n2183), .I1(n99), .CO(n28424));
    SB_LUT4 i8_4_lut_adj_1717 (.I0(n11_adj_4501), .I1(n16_adj_4499), .I2(n1649_adj_4528), 
            .I3(n1650_adj_4529), .O(n1679));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i8_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2266_2_lut (.I0(GND_net), .I1(n663), .I2(n558), .I3(VCC_net), 
            .O(n5959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2266_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2266_2 (.CI(VCC_net), .I0(n663), .I1(n558), .CO(n28423));
    SB_LUT4 add_2265_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n28422), 
            .O(n5925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2265_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n28421), 
            .O(n5926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_22_lut (.I0(GND_net), .I1(n2739), .I2(VCC_net), 
            .I3(n28886), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_16 (.CI(n28421), .I0(n2070), .I1(n86), .CO(n28422));
    SB_LUT4 add_2265_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n28420), 
            .O(n5927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_15 (.CI(n28420), .I0(n2071), .I1(n87), .CO(n28421));
    SB_CARRY rem_4_add_1854_22 (.CI(n28886), .I0(n2739), .I1(VCC_net), 
            .CO(n28887));
    SB_LUT4 add_2265_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n28419), 
            .O(n5928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_14 (.CI(n28419), .I0(n2072), .I1(n88), .CO(n28420));
    SB_LUT4 div_46_i1769_3_lut_3_lut (.I0(n2642), .I1(n6063), .I2(n2633), 
            .I3(GND_net), .O(n2714_adj_4421));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2265_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n28418), 
            .O(n5929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_13 (.CI(n28418), .I0(n2073), .I1(n89), .CO(n28419));
    SB_LUT4 rem_4_add_782_8_lut (.I0(GND_net), .I1(n1152), .I2(VCC_net), 
            .I3(n27979), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2265_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n28417), 
            .O(n5930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_12 (.CI(n28417), .I0(n2074), .I1(n90), .CO(n28418));
    SB_LUT4 i12915_3_lut (.I0(quadA_debounced_adj_4372), .I1(reg_B_adj_5064[1]), 
            .I2(n36606), .I3(GND_net), .O(n17597));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1754_3_lut_3_lut (.I0(n2642), .I1(n6048), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1756_3_lut_3_lut (.I0(n2642), .I1(n6050), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1757_3_lut_3_lut (.I0(n2642), .I1(n6051), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1755_3_lut_3_lut (.I0(n2642), .I1(n6049), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1854_21_lut (.I0(GND_net), .I1(n2740), .I2(VCC_net), 
            .I3(n28885), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_21 (.CI(n28885), .I0(n2740), .I1(VCC_net), 
            .CO(n28886));
    SB_LUT4 add_2265_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n28416), 
            .O(n5931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_11 (.CI(n28416), .I0(n2075), .I1(n91), .CO(n28417));
    SB_LUT4 add_2265_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n28415), 
            .O(n5932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_10 (.CI(n28415), .I0(n2076), .I1(n92), .CO(n28416));
    SB_LUT4 add_2265_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n28414), 
            .O(n5933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_9 (.CI(n28414), .I0(n2077), .I1(n93), .CO(n28415));
    SB_LUT4 add_2265_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n28413), 
            .O(n5934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_8 (.CI(n28413), .I0(n2078), .I1(n94), .CO(n28414));
    SB_LUT4 add_2265_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n28412), 
            .O(n5935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF communication_counter_1176__i2 (.Q(communication_counter[2]), .C(LED_c), 
           .D(n163));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_CARRY add_2265_7 (.CI(n28412), .I0(n2079), .I1(n95), .CO(n28413));
    SB_LUT4 rem_4_add_1854_20_lut (.I0(GND_net), .I1(n2741), .I2(VCC_net), 
            .I3(n28884), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_20 (.CI(n28884), .I0(n2741), .I1(VCC_net), 
            .CO(n28885));
    SB_LUT4 div_46_i1758_3_lut_3_lut (.I0(n2642), .I1(n6052), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2265_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n28411), 
            .O(n5936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_19_lut (.I0(GND_net), .I1(n2742), .I2(VCC_net), 
            .I3(n28883), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_6 (.CI(n28411), .I0(n2080), .I1(n96), .CO(n28412));
    SB_LUT4 add_2265_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n28410), 
            .O(n5937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_19 (.CI(n28883), .I0(n2742), .I1(VCC_net), 
            .CO(n28884));
    SB_LUT4 div_46_i1761_3_lut_3_lut (.I0(n2642), .I1(n6055), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1854_18_lut (.I0(GND_net), .I1(n2743), .I2(VCC_net), 
            .I3(n28882), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_18 (.CI(n28882), .I0(n2743), .I1(VCC_net), 
            .CO(n28883));
    SB_CARRY add_2265_5 (.CI(n28410), .I0(n2081), .I1(n97), .CO(n28411));
    SB_LUT4 rem_4_add_1854_17_lut (.I0(GND_net), .I1(n2744), .I2(VCC_net), 
            .I3(n28881), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_8 (.CI(n27979), .I0(n1152), .I1(VCC_net), .CO(n27980));
    SB_CARRY rem_4_add_1854_17 (.CI(n28881), .I0(n2744), .I1(VCC_net), 
            .CO(n28882));
    SB_LUT4 rem_4_add_1854_16_lut (.I0(GND_net), .I1(n2745), .I2(VCC_net), 
            .I3(n28880), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_16 (.CI(n28880), .I0(n2745), .I1(VCC_net), 
            .CO(n28881));
    SB_LUT4 div_46_i1762_3_lut_3_lut (.I0(n2642), .I1(n6056), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2265_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n28409), 
            .O(n5938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_15_lut (.I0(GND_net), .I1(n2746), .I2(VCC_net), 
            .I3(n28879), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_7_lut (.I0(GND_net), .I1(n1153), .I2(VCC_net), 
            .I3(n27978), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_4 (.CI(n28409), .I0(n2082), .I1(n98), .CO(n28410));
    SB_CARRY rem_4_add_1854_15 (.CI(n28879), .I0(n2746), .I1(VCC_net), 
            .CO(n28880));
    SB_LUT4 rem_4_add_1854_14_lut (.I0(GND_net), .I1(n2747), .I2(VCC_net), 
            .I3(n28878), .O(n2814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2265_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n28408), 
            .O(n5939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2265_3 (.CI(n28408), .I0(n2083), .I1(n99), .CO(n28409));
    SB_CARRY rem_4_add_1854_14 (.CI(n28878), .I0(n2747), .I1(VCC_net), 
            .CO(n28879));
    SB_LUT4 rem_4_add_1854_13_lut (.I0(GND_net), .I1(n2748), .I2(VCC_net), 
            .I3(n28877), .O(n2815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2265_2_lut (.I0(GND_net), .I1(n662), .I2(n558), .I3(VCC_net), 
            .O(n5940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2265_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_13 (.CI(n28877), .I0(n2748), .I1(VCC_net), 
            .CO(n28878));
    SB_CARRY add_2265_2 (.CI(VCC_net), .I0(n662), .I1(n558), .CO(n28408));
    SB_LUT4 add_2264_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n28407), 
            .O(n5908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_12_lut (.I0(GND_net), .I1(n2749), .I2(VCC_net), 
            .I3(n28876), .O(n2816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_12 (.CI(n28876), .I0(n2749), .I1(VCC_net), 
            .CO(n28877));
    SB_LUT4 add_2264_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n28406), 
            .O(n5909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_15 (.CI(n28406), .I0(n1968), .I1(n87), .CO(n28407));
    SB_LUT4 rem_4_add_1854_11_lut (.I0(GND_net), .I1(n2750), .I2(VCC_net), 
            .I3(n28875), .O(n2817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_11 (.CI(n28875), .I0(n2750), .I1(VCC_net), 
            .CO(n28876));
    SB_LUT4 rem_4_add_1854_10_lut (.I0(GND_net), .I1(n2751), .I2(VCC_net), 
            .I3(n28874), .O(n2818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2264_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n28405), 
            .O(n5910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_14 (.CI(n28405), .I0(n1969), .I1(n88), .CO(n28406));
    SB_LUT4 add_2264_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n28404), 
            .O(n5911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_10 (.CI(n28874), .I0(n2751), .I1(VCC_net), 
            .CO(n28875));
    SB_LUT4 rem_4_add_1854_9_lut (.I0(GND_net), .I1(n2752), .I2(VCC_net), 
            .I3(n28873), .O(n2819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_7 (.CI(n27978), .I0(n1153), .I1(VCC_net), .CO(n27979));
    SB_DFF communication_counter_1176__i3 (.Q(communication_counter[3]), .C(LED_c), 
           .D(n162));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i4 (.Q(communication_counter[4]), .C(LED_c), 
           .D(n161));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i5 (.Q(communication_counter[5]), .C(LED_c), 
           .D(n160));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i6 (.Q(communication_counter[6]), .C(LED_c), 
           .D(n159));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i7 (.Q(communication_counter[7]), .C(LED_c), 
           .D(n158));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i8 (.Q(communication_counter[8]), .C(LED_c), 
           .D(n157));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i9 (.Q(communication_counter[9]), .C(LED_c), 
           .D(n156));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i10 (.Q(communication_counter[10]), 
           .C(LED_c), .D(n155));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i11 (.Q(communication_counter[11]), 
           .C(LED_c), .D(n154));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i12 (.Q(communication_counter[12]), 
           .C(LED_c), .D(n153));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i13 (.Q(communication_counter[13]), 
           .C(LED_c), .D(n152));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i14 (.Q(communication_counter[14]), 
           .C(LED_c), .D(n151));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i15 (.Q(communication_counter[15]), 
           .C(LED_c), .D(n150));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i16 (.Q(communication_counter[16]), 
           .C(LED_c), .D(n149));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i17 (.Q(communication_counter[17]), 
           .C(LED_c), .D(n148));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i18 (.Q(communication_counter[18]), 
           .C(LED_c), .D(n147));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i19 (.Q(communication_counter[19]), 
           .C(LED_c), .D(n146));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i20 (.Q(communication_counter[20]), 
           .C(LED_c), .D(n145));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i21 (.Q(communication_counter[21]), 
           .C(LED_c), .D(n144));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i22 (.Q(communication_counter[22]), 
           .C(LED_c), .D(n143));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i23 (.Q(communication_counter[23]), 
           .C(LED_c), .D(n142));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i24 (.Q(communication_counter[24]), 
           .C(LED_c), .D(n141));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i25 (.Q(communication_counter[25]), 
           .C(LED_c), .D(n140));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i26 (.Q(communication_counter[26]), 
           .C(LED_c), .D(n139));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i27 (.Q(communication_counter[27]), 
           .C(LED_c), .D(n138));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i28 (.Q(communication_counter[28]), 
           .C(LED_c), .D(n137));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i29 (.Q(communication_counter[29]), 
           .C(LED_c), .D(n136));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i30 (.Q(communication_counter[30]), 
           .C(LED_c), .D(n135));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_DFF communication_counter_1176__i31 (.Q(communication_counter[31]), 
           .C(LED_c), .D(n134));   // verilog/TinyFPGA_B.v(74[28:51])
    SB_LUT4 div_46_i1759_3_lut_3_lut (.I0(n2642), .I1(n6053), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2264_13 (.CI(n28404), .I0(n1970), .I1(n89), .CO(n28405));
    SB_CARRY rem_4_add_1854_9 (.CI(n28873), .I0(n2752), .I1(VCC_net), 
            .CO(n28874));
    SB_LUT4 rem_4_add_1854_8_lut (.I0(GND_net), .I1(n2753), .I2(VCC_net), 
            .I3(n28872), .O(n2820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_8 (.CI(n28872), .I0(n2753), .I1(VCC_net), 
            .CO(n28873));
    SB_LUT4 rem_4_add_1854_7_lut (.I0(GND_net), .I1(n2754), .I2(GND_net), 
            .I3(n28871), .O(n2821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2264_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n28403), 
            .O(n5912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_7 (.CI(n28871), .I0(n2754), .I1(GND_net), 
            .CO(n28872));
    SB_LUT4 rem_4_add_1854_6_lut (.I0(GND_net), .I1(n2755), .I2(GND_net), 
            .I3(n28870), .O(n2822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_12 (.CI(n28403), .I0(n1971), .I1(n90), .CO(n28404));
    SB_CARRY rem_4_add_1854_6 (.CI(n28870), .I0(n2755), .I1(GND_net), 
            .CO(n28871));
    SB_LUT4 add_2264_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n28402), 
            .O(n5913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_6_lut (.I0(GND_net), .I1(n1154), .I2(GND_net), 
            .I3(n27977), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_6 (.CI(n27977), .I0(n1154), .I1(GND_net), .CO(n27978));
    SB_CARRY add_2264_11 (.CI(n28402), .I0(n1972), .I1(n91), .CO(n28403));
    SB_LUT4 add_2264_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n28401), 
            .O(n5914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_10 (.CI(n28401), .I0(n1973), .I1(n92), .CO(n28402));
    SB_LUT4 rem_4_add_1854_5_lut (.I0(GND_net), .I1(n2756), .I2(VCC_net), 
            .I3(n28869), .O(n2823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_5 (.CI(n28869), .I0(n2756), .I1(VCC_net), 
            .CO(n28870));
    SB_LUT4 rem_4_add_1854_4_lut (.I0(GND_net), .I1(n2757), .I2(VCC_net), 
            .I3(n28868), .O(n2824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2264_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n28400), 
            .O(n5915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_4 (.CI(n28868), .I0(n2757), .I1(VCC_net), 
            .CO(n28869));
    SB_LUT4 rem_4_add_1854_3_lut (.I0(GND_net), .I1(n2758), .I2(GND_net), 
            .I3(n28867), .O(n2825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_9 (.CI(n28400), .I0(n1974), .I1(n93), .CO(n28401));
    SB_LUT4 add_2264_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n28399), 
            .O(n5916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1760_3_lut_3_lut (.I0(n2642), .I1(n6054), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2264_8 (.CI(n28399), .I0(n1975), .I1(n94), .CO(n28400));
    SB_LUT4 add_2264_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n28398), 
            .O(n5917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i889_3_lut_3_lut (.I0(n1316), .I1(n5833), .I2(n1298), 
            .I3(GND_net), .O(n1418));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i889_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1764_3_lut_3_lut (.I0(n2642), .I1(n6058), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2264_7 (.CI(n28398), .I0(n1976), .I1(n95), .CO(n28399));
    SB_LUT4 add_2264_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n28397), 
            .O(n5918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1765_3_lut_3_lut (.I0(n2642), .I1(n6059), .I2(n2629), 
            .I3(GND_net), .O(n2710_adj_4419));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2264_6 (.CI(n28397), .I0(n1977), .I1(n96), .CO(n28398));
    SB_LUT4 add_2264_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n28396), 
            .O(n5919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_5 (.CI(n28396), .I0(n1978), .I1(n97), .CO(n28397));
    SB_LUT4 add_2264_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n28395), 
            .O(n5920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_4 (.CI(n28395), .I0(n1979), .I1(n98), .CO(n28396));
    SB_LUT4 add_2264_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n28394), 
            .O(n5921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_3 (.CI(n28394), .I0(n1980), .I1(n99), .CO(n28395));
    SB_CARRY rem_4_add_1854_3 (.CI(n28867), .I0(n2758), .I1(GND_net), 
            .CO(n28868));
    SB_CARRY rem_4_add_1854_2 (.CI(VCC_net), .I0(n2858), .I1(VCC_net), 
            .CO(n28867));
    SB_LUT4 div_46_i1766_3_lut_3_lut (.I0(n2642), .I1(n6060), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4596), .I3(n28866), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2264_2_lut (.I0(GND_net), .I1(n661), .I2(n558), .I3(VCC_net), 
            .O(n5922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2264_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_5_lut (.I0(GND_net), .I1(n1155), .I2(GND_net), 
            .I3(n27976), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2264_2 (.CI(VCC_net), .I0(n661), .I1(n558), .CO(n28394));
    SB_LUT4 add_2263_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n28393), 
            .O(n5892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4597), .I3(n28865), .O(n3_adj_4382)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2263_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n28392), 
            .O(n5893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_24 (.CI(n28865), .I0(GND_net), .I1(n3_adj_4597), 
            .CO(n28866));
    SB_LUT4 div_46_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4598), .I3(n28864), .O(n4_adj_4356)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_14 (.CI(n28392), .I0(n1863), .I1(n88), .CO(n28393));
    SB_CARRY div_46_unary_minus_2_add_3_23 (.CI(n28864), .I0(GND_net), .I1(n4_adj_4598), 
            .CO(n28865));
    SB_LUT4 add_2263_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n28391), 
            .O(n5894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_13 (.CI(n28391), .I0(n1864), .I1(n89), .CO(n28392));
    SB_LUT4 add_2263_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n28390), 
            .O(n5895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4599), .I3(n28863), .O(n5_adj_4343)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_22 (.CI(n28863), .I0(GND_net), .I1(n5_adj_4599), 
            .CO(n28864));
    SB_LUT4 div_46_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4600), .I3(n28862), .O(n6_adj_4367)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_21 (.CI(n28862), .I0(GND_net), .I1(n6_adj_4600), 
            .CO(n28863));
    SB_LUT4 div_46_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4601), .I3(n28861), .O(n7_adj_4376)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_20 (.CI(n28861), .I0(GND_net), .I1(n7_adj_4601), 
            .CO(n28862));
    SB_LUT4 div_46_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4602), .I3(n28860), .O(n8_adj_4381)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_19 (.CI(n28860), .I0(GND_net), .I1(n8_adj_4602), 
            .CO(n28861));
    SB_LUT4 div_46_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4603), .I3(n28859), .O(n9_adj_4359)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_12 (.CI(n28390), .I0(n1865), .I1(n90), .CO(n28391));
    SB_CARRY div_46_unary_minus_2_add_3_18 (.CI(n28859), .I0(GND_net), .I1(n9_adj_4603), 
            .CO(n28860));
    SB_LUT4 rem_4_add_983_13_lut (.I0(n1481), .I1(n1448), .I2(VCC_net), 
            .I3(n29111), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2263_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n28389), 
            .O(n5896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_12_lut (.I0(GND_net), .I1(n1449), .I2(VCC_net), 
            .I3(n29110), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_12 (.CI(n29110), .I0(n1449), .I1(VCC_net), 
            .CO(n29111));
    SB_LUT4 div_46_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4604), .I3(n28858), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_11_lut (.I0(GND_net), .I1(n1450), .I2(VCC_net), 
            .I3(n29109), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_17 (.CI(n28858), .I0(GND_net), .I1(n10_adj_4604), 
            .CO(n28859));
    SB_LUT4 div_46_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4605), .I3(n28857), .O(n11_adj_4344)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_16 (.CI(n28857), .I0(GND_net), .I1(n11_adj_4605), 
            .CO(n28858));
    SB_LUT4 div_46_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4606), .I3(n28856), .O(n12_adj_4345)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_11 (.CI(n28389), .I0(n1866), .I1(n91), .CO(n28390));
    SB_CARRY rem_4_add_983_11 (.CI(n29109), .I0(n1450), .I1(VCC_net), 
            .CO(n29110));
    SB_CARRY div_46_unary_minus_2_add_3_15 (.CI(n28856), .I0(GND_net), .I1(n12_adj_4606), 
            .CO(n28857));
    SB_LUT4 add_2263_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n28388), 
            .O(n5897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_10 (.CI(n28388), .I0(n1867), .I1(n92), .CO(n28389));
    SB_LUT4 add_2263_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n28387), 
            .O(n5898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4607), .I3(n28855), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_14 (.CI(n28855), .I0(GND_net), .I1(n13_adj_4607), 
            .CO(n28856));
    SB_LUT4 rem_4_add_983_10_lut (.I0(GND_net), .I1(n1451), .I2(VCC_net), 
            .I3(n29108), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_10 (.CI(n29108), .I0(n1451), .I1(VCC_net), 
            .CO(n29109));
    SB_LUT4 rem_4_add_983_9_lut (.I0(GND_net), .I1(n1452), .I2(VCC_net), 
            .I3(n29107), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4608), .I3(n28854), .O(n14_adj_4377)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_13 (.CI(n28854), .I0(GND_net), .I1(n14_adj_4608), 
            .CO(n28855));
    SB_CARRY rem_4_add_983_9 (.CI(n29107), .I0(n1452), .I1(VCC_net), .CO(n29108));
    SB_LUT4 rem_4_add_983_8_lut (.I0(GND_net), .I1(n1453), .I2(VCC_net), 
            .I3(n29106), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4609), .I3(n28853), .O(n15_adj_4320)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_8 (.CI(n29106), .I0(n1453), .I1(VCC_net), .CO(n29107));
    SB_CARRY div_46_unary_minus_2_add_3_12 (.CI(n28853), .I0(GND_net), .I1(n15_adj_4609), 
            .CO(n28854));
    SB_LUT4 rem_4_add_983_7_lut (.I0(GND_net), .I1(n1454), .I2(GND_net), 
            .I3(n29105), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4610), .I3(n28852), .O(n16_adj_4378)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_11 (.CI(n28852), .I0(GND_net), .I1(n16_adj_4610), 
            .CO(n28853));
    SB_LUT4 i12596_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n13195), .I3(GND_net), .O(n17278));   // verilog/coms.v(126[12] 289[6])
    defparam i12596_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_983_7 (.CI(n29105), .I0(n1454), .I1(GND_net), .CO(n29106));
    SB_LUT4 div_46_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4611), .I3(n28851), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1718 (.I0(bit_ctr[19]), .I1(n40174), .I2(n4385), 
            .I3(GND_net), .O(n33329));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1718.LUT_INIT = 16'hacac;
    SB_CARRY add_2263_9 (.CI(n28387), .I0(n1868), .I1(n93), .CO(n28388));
    SB_LUT4 div_46_i1767_3_lut_3_lut (.I0(n2642), .I1(n6061), .I2(n2631), 
            .I3(GND_net), .O(n2712_adj_4420));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2263_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n28386), 
            .O(n5899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_6_lut (.I0(GND_net), .I1(n1455), .I2(GND_net), 
            .I3(n29104), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_6 (.CI(n29104), .I0(n1455), .I1(GND_net), .CO(n29105));
    SB_CARRY div_46_unary_minus_2_add_3_10 (.CI(n28851), .I0(GND_net), .I1(n17_adj_4611), 
            .CO(n28852));
    SB_LUT4 div_46_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4612), .I3(n28850), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12857_3_lut (.I0(encoder1_position[14]), .I1(n2900), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17539));   // quad.v(35[10] 41[6])
    defparam i12857_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2263_8 (.CI(n28386), .I0(n1869), .I1(n94), .CO(n28387));
    SB_LUT4 rem_4_add_983_5_lut (.I0(GND_net), .I1(n1456), .I2(VCC_net), 
            .I3(n29103), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_5 (.CI(n29103), .I0(n1456), .I1(VCC_net), .CO(n29104));
    SB_CARRY rem_4_add_782_5 (.CI(n27976), .I0(n1155), .I1(GND_net), .CO(n27977));
    SB_CARRY div_46_unary_minus_2_add_3_9 (.CI(n28850), .I0(GND_net), .I1(n18_adj_4612), 
            .CO(n28851));
    SB_LUT4 add_2263_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n28385), 
            .O(n5900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4613), .I3(n28849), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_8 (.CI(n28849), .I0(GND_net), .I1(n19_adj_4613), 
            .CO(n28850));
    SB_CARRY add_2263_7 (.CI(n28385), .I0(n1870), .I1(n95), .CO(n28386));
    SB_LUT4 rem_4_add_983_4_lut (.I0(GND_net), .I1(n1457), .I2(VCC_net), 
            .I3(n29102), .O(n1524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_4_lut (.I0(GND_net), .I1(n1156), .I2(VCC_net), 
            .I3(n27975), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1775_3_lut_3_lut (.I0(n2642), .I1(n6069), .I2(n668), 
            .I3(GND_net), .O(n2720_adj_4424));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4614), .I3(n28848), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_4 (.CI(n29102), .I0(n1457), .I1(VCC_net), .CO(n29103));
    SB_LUT4 add_2263_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n28384), 
            .O(n5901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_7 (.CI(n28848), .I0(GND_net), .I1(n20_adj_4614), 
            .CO(n28849));
    SB_LUT4 rem_4_add_983_3_lut (.I0(GND_net), .I1(n1458), .I2(GND_net), 
            .I3(n29101), .O(n1525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4615), .I3(n28847), .O(n21_adj_4392)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_6 (.CI(n28847), .I0(GND_net), .I1(n21_adj_4615), 
            .CO(n28848));
    SB_CARRY rem_4_add_983_3 (.CI(n29101), .I0(n1458), .I1(GND_net), .CO(n29102));
    SB_CARRY rem_4_add_983_2 (.CI(VCC_net), .I0(n1558), .I1(VCC_net), 
            .CO(n29101));
    SB_LUT4 div_46_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4616), .I3(n28846), .O(n22_adj_4357)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_14_lut (.I0(n1580), .I1(n1547), .I2(VCC_net), 
            .I3(n29100), .O(n1646_adj_4525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2263_6 (.CI(n28384), .I0(n1871), .I1(n96), .CO(n28385));
    SB_CARRY div_46_unary_minus_2_add_3_5 (.CI(n28846), .I0(GND_net), .I1(n22_adj_4616), 
            .CO(n28847));
    SB_LUT4 rem_4_add_1050_13_lut (.I0(GND_net), .I1(n1548), .I2(VCC_net), 
            .I3(n29099), .O(n1615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4617), .I3(n28845), .O(n23_adj_4393)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_13 (.CI(n29099), .I0(n1548), .I1(VCC_net), 
            .CO(n29100));
    SB_LUT4 add_2263_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n28383), 
            .O(n5902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_4 (.CI(n28845), .I0(GND_net), .I1(n23_adj_4617), 
            .CO(n28846));
    SB_LUT4 rem_4_add_1050_12_lut (.I0(GND_net), .I1(n1549), .I2(VCC_net), 
            .I3(n29098), .O(n1616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_5 (.CI(n28383), .I0(n1872), .I1(n97), .CO(n28384));
    SB_LUT4 div_46_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4618), .I3(n28844), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_12 (.CI(n29098), .I0(n1549), .I1(VCC_net), 
            .CO(n29099));
    SB_CARRY div_46_unary_minus_2_add_3_3 (.CI(n28844), .I0(GND_net), .I1(n24_adj_4618), 
            .CO(n28845));
    SB_LUT4 add_2263_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n28382), 
            .O(n5903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4619), .I3(VCC_net), .O(n25_adj_4358)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_4 (.CI(n28382), .I0(n1873), .I1(n98), .CO(n28383));
    SB_LUT4 add_2263_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n28381), 
            .O(n5904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_3 (.CI(n28381), .I0(n1874), .I1(n99), .CO(n28382));
    SB_LUT4 add_2263_2_lut (.I0(GND_net), .I1(n660), .I2(n558), .I3(VCC_net), 
            .O(n5905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2263_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2263_2 (.CI(VCC_net), .I0(n660), .I1(n558), .CO(n28381));
    SB_LUT4 div_46_i1768_3_lut_3_lut (.I0(n2642), .I1(n6062), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1772_3_lut_3_lut (.I0(n2642), .I1(n6066), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_46_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4619), 
            .CO(n28844));
    SB_LUT4 add_2262_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n28380), 
            .O(n5877)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2262_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n28379), 
            .O(n5878)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2262_13 (.CI(n28379), .I0(n1755), .I1(n89), .CO(n28380));
    SB_LUT4 add_2262_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n28378), 
            .O(n5879)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12597_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n13195), .I3(GND_net), .O(n17279));   // verilog/coms.v(126[12] 289[6])
    defparam i12597_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_782_4 (.CI(n27975), .I0(n1156), .I1(VCC_net), .CO(n27976));
    SB_CARRY add_2262_12 (.CI(n28378), .I0(n1756), .I1(n90), .CO(n28379));
    SB_LUT4 add_2262_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n28377), 
            .O(n5880)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2262_11 (.CI(n28377), .I0(n1757), .I1(n91), .CO(n28378));
    SB_LUT4 add_2262_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n28376), 
            .O(n5881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2262_10 (.CI(n28376), .I0(n1758), .I1(n92), .CO(n28377));
    SB_LUT4 i12598_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n13195), .I3(GND_net), .O(n17280));   // verilog/coms.v(126[12] 289[6])
    defparam i12598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2262_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n28375), 
            .O(n5882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2262_9 (.CI(n28375), .I0(n1759), .I1(n93), .CO(n28376));
    SB_LUT4 i12856_3_lut (.I0(encoder1_position[13]), .I1(n2901), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17538));   // quad.v(35[10] 41[6])
    defparam i12856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2262_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n28374), 
            .O(n5883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2262_8 (.CI(n28374), .I0(n1760), .I1(n94), .CO(n28375));
    SB_LUT4 i12599_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n13195), .I3(GND_net), .O(n17281));   // verilog/coms.v(126[12] 289[6])
    defparam i12599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1763_3_lut_3_lut (.I0(n2642), .I1(n6057), .I2(n2627), 
            .I3(GND_net), .O(n2708_adj_4418));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12855_3_lut (.I0(encoder1_position[12]), .I1(n2902), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17537));   // quad.v(35[10] 41[6])
    defparam i12855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2262_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n28373), 
            .O(n5884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12854_3_lut (.I0(encoder1_position[11]), .I1(n2903), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17536));   // quad.v(35[10] 41[6])
    defparam i12854_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2262_7 (.CI(n28373), .I0(n1761), .I1(n95), .CO(n28374));
    SB_LUT4 i12853_3_lut (.I0(encoder1_position[10]), .I1(n2904), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17535));   // quad.v(35[10] 41[6])
    defparam i12853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2262_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n28372), 
            .O(n5885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_11_lut (.I0(GND_net), .I1(n1550), .I2(VCC_net), 
            .I3(n29097), .O(n1617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4572), .I3(n28843), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2262_6 (.CI(n28372), .I0(n1762), .I1(n96), .CO(n28373));
    SB_LUT4 i12852_3_lut (.I0(encoder1_position[9]), .I1(n2905), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17534));   // quad.v(35[10] 41[6])
    defparam i12852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2262_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n28371), 
            .O(n5886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2262_5 (.CI(n28371), .I0(n1763), .I1(n97), .CO(n28372));
    SB_LUT4 add_2262_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n28370), 
            .O(n5887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_11 (.CI(n29097), .I0(n1550), .I1(VCC_net), 
            .CO(n29098));
    SB_CARRY add_2262_4 (.CI(n28370), .I0(n1764), .I1(n98), .CO(n28371));
    SB_LUT4 rem_4_add_1050_10_lut (.I0(GND_net), .I1(n1551), .I2(VCC_net), 
            .I3(n29096), .O(n1618)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4573), .I3(n28842), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_10 (.CI(n29096), .I0(n1551), .I1(VCC_net), 
            .CO(n29097));
    SB_LUT4 add_2262_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n28369), 
            .O(n5888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_24 (.CI(n28842), .I0(GND_net), .I1(n3_adj_4573), 
            .CO(n28843));
    SB_CARRY add_2262_3 (.CI(n28369), .I0(n1765), .I1(n99), .CO(n28370));
    SB_LUT4 add_2262_2_lut (.I0(GND_net), .I1(n659), .I2(n558), .I3(VCC_net), 
            .O(n5889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2262_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2262_2 (.CI(VCC_net), .I0(n659), .I1(n558), .CO(n28369));
    SB_LUT4 add_2261_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n28368), 
            .O(n5863)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1770_3_lut_3_lut (.I0(n2642), .I1(n6064), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4574), .I3(n28841), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2261_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n28367), 
            .O(n5864)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_12 (.CI(n28367), .I0(n1644), .I1(n90), .CO(n28368));
    SB_LUT4 add_2261_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n28366), 
            .O(n5865)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_9_lut (.I0(GND_net), .I1(n1552), .I2(VCC_net), 
            .I3(n29095), .O(n1619)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_23 (.CI(n28841), .I0(GND_net), .I1(n4_adj_4574), 
            .CO(n28842));
    SB_CARRY add_2261_11 (.CI(n28366), .I0(n1645), .I1(n91), .CO(n28367));
    SB_LUT4 div_46_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4575), .I3(n28840), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_9 (.CI(n29095), .I0(n1552), .I1(VCC_net), 
            .CO(n29096));
    SB_LUT4 add_2261_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n28365), 
            .O(n5866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_8_lut (.I0(GND_net), .I1(n1553_adj_4533), .I2(VCC_net), 
            .I3(n29094), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_10 (.CI(n28365), .I0(n1646), .I1(n92), .CO(n28366));
    SB_CARRY div_46_unary_minus_4_add_3_22 (.CI(n28840), .I0(GND_net), .I1(n5_adj_4575), 
            .CO(n28841));
    SB_LUT4 div_46_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4576), .I3(n28839), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2261_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n28364), 
            .O(n5867)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1719 (.I0(bit_ctr[11]), .I1(n40176), .I2(n4385), 
            .I3(GND_net), .O(n33333));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1719.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1050_8 (.CI(n29094), .I0(n1553_adj_4533), .I1(VCC_net), 
            .CO(n29095));
    SB_CARRY add_2261_9 (.CI(n28364), .I0(n1647), .I1(n93), .CO(n28365));
    SB_LUT4 add_2261_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n28363), 
            .O(n5868)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_8 (.CI(n28363), .I0(n1648), .I1(n94), .CO(n28364));
    SB_LUT4 add_2261_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n28362), 
            .O(n5869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_7 (.CI(n28362), .I0(n1649), .I1(n95), .CO(n28363));
    SB_CARRY div_46_unary_minus_4_add_3_21 (.CI(n28839), .I0(GND_net), .I1(n6_adj_4576), 
            .CO(n28840));
    SB_LUT4 rem_4_i1053_3_lut (.I0(n1548), .I1(n1615), .I2(n1580), .I3(GND_net), 
            .O(n1647_adj_4526));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1050_7_lut (.I0(GND_net), .I1(n1554_adj_4534), .I2(GND_net), 
            .I3(n29093), .O(n1621)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2261_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n28361), 
            .O(n5870)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_6 (.CI(n28361), .I0(n1650), .I1(n96), .CO(n28362));
    SB_LUT4 add_2261_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n28360), 
            .O(n5871)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4577), .I3(n28838), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_7 (.CI(n29093), .I0(n1554_adj_4534), .I1(GND_net), 
            .CO(n29094));
    SB_CARRY div_46_unary_minus_4_add_3_20 (.CI(n28838), .I0(GND_net), .I1(n7_adj_4577), 
            .CO(n28839));
    SB_CARRY add_2261_5 (.CI(n28360), .I0(n1651), .I1(n97), .CO(n28361));
    SB_LUT4 add_2261_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n28359), 
            .O(n5872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1774_3_lut_3_lut (.I0(n2642), .I1(n6068), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1050_6_lut (.I0(GND_net), .I1(n1555), .I2(GND_net), 
            .I3(n29092), .O(n1622)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_6 (.CI(n29092), .I0(n1555), .I1(GND_net), 
            .CO(n29093));
    SB_LUT4 div_46_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4578), .I3(n28837), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_4 (.CI(n28359), .I0(n1652), .I1(n98), .CO(n28360));
    SB_LUT4 add_2261_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n28358), 
            .O(n5873)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_3 (.CI(n28358), .I0(n1653), .I1(n99), .CO(n28359));
    SB_LUT4 div_46_i1773_3_lut_3_lut (.I0(n2642), .I1(n6067), .I2(n2637), 
            .I3(GND_net), .O(n2718_adj_4423));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2261_2_lut (.I0(GND_net), .I1(n658), .I2(n558), .I3(VCC_net), 
            .O(n5874)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2261_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2261_2 (.CI(VCC_net), .I0(n658), .I1(n558), .CO(n28358));
    SB_LUT4 rem_4_add_1050_5_lut (.I0(GND_net), .I1(n1556), .I2(VCC_net), 
            .I3(n29091), .O(n1623)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_19 (.CI(n28837), .I0(GND_net), .I1(n8_adj_4578), 
            .CO(n28838));
    SB_LUT4 add_2260_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n28357), 
            .O(n5850)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4579), .I3(n28836), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2260_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n28356), 
            .O(n5851)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2260_11 (.CI(n28356), .I0(n1530), .I1(n91), .CO(n28357));
    SB_LUT4 add_2260_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n28355), 
            .O(n5852)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2260_10 (.CI(n28355), .I0(n1531), .I1(n92), .CO(n28356));
    SB_LUT4 add_2260_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n28354), 
            .O(n5853)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2260_9 (.CI(n28354), .I0(n1532), .I1(n93), .CO(n28355));
    SB_LUT4 add_2260_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n28353), 
            .O(n5854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_18 (.CI(n28836), .I0(GND_net), .I1(n9_adj_4579), 
            .CO(n28837));
    SB_CARRY add_2260_8 (.CI(n28353), .I0(n1533), .I1(n94), .CO(n28354));
    SB_LUT4 div_46_i1771_3_lut_3_lut (.I0(n2642), .I1(n6065), .I2(n2635), 
            .I3(GND_net), .O(n2716_adj_4422));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1050_5 (.CI(n29091), .I0(n1556), .I1(VCC_net), 
            .CO(n29092));
    SB_LUT4 div_46_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4580), .I3(n28835), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2260_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n28352), 
            .O(n5855)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_4_lut (.I0(GND_net), .I1(n1557), .I2(VCC_net), 
            .I3(n29090), .O(n1624)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_17 (.CI(n28835), .I0(GND_net), .I1(n10_adj_4580), 
            .CO(n28836));
    SB_CARRY add_2260_7 (.CI(n28352), .I0(n1534), .I1(n95), .CO(n28353));
    SB_LUT4 add_2260_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n28351), 
            .O(n5856)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2260_6 (.CI(n28351), .I0(n1535), .I1(n96), .CO(n28352));
    SB_CARRY rem_4_add_1050_4 (.CI(n29090), .I0(n1557), .I1(VCC_net), 
            .CO(n29091));
    SB_LUT4 div_46_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4581), .I3(n28834), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2260_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n28350), 
            .O(n5857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2260_5 (.CI(n28350), .I0(n1536), .I1(n97), .CO(n28351));
    SB_LUT4 add_2260_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n28349), 
            .O(n5858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2260_4 (.CI(n28349), .I0(n1537), .I1(n98), .CO(n28350));
    SB_LUT4 rem_4_add_1050_3_lut (.I0(GND_net), .I1(n1558), .I2(GND_net), 
            .I3(n29089), .O(n1625)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2260_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n28348), 
            .O(n5859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_16 (.CI(n28834), .I0(GND_net), .I1(n11_adj_4581), 
            .CO(n28835));
    SB_CARRY rem_4_add_1050_3 (.CI(n29089), .I0(n1558), .I1(GND_net), 
            .CO(n29090));
    SB_CARRY add_2260_3 (.CI(n28348), .I0(n1538), .I1(n99), .CO(n28349));
    SB_LUT4 div_46_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4582), .I3(n28833), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_15 (.CI(n28833), .I0(GND_net), .I1(n12_adj_4582), 
            .CO(n28834));
    SB_LUT4 add_2260_2_lut (.I0(GND_net), .I1(n657), .I2(n558), .I3(VCC_net), 
            .O(n5860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2260_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2260_2 (.CI(VCC_net), .I0(n657), .I1(n558), .CO(n28348));
    SB_LUT4 add_2259_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n28347), 
            .O(n5838)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_2 (.CI(VCC_net), .I0(n1658), .I1(VCC_net), 
            .CO(n29089));
    SB_LUT4 rem_4_add_1117_15_lut (.I0(n1679), .I1(n1646_adj_4525), .I2(VCC_net), 
            .I3(n29088), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4583), .I3(n28832), .O(n63_adj_4324)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2259_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n28346), 
            .O(n5839)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2259_10 (.CI(n28346), .I0(n1413), .I1(n92), .CO(n28347));
    SB_LUT4 add_2259_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n28345), 
            .O(n5840)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_14_lut (.I0(GND_net), .I1(n1647_adj_4526), .I2(VCC_net), 
            .I3(n29087), .O(n1714)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_14 (.CI(n28832), .I0(GND_net), .I1(n13_adj_4583), 
            .CO(n28833));
    SB_CARRY add_2259_9 (.CI(n28345), .I0(n1414), .I1(n93), .CO(n28346));
    SB_LUT4 add_2259_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n28344), 
            .O(n5841)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2259_8 (.CI(n28344), .I0(n1415), .I1(n94), .CO(n28345));
    SB_LUT4 div_46_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4584), .I3(n28831), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2259_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n28343), 
            .O(n5842)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2259_7 (.CI(n28343), .I0(n1416), .I1(n95), .CO(n28344));
    SB_LUT4 add_2259_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n28342), 
            .O(n5843)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2259_6 (.CI(n28342), .I0(n1417), .I1(n96), .CO(n28343));
    SB_LUT4 add_2259_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n28341), 
            .O(n5844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2259_5 (.CI(n28341), .I0(n1418), .I1(n97), .CO(n28342));
    SB_LUT4 add_2259_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n28340), 
            .O(n5845)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_14 (.CI(n29087), .I0(n1647_adj_4526), .I1(VCC_net), 
            .CO(n29088));
    SB_CARRY div_46_unary_minus_4_add_3_13 (.CI(n28831), .I0(GND_net), .I1(n14_adj_4584), 
            .CO(n28832));
    SB_CARRY add_2259_4 (.CI(n28340), .I0(n1419), .I1(n98), .CO(n28341));
    SB_LUT4 add_2259_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n28339), 
            .O(n5846)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_13_lut (.I0(GND_net), .I1(n1648_adj_4527), .I2(VCC_net), 
            .I3(n29086), .O(n1715)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4585), .I3(n28830), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2259_3 (.CI(n28339), .I0(n1420), .I1(n99), .CO(n28340));
    SB_CARRY rem_4_add_1117_13 (.CI(n29086), .I0(n1648_adj_4527), .I1(VCC_net), 
            .CO(n29087));
    SB_CARRY div_46_unary_minus_4_add_3_12 (.CI(n28830), .I0(GND_net), .I1(n15_adj_4585), 
            .CO(n28831));
    SB_LUT4 add_2259_2_lut (.I0(GND_net), .I1(n656), .I2(n558), .I3(VCC_net), 
            .O(n5847)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2259_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2259_2 (.CI(VCC_net), .I0(n656), .I1(n558), .CO(n28339));
    SB_LUT4 add_2258_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n28338), 
            .O(n5827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2258_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n28337), 
            .O(n5828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12600_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n13195), .I3(GND_net), .O(n17282));   // verilog/coms.v(126[12] 289[6])
    defparam i12600_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2258_9 (.CI(n28337), .I0(n1293), .I1(n93), .CO(n28338));
    SB_LUT4 rem_4_add_1117_12_lut (.I0(GND_net), .I1(n1649_adj_4528), .I2(VCC_net), 
            .I3(n29085), .O(n1716)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4586), .I3(n28829), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2258_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n28336), 
            .O(n5829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2258_8 (.CI(n28336), .I0(n1294), .I1(n94), .CO(n28337));
    SB_CARRY div_46_unary_minus_4_add_3_11 (.CI(n28829), .I0(GND_net), .I1(n16_adj_4586), 
            .CO(n28830));
    SB_LUT4 add_2258_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n28335), 
            .O(n5830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2258_7 (.CI(n28335), .I0(n1295), .I1(n95), .CO(n28336));
    SB_LUT4 add_2258_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n28334), 
            .O(n5831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2258_6 (.CI(n28334), .I0(n1296), .I1(n96), .CO(n28335));
    SB_LUT4 add_2258_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n28333), 
            .O(n5832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2258_5 (.CI(n28333), .I0(n1297), .I1(n97), .CO(n28334));
    SB_LUT4 add_2258_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n28332), 
            .O(n5833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_3_lut_adj_1720 (.I0(bit_ctr[10]), .I1(n40175), .I2(n4385), 
            .I3(GND_net), .O(n33331));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1720.LUT_INIT = 16'hacac;
    SB_CARRY add_2258_4 (.CI(n28332), .I0(n1298), .I1(n98), .CO(n28333));
    SB_CARRY rem_4_add_1117_12 (.CI(n29085), .I0(n1649_adj_4528), .I1(VCC_net), 
            .CO(n29086));
    SB_LUT4 div_46_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4587), .I3(n28828), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_11_lut (.I0(GND_net), .I1(n1650_adj_4529), .I2(VCC_net), 
            .I3(n29084), .O(n1717)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_10 (.CI(n28828), .I0(GND_net), .I1(n17_adj_4587), 
            .CO(n28829));
    SB_LUT4 i12347_3_lut (.I0(n16772), .I1(r_Bit_Index_adj_5055[0]), .I2(n16641), 
            .I3(GND_net), .O(n17029));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12347_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i12866_3_lut (.I0(encoder1_position[23]), .I1(n2891), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17548));   // quad.v(35[10] 41[6])
    defparam i12866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2258_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n28331), 
            .O(n5834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12865_3_lut (.I0(encoder1_position[22]), .I1(n2892), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17547));   // quad.v(35[10] 41[6])
    defparam i12865_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1117_11 (.CI(n29084), .I0(n1650_adj_4529), .I1(VCC_net), 
            .CO(n29085));
    SB_LUT4 rem_4_add_1117_10_lut (.I0(GND_net), .I1(n1651_adj_4530), .I2(VCC_net), 
            .I3(n29083), .O(n1718)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_10 (.CI(n29083), .I0(n1651_adj_4530), .I1(VCC_net), 
            .CO(n29084));
    SB_LUT4 div_46_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4588), .I3(n28827), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2258_3 (.CI(n28331), .I0(n1299), .I1(n99), .CO(n28332));
    SB_LUT4 add_2258_2_lut (.I0(GND_net), .I1(n655), .I2(n558), .I3(VCC_net), 
            .O(n5835)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2258_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2258_2 (.CI(VCC_net), .I0(n655), .I1(n558), .CO(n28331));
    SB_LUT4 add_2257_9_lut (.I0(GND_net), .I1(n1169_adj_4409), .I2(n93), 
            .I3(n28330), .O(n5817)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2257_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n28329), 
            .O(n5818)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_9 (.CI(n28827), .I0(GND_net), .I1(n18_adj_4588), 
            .CO(n28828));
    SB_LUT4 rem_4_add_1117_9_lut (.I0(GND_net), .I1(n1652_adj_4531), .I2(VCC_net), 
            .I3(n29082), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_9 (.CI(n29082), .I0(n1652_adj_4531), .I1(VCC_net), 
            .CO(n29083));
    SB_LUT4 div_46_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4589), .I3(n28826), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2257_8 (.CI(n28329), .I0(n1170), .I1(n94), .CO(n28330));
    SB_LUT4 add_2257_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n28328), 
            .O(n5819)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_8_lut (.I0(GND_net), .I1(n1653_adj_4532), .I2(VCC_net), 
            .I3(n29081), .O(n1720)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2257_7 (.CI(n28328), .I0(n1171), .I1(n95), .CO(n28329));
    SB_LUT4 add_2257_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n28327), 
            .O(n5820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2257_6 (.CI(n28327), .I0(n1172), .I1(n96), .CO(n28328));
    SB_LUT4 add_2257_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n28326), 
            .O(n5821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_8 (.CI(n28826), .I0(GND_net), .I1(n19_adj_4589), 
            .CO(n28827));
    SB_LUT4 div_46_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4590), .I3(n28825), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2257_5 (.CI(n28326), .I0(n1173), .I1(n97), .CO(n28327));
    SB_CARRY rem_4_add_1117_8 (.CI(n29081), .I0(n1653_adj_4532), .I1(VCC_net), 
            .CO(n29082));
    SB_CARRY div_46_unary_minus_4_add_3_7 (.CI(n28825), .I0(GND_net), .I1(n20_adj_4590), 
            .CO(n28826));
    SB_LUT4 rem_4_add_1117_7_lut (.I0(GND_net), .I1(n1654), .I2(GND_net), 
            .I3(n29080), .O(n1721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_7 (.CI(n29080), .I0(n1654), .I1(GND_net), 
            .CO(n29081));
    SB_LUT4 i12601_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n13195), .I3(GND_net), .O(n17283));   // verilog/coms.v(126[12] 289[6])
    defparam i12601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4591), .I3(n28824), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2257_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n28325), 
            .O(n5822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_6 (.CI(n28824), .I0(GND_net), .I1(n21_adj_4591), 
            .CO(n28825));
    SB_CARRY add_2257_4 (.CI(n28325), .I0(n1174), .I1(n98), .CO(n28326));
    SB_LUT4 add_2257_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n28324), 
            .O(n5823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12602_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n13195), .I3(GND_net), .O(n17284));   // verilog/coms.v(126[12] 289[6])
    defparam i12602_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2257_3 (.CI(n28324), .I0(n1175), .I1(n99), .CO(n28325));
    SB_LUT4 add_2257_2_lut (.I0(GND_net), .I1(n654), .I2(n558), .I3(VCC_net), 
            .O(n5824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2257_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_6_lut (.I0(GND_net), .I1(n1655), .I2(GND_net), 
            .I3(n29079), .O(n1722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_6 (.CI(n29079), .I0(n1655), .I1(GND_net), 
            .CO(n29080));
    SB_LUT4 div_46_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4592), .I3(n28823), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_5 (.CI(n28823), .I0(GND_net), .I1(n22_adj_4592), 
            .CO(n28824));
    SB_CARRY add_2257_2 (.CI(VCC_net), .I0(n654), .I1(n558), .CO(n28324));
    SB_LUT4 i12864_3_lut (.I0(encoder1_position[21]), .I1(n2893), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17546));   // quad.v(35[10] 41[6])
    defparam i12864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2256_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n28323), 
            .O(n5808)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2256_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12863_3_lut (.I0(encoder1_position[20]), .I1(n2894), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17545));   // quad.v(35[10] 41[6])
    defparam i12863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_5_lut (.I0(GND_net), .I1(n1656), .I2(VCC_net), 
            .I3(n29078), .O(n1723)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4593), .I3(n28822), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2256_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n28322), 
            .O(n5809)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2256_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2256_7 (.CI(n28322), .I0(n1044), .I1(n95), .CO(n28323));
    SB_LUT4 i12862_3_lut (.I0(encoder1_position[19]), .I1(n2895), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17544));   // quad.v(35[10] 41[6])
    defparam i12862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2256_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n28321), 
            .O(n5810)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2256_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12861_3_lut (.I0(encoder1_position[18]), .I1(n2896), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17543));   // quad.v(35[10] 41[6])
    defparam i12861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12603_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n13195), .I3(GND_net), .O(n17285));   // verilog/coms.v(126[12] 289[6])
    defparam i12603_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1117_5 (.CI(n29078), .I0(n1656), .I1(VCC_net), 
            .CO(n29079));
    SB_CARRY div_46_unary_minus_4_add_3_4 (.CI(n28822), .I0(GND_net), .I1(n23_adj_4593), 
            .CO(n28823));
    SB_CARRY add_2256_6 (.CI(n28321), .I0(n1045), .I1(n96), .CO(n28322));
    SB_LUT4 add_2256_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n28320), 
            .O(n5811)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2256_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2256_5 (.CI(n28320), .I0(n1046), .I1(n97), .CO(n28321));
    SB_LUT4 add_2256_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n28319), 
            .O(n5812)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2256_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12860_3_lut (.I0(encoder1_position[17]), .I1(n2897), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n17542));   // quad.v(35[10] 41[6])
    defparam i12860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_4_lut (.I0(GND_net), .I1(n1657), .I2(VCC_net), 
            .I3(n29077), .O(n1724)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4594), .I3(n28821), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2256_4 (.CI(n28319), .I0(n1047), .I1(n98), .CO(n28320));
    SB_LUT4 i22_3_lut_adj_1721 (.I0(bit_ctr[21]), .I1(n40182), .I2(n4385), 
            .I3(GND_net), .O(n33351));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1721.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1117_4 (.CI(n29077), .I0(n1657), .I1(VCC_net), 
            .CO(n29078));
    SB_CARRY div_46_unary_minus_4_add_3_3 (.CI(n28821), .I0(GND_net), .I1(n24_adj_4594), 
            .CO(n28822));
    SB_LUT4 rem_4_add_1117_3_lut (.I0(GND_net), .I1(n1658), .I2(GND_net), 
            .I3(n29076), .O(n1725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4595), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2256_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n28318), 
            .O(n5813)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2256_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2256_3 (.CI(n28318), .I0(n1048), .I1(n99), .CO(n28319));
    SB_LUT4 add_2256_2_lut (.I0(GND_net), .I1(n653), .I2(n558), .I3(VCC_net), 
            .O(n5814)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2256_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_782_3_lut (.I0(GND_net), .I1(n1157), .I2(VCC_net), 
            .I3(n27974), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_3 (.CI(n29076), .I0(n1658), .I1(GND_net), 
            .CO(n29077));
    SB_CARRY div_46_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4595), 
            .CO(n28821));
    SB_CARRY rem_4_add_782_3 (.CI(n27974), .I0(n1157), .I1(VCC_net), .CO(n27975));
    SB_LUT4 i12604_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n13195), .I3(GND_net), .O(n17286));   // verilog/coms.v(126[12] 289[6])
    defparam i12604_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2256_2 (.CI(VCC_net), .I0(n653), .I1(n558), .CO(n28318));
    SB_LUT4 rem_4_add_782_2_lut (.I0(GND_net), .I1(n1158), .I2(GND_net), 
            .I3(VCC_net), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2255_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n28317), 
            .O(n5800)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2255_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2255_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n28316), 
            .O(n5801)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2255_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2255_6 (.CI(n28316), .I0(n915), .I1(n96), .CO(n28317));
    SB_LUT4 add_2255_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n28315), 
            .O(n5802)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2255_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2255_5 (.CI(n28315), .I0(n916), .I1(n97), .CO(n28316));
    SB_LUT4 add_2255_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n28314), 
            .O(n5803)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2255_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2255_4 (.CI(n28314), .I0(n917), .I1(n98), .CO(n28315));
    SB_CARRY rem_4_add_1117_2 (.CI(VCC_net), .I0(n1758_adj_4498), .I1(VCC_net), 
            .CO(n29076));
    SB_LUT4 rem_4_add_1921_27_lut (.I0(n2867), .I1(n2834), .I2(VCC_net), 
            .I3(n28820), .O(n2933)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_782_2 (.CI(VCC_net), .I0(n1158), .I1(GND_net), 
            .CO(n27974));
    SB_LUT4 rem_4_add_1184_16_lut (.I0(n1778_adj_4500), .I1(n1745), .I2(VCC_net), 
            .I3(n29075), .O(n1844)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1921_26_lut (.I0(GND_net), .I1(n2835), .I2(VCC_net), 
            .I3(n28819), .O(n2902_adj_4473)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_15_lut (.I0(GND_net), .I1(n1746), .I2(VCC_net), 
            .I3(n29074), .O(n1813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_26 (.CI(n28819), .I0(n2835), .I1(VCC_net), 
            .CO(n28820));
    SB_LUT4 add_2255_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n28313), 
            .O(n5804)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2255_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2255_3 (.CI(n28313), .I0(n918), .I1(n99), .CO(n28314));
    SB_LUT4 add_2255_2_lut (.I0(GND_net), .I1(n652), .I2(n558), .I3(VCC_net), 
            .O(n5805)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2255_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2255_2 (.CI(VCC_net), .I0(n652), .I1(n558), .CO(n28313));
    SB_LUT4 rem_4_add_1921_25_lut (.I0(GND_net), .I1(n2836), .I2(VCC_net), 
            .I3(n28818), .O(n2903_adj_4472)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_15 (.CI(n29074), .I0(n1746), .I1(VCC_net), 
            .CO(n29075));
    SB_CARRY rem_4_add_1921_25 (.CI(n28818), .I0(n2836), .I1(VCC_net), 
            .CO(n28819));
    SB_LUT4 rem_4_add_1184_14_lut (.I0(GND_net), .I1(n1747), .I2(VCC_net), 
            .I3(n29073), .O(n1814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_24_lut (.I0(GND_net), .I1(n2837), .I2(VCC_net), 
            .I3(n28817), .O(n2904_adj_4471)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_14 (.CI(n29073), .I0(n1747), .I1(VCC_net), 
            .CO(n29074));
    SB_CARRY rem_4_add_1921_24 (.CI(n28817), .I0(n2837), .I1(VCC_net), 
            .CO(n28818));
    GND i1 (.Y(GND_net));
    SB_LUT4 rem_4_add_1184_13_lut (.I0(GND_net), .I1(n1748), .I2(VCC_net), 
            .I3(n29072), .O(n1815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_23_lut (.I0(GND_net), .I1(n2838), .I2(VCC_net), 
            .I3(n28816), .O(n2905_adj_4470)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12477_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17159));   // verilog/coms.v(126[12] 289[6])
    defparam i12477_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_13 (.CI(n29072), .I0(n1748), .I1(VCC_net), 
            .CO(n29073));
    SB_LUT4 i12478_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17160));   // verilog/coms.v(126[12] 289[6])
    defparam i12478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1184_12_lut (.I0(GND_net), .I1(n1749), .I2(VCC_net), 
            .I3(n29071), .O(n1816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_23 (.CI(n28816), .I0(n2838), .I1(VCC_net), 
            .CO(n28817));
    SB_LUT4 rem_4_add_1921_22_lut (.I0(GND_net), .I1(n2839), .I2(VCC_net), 
            .I3(n28815), .O(n2906_adj_4319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_12 (.CI(n29071), .I0(n1749), .I1(VCC_net), 
            .CO(n29072));
    SB_LUT4 rem_4_add_1184_11_lut (.I0(GND_net), .I1(n1750), .I2(VCC_net), 
            .I3(n29070), .O(n1817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_22 (.CI(n28815), .I0(n2839), .I1(VCC_net), 
            .CO(n28816));
    SB_LUT4 rem_4_add_1921_21_lut (.I0(GND_net), .I1(n2840), .I2(VCC_net), 
            .I3(n28814), .O(n2907_adj_4451)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_11 (.CI(n29070), .I0(n1750), .I1(VCC_net), 
            .CO(n29071));
    SB_LUT4 i12479_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17161));   // verilog/coms.v(126[12] 289[6])
    defparam i12479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12480_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17162));   // verilog/coms.v(126[12] 289[6])
    defparam i12480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12481_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17163));   // verilog/coms.v(126[12] 289[6])
    defparam i12481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12482_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17164));   // verilog/coms.v(126[12] 289[6])
    defparam i12482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12483_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n13195), .I3(GND_net), .O(n17165));   // verilog/coms.v(126[12] 289[6])
    defparam i12483_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_21 (.CI(n28814), .I0(n2840), .I1(VCC_net), 
            .CO(n28815));
    SB_LUT4 rem_4_add_1184_10_lut (.I0(GND_net), .I1(n1751), .I2(VCC_net), 
            .I3(n29069), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12605_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n13195), .I3(GND_net), .O(n17287));   // verilog/coms.v(126[12] 289[6])
    defparam i12605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12487_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n13195), .I3(GND_net), .O(n17169));   // verilog/coms.v(126[12] 289[6])
    defparam i12487_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_10 (.CI(n29069), .I0(n1751), .I1(VCC_net), 
            .CO(n29070));
    SB_LUT4 rem_4_add_1921_20_lut (.I0(GND_net), .I1(n2841), .I2(VCC_net), 
            .I3(n28813), .O(n2908_adj_4450)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_9_lut (.I0(GND_net), .I1(n1752), .I2(VCC_net), 
            .I3(n29068), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_20 (.CI(n28813), .I0(n2841), .I1(VCC_net), 
            .CO(n28814));
    SB_LUT4 i22_3_lut_adj_1722 (.I0(bit_ctr[14]), .I1(n40181), .I2(n4385), 
            .I3(GND_net), .O(n33349));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1722.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1184_9 (.CI(n29068), .I0(n1752), .I1(VCC_net), 
            .CO(n29069));
    SB_LUT4 rem_4_add_1921_19_lut (.I0(GND_net), .I1(n2842), .I2(VCC_net), 
            .I3(n28812), .O(n2909_adj_4449)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33843_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24853), .I3(start), .O(n40201));
    defparam i33843_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 rem_4_add_1184_8_lut (.I0(GND_net), .I1(n1753), .I2(VCC_net), 
            .I3(n29067), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_19 (.CI(n28812), .I0(n2842), .I1(VCC_net), 
            .CO(n28813));
    SB_LUT4 rem_4_add_1921_18_lut (.I0(GND_net), .I1(n2843), .I2(VCC_net), 
            .I3(n28811), .O(n2910_adj_4448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12488_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n13195), .I3(GND_net), .O(n17170));   // verilog/coms.v(126[12] 289[6])
    defparam i12488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_33_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(n2_adj_4965), .I3(n29951), .O(n746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_unary_minus_2_add_3_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4966), .I3(n29950), .O(n3_adj_4514)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_8 (.CI(n29067), .I0(n1753), .I1(VCC_net), 
            .CO(n29068));
    SB_LUT4 i2_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24853), .I3(state[1]), .O(n36917));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 rem_4_add_1184_7_lut (.I0(GND_net), .I1(n1754_adj_4494), .I2(GND_net), 
            .I3(n29066), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_18 (.CI(n28811), .I0(n2843), .I1(VCC_net), 
            .CO(n28812));
    SB_LUT4 i22_3_lut_adj_1723 (.I0(bit_ctr[13]), .I1(n40180), .I2(n4385), 
            .I3(GND_net), .O(n33347));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1723.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_32 (.CI(n29950), .I0(GND_net), .I1(n3_adj_4966), 
            .CO(n29951));
    SB_CARRY rem_4_add_1184_7 (.CI(n29066), .I0(n1754_adj_4494), .I1(GND_net), 
            .CO(n29067));
    SB_LUT4 i12489_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n13195), .I3(GND_net), .O(n17171));   // verilog/coms.v(126[12] 289[6])
    defparam i12489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1184_6_lut (.I0(GND_net), .I1(n1755_adj_4495), .I2(GND_net), 
            .I3(n29065), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_17_lut (.I0(GND_net), .I1(n2844), .I2(VCC_net), 
            .I3(n28810), .O(n2911_adj_4447)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_6 (.CI(n29065), .I0(n1755_adj_4495), .I1(GND_net), 
            .CO(n29066));
    SB_CARRY rem_4_add_1921_17 (.CI(n28810), .I0(n2844), .I1(VCC_net), 
            .CO(n28811));
    SB_LUT4 rem_4_add_1184_5_lut (.I0(GND_net), .I1(n1756_adj_4496), .I2(VCC_net), 
            .I3(n29064), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_5 (.CI(n29064), .I0(n1756_adj_4496), .I1(VCC_net), 
            .CO(n29065));
    SB_LUT4 rem_4_add_1921_16_lut (.I0(GND_net), .I1(n2845), .I2(VCC_net), 
            .I3(n28809), .O(n2912_adj_4446)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_16 (.CI(n28809), .I0(n2845), .I1(VCC_net), 
            .CO(n28810));
    SB_LUT4 rem_4_unary_minus_2_add_3_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4967), .I3(n29949), .O(n4_adj_4513)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_4_lut (.I0(GND_net), .I1(n1757_adj_4497), .I2(VCC_net), 
            .I3(n29063), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_31 (.CI(n29949), .I0(GND_net), .I1(n4_adj_4967), 
            .CO(n29950));
    SB_LUT4 rem_4_add_1921_15_lut (.I0(GND_net), .I1(n2846), .I2(VCC_net), 
            .I3(n28808), .O(n2913_adj_4445)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4968), .I3(n29948), .O(n5_adj_4512)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_30 (.CI(n29948), .I0(GND_net), .I1(n5_adj_4968), 
            .CO(n29949));
    SB_LUT4 rem_4_unary_minus_2_add_3_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4969), .I3(n29947), .O(n6_adj_4511)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_29 (.CI(n29947), .I0(GND_net), .I1(n6_adj_4969), 
            .CO(n29948));
    SB_LUT4 rem_4_unary_minus_2_add_3_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4970), .I3(n29946), .O(n7_adj_4510)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_28 (.CI(n29946), .I0(GND_net), .I1(n7_adj_4970), 
            .CO(n29947));
    SB_LUT4 rem_4_unary_minus_2_add_3_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4971), .I3(n29945), .O(n8_adj_4509)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1724 (.I0(n1746), .I1(n1747), .I2(n1745), .I3(n1748), 
            .O(n16_adj_4412));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i6_4_lut_adj_1724.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_unary_minus_2_add_3_27 (.CI(n29945), .I0(GND_net), .I1(n8_adj_4971), 
            .CO(n29946));
    SB_LUT4 rem_4_unary_minus_2_add_3_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4972), .I3(n29944), .O(n9_adj_4508)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_26 (.CI(n29944), .I0(GND_net), .I1(n9_adj_4972), 
            .CO(n29945));
    SB_LUT4 rem_4_unary_minus_2_add_3_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4973), .I3(n29943), .O(n10_adj_4507)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_25 (.CI(n29943), .I0(GND_net), .I1(n10_adj_4973), 
            .CO(n29944));
    SB_CARRY rem_4_add_1184_4 (.CI(n29063), .I0(n1757_adj_4497), .I1(VCC_net), 
            .CO(n29064));
    SB_LUT4 rem_4_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4974), .I3(n29942), .O(n11_adj_4506)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_24 (.CI(n29942), .I0(GND_net), .I1(n11_adj_4974), 
            .CO(n29943));
    SB_CARRY rem_4_add_1921_15 (.CI(n28808), .I0(n2846), .I1(VCC_net), 
            .CO(n28809));
    SB_LUT4 rem_4_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4975), .I3(n29941), .O(n12_adj_4505)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_23 (.CI(n29941), .I0(GND_net), .I1(n12_adj_4975), 
            .CO(n29942));
    SB_LUT4 rem_4_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4976), .I3(n29940), .O(n13_adj_4504)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_14_lut (.I0(GND_net), .I1(n2847), .I2(VCC_net), 
            .I3(n28807), .O(n2914_adj_4444)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_3_lut (.I0(GND_net), .I1(n1758_adj_4498), .I2(GND_net), 
            .I3(n29062), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_22 (.CI(n29940), .I0(GND_net), .I1(n13_adj_4976), 
            .CO(n29941));
    SB_LUT4 rem_4_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4977), .I3(n29939), .O(n14_adj_4469)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_14 (.CI(n28807), .I0(n2847), .I1(VCC_net), 
            .CO(n28808));
    SB_CARRY rem_4_unary_minus_2_add_3_21 (.CI(n29939), .I0(GND_net), .I1(n14_adj_4977), 
            .CO(n29940));
    SB_CARRY rem_4_add_1184_3 (.CI(n29062), .I0(n1758_adj_4498), .I1(GND_net), 
            .CO(n29063));
    SB_LUT4 rem_4_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4978), .I3(n29938), .O(n15_adj_4468)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_20 (.CI(n29938), .I0(GND_net), .I1(n15_adj_4978), 
            .CO(n29939));
    SB_LUT4 rem_4_add_1921_13_lut (.I0(GND_net), .I1(n2848), .I2(VCC_net), 
            .I3(n28806), .O(n2915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4979), .I3(n29937), .O(n16_adj_4467)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1725 (.I0(n1756_adj_4496), .I1(n1757_adj_4497), 
            .I2(n1758_adj_4498), .I3(GND_net), .O(n35564));
    defparam i1_3_lut_adj_1725.LUT_INIT = 16'hfefe;
    SB_CARRY rem_4_unary_minus_2_add_3_19 (.CI(n29937), .I0(GND_net), .I1(n16_adj_4979), 
            .CO(n29938));
    SB_LUT4 rem_4_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4980), .I3(n29936), .O(n17_adj_4466)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_2 (.CI(VCC_net), .I0(n1858), .I1(VCC_net), 
            .CO(n29062));
    SB_CARRY rem_4_add_1921_13 (.CI(n28806), .I0(n2848), .I1(VCC_net), 
            .CO(n28807));
    SB_LUT4 i8_3_lut (.I0(n1753), .I1(n16_adj_4412), .I2(n1751), .I3(GND_net), 
            .O(n18_adj_4411));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_1251_17_lut (.I0(n1844), .I1(n1844), .I2(n1877), 
            .I3(n29061), .O(n1943)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_1921_12_lut (.I0(GND_net), .I1(n2849), .I2(VCC_net), 
            .I3(n28805), .O(n2916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1726 (.I0(n1754_adj_4494), .I1(n1749), .I2(n35564), 
            .I3(n1755_adj_4495), .O(n13_adj_4413));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i3_4_lut_adj_1726.LUT_INIT = 16'heccc;
    SB_LUT4 i22_3_lut_adj_1727 (.I0(bit_ctr[12]), .I1(n40179), .I2(n4385), 
            .I3(GND_net), .O(n33343));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1727.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_unary_minus_2_add_3_18 (.CI(n29936), .I0(GND_net), .I1(n17_adj_4980), 
            .CO(n29937));
    SB_LUT4 rem_4_add_1251_16_lut (.I0(n1845), .I1(n1845), .I2(n1877), 
            .I3(n29060), .O(n1944)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4981), .I3(n29935), .O(n18_adj_4465)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_12 (.CI(n28805), .I0(n2849), .I1(VCC_net), 
            .CO(n28806));
    SB_CARRY rem_4_unary_minus_2_add_3_17 (.CI(n29935), .I0(GND_net), .I1(n18_adj_4981), 
            .CO(n29936));
    SB_LUT4 rem_4_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4982), .I3(n29934), .O(n19_adj_4464)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_16 (.CI(n29934), .I0(GND_net), .I1(n19_adj_4982), 
            .CO(n29935));
    SB_LUT4 rem_4_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4983), .I3(n29933), .O(n20_adj_4463)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_15 (.CI(n29933), .I0(GND_net), .I1(n20_adj_4983), 
            .CO(n29934));
    SB_LUT4 rem_4_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4984), .I3(n29932), .O(n21_adj_4462)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_14 (.CI(n29932), .I0(GND_net), .I1(n21_adj_4984), 
            .CO(n29933));
    SB_LUT4 rem_4_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4985), .I3(n29931), .O(n22_adj_4461)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_13 (.CI(n29931), .I0(GND_net), .I1(n22_adj_4985), 
            .CO(n29932));
    SB_LUT4 rem_4_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4986), .I3(n29930), .O(n23_adj_4460)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_12 (.CI(n29930), .I0(GND_net), .I1(n23_adj_4986), 
            .CO(n29931));
    SB_LUT4 rem_4_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4987), .I3(n29929), .O(n24_adj_4459)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_11 (.CI(n29929), .I0(GND_net), .I1(n24_adj_4987), 
            .CO(n29930));
    SB_LUT4 rem_4_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4988), .I3(n29928), .O(n25_adj_4458)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_10 (.CI(n29928), .I0(GND_net), .I1(n25_adj_4988), 
            .CO(n29929));
    SB_LUT4 rem_4_add_1921_11_lut (.I0(GND_net), .I1(n2850), .I2(VCC_net), 
            .I3(n28804), .O(n2917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26_adj_4989), .I3(n29927), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_9 (.CI(n29927), .I0(GND_net), .I1(n26_adj_4989), 
            .CO(n29928));
    SB_LUT4 rem_4_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n27_adj_4990), .I3(n29926), .O(n27_adj_4457)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_8 (.CI(n29926), .I0(GND_net), .I1(n27_adj_4990), 
            .CO(n29927));
    SB_LUT4 rem_4_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n28_adj_4991), .I3(n29925), .O(n28_adj_4456)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_7 (.CI(n29925), .I0(GND_net), .I1(n28_adj_4991), 
            .CO(n29926));
    SB_LUT4 rem_4_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n29_adj_4992), .I3(n29924), .O(n29_adj_4455)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_6 (.CI(n29924), .I0(GND_net), .I1(n29_adj_4992), 
            .CO(n29925));
    SB_CARRY rem_4_add_1251_16 (.CI(n29060), .I0(n1845), .I1(n1877), .CO(n29061));
    SB_LUT4 rem_4_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n30_adj_4993), .I3(n29923), .O(n30_adj_4454)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_11 (.CI(n28804), .I0(n2850), .I1(VCC_net), 
            .CO(n28805));
    SB_CARRY rem_4_unary_minus_2_add_3_5 (.CI(n29923), .I0(GND_net), .I1(n30_adj_4993), 
            .CO(n29924));
    SB_LUT4 rem_4_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n31_adj_4994), .I3(n29922), .O(n31_adj_4453)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_10_lut (.I0(n1283), .I1(n1250), .I2(VCC_net), 
            .I3(n28258), .O(n1349)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_unary_minus_2_add_3_4 (.CI(n29922), .I0(GND_net), .I1(n31_adj_4994), 
            .CO(n29923));
    SB_LUT4 rem_4_add_1251_15_lut (.I0(n1846), .I1(n1846), .I2(n1877), 
            .I3(n29059), .O(n1945)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n32_adj_4995), .I3(n29921), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_3 (.CI(n29921), .I0(GND_net), .I1(n32_adj_4995), 
            .CO(n29922));
    SB_LUT4 rem_4_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n33_adj_4996), .I3(VCC_net), .O(n33_adj_4452)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_10_lut (.I0(GND_net), .I1(n2851), .I2(VCC_net), 
            .I3(n28803), .O(n2918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n33_adj_4996), 
            .CO(n29921));
    SB_LUT4 rem_4_add_849_9_lut (.I0(GND_net), .I1(n1251), .I2(VCC_net), 
            .I3(n28257), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12490_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n13195), .I3(GND_net), .O(n17172));   // verilog/coms.v(126[12] 289[6])
    defparam i12490_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF blink_53 (.Q(blink), .C(LED_c), .D(blink_N_255));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    SB_CARRY rem_4_add_1921_10 (.CI(n28803), .I0(n2851), .I1(VCC_net), 
            .CO(n28804));
    SB_CARRY rem_4_add_1251_15 (.CI(n29059), .I0(n1846), .I1(n1877), .CO(n29060));
    SB_CARRY rem_4_add_849_9 (.CI(n28257), .I0(n1251), .I1(VCC_net), .CO(n28258));
    SB_LUT4 rem_4_add_1921_9_lut (.I0(GND_net), .I1(n2852), .I2(VCC_net), 
            .I3(n28802), .O(n2919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_14_lut (.I0(n1847), .I1(n1847), .I2(n1877), 
            .I3(n29058), .O(n1946)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_849_8_lut (.I0(GND_net), .I1(n1252), .I2(VCC_net), 
            .I3(n28256), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_9 (.CI(n28802), .I0(n2852), .I1(VCC_net), 
            .CO(n28803));
    SB_CARRY rem_4_add_849_8 (.CI(n28256), .I0(n1252), .I1(VCC_net), .CO(n28257));
    SB_LUT4 rem_4_add_1921_8_lut (.I0(GND_net), .I1(n2853), .I2(VCC_net), 
            .I3(n28801), .O(n2920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_7_lut (.I0(GND_net), .I1(n1253), .I2(VCC_net), 
            .I3(n28255), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_14 (.CI(n29058), .I0(n1847), .I1(n1877), .CO(n29059));
    SB_CARRY rem_4_add_1921_8 (.CI(n28801), .I0(n2853), .I1(VCC_net), 
            .CO(n28802));
    SB_CARRY rem_4_add_849_7 (.CI(n28255), .I0(n1253), .I1(VCC_net), .CO(n28256));
    SB_LUT4 rem_4_add_1251_13_lut (.I0(n1848), .I1(n1848), .I2(n1877), 
            .I3(n29057), .O(n1947)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_849_6_lut (.I0(GND_net), .I1(n1254), .I2(GND_net), 
            .I3(n28254), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_7_lut (.I0(GND_net), .I1(n2854), .I2(GND_net), 
            .I3(n28800), .O(n2921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_13 (.CI(n29057), .I0(n1848), .I1(n1877), .CO(n29058));
    SB_CARRY rem_4_add_849_6 (.CI(n28254), .I0(n1254), .I1(GND_net), .CO(n28255));
    SB_CARRY rem_4_add_1921_7 (.CI(n28800), .I0(n2854), .I1(GND_net), 
            .CO(n28801));
    SB_LUT4 i12491_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n13195), .I3(GND_net), .O(n17173));   // verilog/coms.v(126[12] 289[6])
    defparam i12491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12492_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n13195), .I3(GND_net), .O(n17174));   // verilog/coms.v(126[12] 289[6])
    defparam i12492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1251_12_lut (.I0(n1849), .I1(n1849), .I2(n1877), 
            .I3(n29056), .O(n1948)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1251_12 (.CI(n29056), .I0(n1849), .I1(n1877), .CO(n29057));
    SB_LUT4 rem_4_add_1921_6_lut (.I0(GND_net), .I1(n2855_adj_4474), .I2(GND_net), 
            .I3(n28799), .O(n2922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_5_lut (.I0(GND_net), .I1(n1255), .I2(GND_net), 
            .I3(n28253), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_6 (.CI(n28799), .I0(n2855_adj_4474), .I1(GND_net), 
            .CO(n28800));
    SB_LUT4 rem_4_add_1251_11_lut (.I0(n1850), .I1(n1850), .I2(n1877), 
            .I3(n29055), .O(n1949)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY rem_4_add_1251_11 (.CI(n29055), .I0(n1850), .I1(n1877), .CO(n29056));
    SB_CARRY rem_4_add_849_5 (.CI(n28253), .I0(n1255), .I1(GND_net), .CO(n28254));
    SB_LUT4 rem_4_add_1251_10_lut (.I0(n1851), .I1(n1851), .I2(n1877), 
            .I3(n29054), .O(n1950)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 rem_4_add_849_4_lut (.I0(GND_net), .I1(n1256), .I2(VCC_net), 
            .I3(n28252), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_5_lut (.I0(GND_net), .I1(n2856), .I2(VCC_net), 
            .I3(n28798), .O(n2923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_4 (.CI(n28252), .I0(n1256), .I1(VCC_net), .CO(n28253));
    SB_LUT4 rem_4_add_849_3_lut (.I0(GND_net), .I1(n1257), .I2(VCC_net), 
            .I3(n28251), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_10 (.CI(n29054), .I0(n1851), .I1(n1877), .CO(n29055));
    SB_CARRY rem_4_add_849_3 (.CI(n28251), .I0(n1257), .I1(VCC_net), .CO(n28252));
    SB_CARRY rem_4_add_1921_5 (.CI(n28798), .I0(n2856), .I1(VCC_net), 
            .CO(n28799));
    SB_LUT4 rem_4_add_849_2_lut (.I0(GND_net), .I1(n1258), .I2(GND_net), 
            .I3(VCC_net), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_2 (.CI(VCC_net), .I0(n1258), .I1(GND_net), 
            .CO(n28251));
    SB_LUT4 rem_4_add_1921_4_lut (.I0(GND_net), .I1(n2857), .I2(VCC_net), 
            .I3(n28797), .O(n2924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_9_lut (.I0(n1852), .I1(n1852), .I2(n1877), 
            .I3(n29053), .O(n1951)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12606_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n13195), .I3(GND_net), .O(n17288));   // verilog/coms.v(126[12] 289[6])
    defparam i12606_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_4 (.CI(n28797), .I0(n2857), .I1(VCC_net), 
            .CO(n28798));
    SB_CARRY rem_4_add_1251_9 (.CI(n29053), .I0(n1852), .I1(n1877), .CO(n29054));
    SB_LUT4 rem_4_add_1921_3_lut (.I0(GND_net), .I1(n2858), .I2(GND_net), 
            .I3(n28796), .O(n2925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_8_lut (.I0(n1853), .I1(n1853), .I2(n1877), 
            .I3(n29052), .O(n1952)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12493_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n13195), .I3(GND_net), .O(n17175));   // verilog/coms.v(126[12] 289[6])
    defparam i12493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12494_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n13195), .I3(GND_net), .O(n17176));   // verilog/coms.v(126[12] 289[6])
    defparam i12494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12495_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n13195), .I3(GND_net), .O(n17177));   // verilog/coms.v(126[12] 289[6])
    defparam i12495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12496_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n13195), .I3(GND_net), .O(n17178));   // verilog/coms.v(126[12] 289[6])
    defparam i12496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12497_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n13195), .I3(GND_net), .O(n17179));   // verilog/coms.v(126[12] 289[6])
    defparam i12497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12498_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n13195), .I3(GND_net), .O(n17180));   // verilog/coms.v(126[12] 289[6])
    defparam i12498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12499_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n13195), .I3(GND_net), .O(n17181));   // verilog/coms.v(126[12] 289[6])
    defparam i12499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12500_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n13195), .I3(GND_net), .O(n17182));   // verilog/coms.v(126[12] 289[6])
    defparam i12500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12501_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n13195), .I3(GND_net), .O(n17183));   // verilog/coms.v(126[12] 289[6])
    defparam i12501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12502_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n13195), .I3(GND_net), .O(n17184));   // verilog/coms.v(126[12] 289[6])
    defparam i12502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12503_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n13195), .I3(GND_net), .O(n17185));   // verilog/coms.v(126[12] 289[6])
    defparam i12503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12504_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n13195), .I3(GND_net), .O(n17186));   // verilog/coms.v(126[12] 289[6])
    defparam i12504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12505_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n13195), .I3(GND_net), .O(n17187));   // verilog/coms.v(126[12] 289[6])
    defparam i12505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12506_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n13195), .I3(GND_net), .O(n17188));   // verilog/coms.v(126[12] 289[6])
    defparam i12506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12507_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n13195), .I3(GND_net), .O(n17189));   // verilog/coms.v(126[12] 289[6])
    defparam i12507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4400));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4399));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4331));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12508_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n13195), .I3(GND_net), .O(n17190));   // verilog/coms.v(126[12] 289[6])
    defparam i12508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4398));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23126_2_lut_3_lut (.I0(n749), .I1(n855), .I2(n748), .I3(GND_net), 
            .O(n6_adj_4410));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i23126_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i585_3_lut_4_lut (.I0(n749), .I1(n855), .I2(n884), .I3(n748), 
            .O(n955));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i585_3_lut_4_lut.LUT_INIT = 16'hef10;
    SB_LUT4 i12320_4_lut (.I0(n16746), .I1(r_Bit_Index[2]), .I2(n4591), 
            .I3(n16635), .O(n17002));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12320_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4397));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4396));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4330));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4395));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12607_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n13195), .I3(GND_net), .O(n17289));   // verilog/coms.v(126[12] 289[6])
    defparam i12607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4364));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1596_3_lut (.I0(n2347), .I1(n2414), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2446));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1591_3_lut (.I0(n2342), .I1(n2409), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2441));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1598_3_lut (.I0(n2349), .I1(n2416), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2448_adj_4570));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1602_3_lut (.I0(n2353), .I1(n2420), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2452_adj_4566));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1599_3_lut (.I0(n2350), .I1(n2417), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2449_adj_4569));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1590_3_lut (.I0(n2341), .I1(n2408), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2440));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1601_3_lut (.I0(n2352), .I1(n2419), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2451_adj_4567));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1600_3_lut (.I0(n2351), .I1(n2418), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2450_adj_4568));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1594_3_lut (.I0(n2345), .I1(n2412), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2444));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1597_3_lut (.I0(n2348), .I1(n2415), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2447_adj_4571));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1607_3_lut (.I0(n2358_adj_4622), .I1(n2425), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2457_adj_4561));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1605_3_lut (.I0(n2356), .I1(n2423), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2455_adj_4563));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1604_3_lut (.I0(n2355), .I1(n2422), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2454_adj_4564));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1592_3_lut (.I0(n2343), .I1(n2410), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2442));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1589_3_lut (.I0(n2340), .I1(n2407), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2439));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1603_3_lut (.I0(n2354), .I1(n2421), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2453_adj_4565));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1595_3_lut (.I0(n2346), .I1(n2413), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2445));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1593_3_lut (.I0(n2344), .I1(n2411), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2443));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1606_3_lut (.I0(n2357_adj_4623), .I1(n2424), .I2(n2372_adj_4620), 
            .I3(GND_net), .O(n2456_adj_4562));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1728 (.I0(n2443), .I1(n2445), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4350));
    defparam i1_2_lut_adj_1728.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1729 (.I0(n2456_adj_4562), .I1(n2458_adj_4560), 
            .I2(GND_net), .I3(GND_net), .O(n37950));
    defparam i1_2_lut_adj_1729.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n2454_adj_4564), .I1(n37950), .I2(n2455_adj_4563), 
            .I3(n2457_adj_4561), .O(n35665));
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'ha080;
    SB_LUT4 i13_4_lut_adj_1731 (.I0(n2453_adj_4565), .I1(n2439), .I2(n2442), 
            .I3(n18_adj_4350), .O(n30_adj_4347));
    defparam i13_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1732 (.I0(n2447_adj_4571), .I1(n2444), .I2(n2450_adj_4568), 
            .I3(n2451_adj_4567), .O(n28_adj_4349));
    defparam i11_4_lut_adj_1732.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1733 (.I0(n35665), .I1(n2440), .I2(n2449_adj_4569), 
            .I3(n2452_adj_4566), .O(n29_adj_4348));
    defparam i12_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1734 (.I0(n2448_adj_4570), .I1(n2438), .I2(n2441), 
            .I3(n2446), .O(n27));
    defparam i10_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1735 (.I0(n27), .I1(n29_adj_4348), .I2(n28_adj_4349), 
            .I3(n30_adj_4347), .O(n2471_adj_4558));
    defparam i16_4_lut_adj_1735.LUT_INIT = 16'hfffe;
    SB_LUT4 i12509_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n13195), .I3(GND_net), .O(n17191));   // verilog/coms.v(126[12] 289[6])
    defparam i12509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12510_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n13195), .I3(GND_net), .O(n17192));   // verilog/coms.v(126[12] 289[6])
    defparam i12510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12511_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n13195), .I3(GND_net), .O(n17193));   // verilog/coms.v(126[12] 289[6])
    defparam i12511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12512_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n13195), .I3(GND_net), .O(n17194));   // verilog/coms.v(126[12] 289[6])
    defparam i12512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12513_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n13195), .I3(GND_net), .O(n17195));   // verilog/coms.v(126[12] 289[6])
    defparam i12513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12514_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n13195), .I3(GND_net), .O(n17196));   // verilog/coms.v(126[12] 289[6])
    defparam i12514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12515_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n13195), .I3(GND_net), .O(n17197));   // verilog/coms.v(126[12] 289[6])
    defparam i12515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i12_3_lut (.I0(communication_counter[11]), .I1(n22_adj_4461), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2458_adj_4560));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12516_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n13195), .I3(GND_net), .O(n17198));   // verilog/coms.v(126[12] 289[6])
    defparam i12516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12517_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n13195), .I3(GND_net), .O(n17199));   // verilog/coms.v(126[12] 289[6])
    defparam i12517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12518_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n13195), .I3(GND_net), .O(n17200));   // verilog/coms.v(126[12] 289[6])
    defparam i12518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12519_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n13195), .I3(GND_net), .O(n17201));   // verilog/coms.v(126[12] 289[6])
    defparam i12519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12520_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n13195), .I3(GND_net), .O(n17202));   // verilog/coms.v(126[12] 289[6])
    defparam i12520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12521_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n13195), .I3(GND_net), .O(n17203));   // verilog/coms.v(126[12] 289[6])
    defparam i12521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12522_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n13195), .I3(GND_net), .O(n17204));   // verilog/coms.v(126[12] 289[6])
    defparam i12522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12523_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n13195), .I3(GND_net), .O(n17205));   // verilog/coms.v(126[12] 289[6])
    defparam i12523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12524_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n13195), .I3(GND_net), .O(n17206));   // verilog/coms.v(126[12] 289[6])
    defparam i12524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12525_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n13195), .I3(GND_net), .O(n17207));   // verilog/coms.v(126[12] 289[6])
    defparam i12525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12526_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n13195), .I3(GND_net), .O(n17208));   // verilog/coms.v(126[12] 289[6])
    defparam i12526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12608_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n13195), .I3(GND_net), .O(n17290));   // verilog/coms.v(126[12] 289[6])
    defparam i12608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4365));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12527_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n13195), .I3(GND_net), .O(n17209));   // verilog/coms.v(126[12] 289[6])
    defparam i12527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12528_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n13195), .I3(GND_net), .O(n17210));   // verilog/coms.v(126[12] 289[6])
    defparam i12528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12529_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n13195), .I3(GND_net), .O(n17211));   // verilog/coms.v(126[12] 289[6])
    defparam i12529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12530_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n13195), .I3(GND_net), .O(n17212));   // verilog/coms.v(126[12] 289[6])
    defparam i12530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12531_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n13195), .I3(GND_net), .O(n17213));   // verilog/coms.v(126[12] 289[6])
    defparam i12531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12532_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n13195), .I3(GND_net), .O(n17214));   // verilog/coms.v(126[12] 289[6])
    defparam i12532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12533_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n13195), .I3(GND_net), .O(n17215));   // verilog/coms.v(126[12] 289[6])
    defparam i12533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34115_3_lut_3_lut (.I0(n392), .I1(n558), .I2(n369), .I3(GND_net), 
            .O(n510));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34115_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i12534_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n13195), .I3(GND_net), .O(n17216));   // verilog/coms.v(126[12] 289[6])
    defparam i12534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12535_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n13195), .I3(GND_net), .O(n17217));   // verilog/coms.v(126[12] 289[6])
    defparam i12535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12536_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n13195), .I3(GND_net), .O(n17218));   // verilog/coms.v(126[12] 289[6])
    defparam i12536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12537_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n13195), .I3(GND_net), .O(n17219));   // verilog/coms.v(126[12] 289[6])
    defparam i12537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12538_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n13195), .I3(GND_net), .O(n17220));   // verilog/coms.v(126[12] 289[6])
    defparam i12538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12539_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n13195), .I3(GND_net), .O(n17221));   // verilog/coms.v(126[12] 289[6])
    defparam i12539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12540_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n13195), .I3(GND_net), .O(n17222));   // verilog/coms.v(126[12] 289[6])
    defparam i12540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12541_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n13195), .I3(GND_net), .O(n17223));   // verilog/coms.v(126[12] 289[6])
    defparam i12541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12542_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n13195), .I3(GND_net), .O(n17224));   // verilog/coms.v(126[12] 289[6])
    defparam i12542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12543_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n13195), .I3(GND_net), .O(n17225));   // verilog/coms.v(126[12] 289[6])
    defparam i12543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12544_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n13195), .I3(GND_net), .O(n17226));   // verilog/coms.v(126[12] 289[6])
    defparam i12544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12545_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n13195), .I3(GND_net), .O(n17227));   // verilog/coms.v(126[12] 289[6])
    defparam i12545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12546_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n13195), .I3(GND_net), .O(n17228));   // verilog/coms.v(126[12] 289[6])
    defparam i12546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12547_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n13195), .I3(GND_net), .O(n17229));   // verilog/coms.v(126[12] 289[6])
    defparam i12547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12548_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n13195), .I3(GND_net), .O(n17230));   // verilog/coms.v(126[12] 289[6])
    defparam i12548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12549_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n13195), .I3(GND_net), .O(n17231));   // verilog/coms.v(126[12] 289[6])
    defparam i12549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12550_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n13195), .I3(GND_net), .O(n17232));   // verilog/coms.v(126[12] 289[6])
    defparam i12550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12551_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n13195), .I3(GND_net), .O(n17233));   // verilog/coms.v(126[12] 289[6])
    defparam i12551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12552_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n13195), .I3(GND_net), .O(n17234));   // verilog/coms.v(126[12] 289[6])
    defparam i12552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12553_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n13195), .I3(GND_net), .O(n17235));   // verilog/coms.v(126[12] 289[6])
    defparam i12553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12554_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n13195), .I3(GND_net), .O(n17236));   // verilog/coms.v(126[12] 289[6])
    defparam i12554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12555_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n13195), .I3(GND_net), .O(n17237));   // verilog/coms.v(126[12] 289[6])
    defparam i12555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4413), .I1(n18_adj_4411), .I2(n1752), 
            .I3(n1750), .O(n1778_adj_4500));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12556_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n13195), .I3(GND_net), .O(n17238));   // verilog/coms.v(126[12] 289[6])
    defparam i12556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12557_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n13195), .I3(GND_net), .O(n17239));   // verilog/coms.v(126[12] 289[6])
    defparam i12557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4329));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12558_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n13195), .I3(GND_net), .O(n17240));   // verilog/coms.v(126[12] 289[6])
    defparam i12558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12609_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n13195), .I3(GND_net), .O(n17291));   // verilog/coms.v(126[12] 289[6])
    defparam i12609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12559_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n13195), .I3(GND_net), .O(n17241));   // verilog/coms.v(126[12] 289[6])
    defparam i12559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12560_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n13195), .I3(GND_net), .O(n17242));   // verilog/coms.v(126[12] 289[6])
    defparam i12560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12561_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n13195), .I3(GND_net), .O(n17243));   // verilog/coms.v(126[12] 289[6])
    defparam i12561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12562_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n13195), .I3(GND_net), .O(n17244));   // verilog/coms.v(126[12] 289[6])
    defparam i12562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12563_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n13195), .I3(GND_net), .O(n17245));   // verilog/coms.v(126[12] 289[6])
    defparam i12563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4366));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12564_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n13195), .I3(GND_net), .O(n17246));   // verilog/coms.v(126[12] 289[6])
    defparam i12564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12565_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n13195), .I3(GND_net), .O(n17247));   // verilog/coms.v(126[12] 289[6])
    defparam i12565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12566_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n13195), 
            .I3(GND_net), .O(n17248));   // verilog/coms.v(126[12] 289[6])
    defparam i12566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12567_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n13195), 
            .I3(GND_net), .O(n17249));   // verilog/coms.v(126[12] 289[6])
    defparam i12567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12568_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n13195), 
            .I3(GND_net), .O(n17250));   // verilog/coms.v(126[12] 289[6])
    defparam i12568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12569_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n13195), 
            .I3(GND_net), .O(n17251));   // verilog/coms.v(126[12] 289[6])
    defparam i12569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12570_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n13195), 
            .I3(GND_net), .O(n17252));   // verilog/coms.v(126[12] 289[6])
    defparam i12570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12571_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n13195), 
            .I3(GND_net), .O(n17253));   // verilog/coms.v(126[12] 289[6])
    defparam i12571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12572_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n13195), 
            .I3(GND_net), .O(n17254));   // verilog/coms.v(126[12] 289[6])
    defparam i12572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12573_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n13195), 
            .I3(GND_net), .O(n17255));   // verilog/coms.v(126[12] 289[6])
    defparam i12573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12610_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n13195), .I3(GND_net), .O(n17292));   // verilog/coms.v(126[12] 289[6])
    defparam i12610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i891_3_lut_3_lut (.I0(n1316), .I1(n5835), .I2(n655), 
            .I3(GND_net), .O(n1420));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i891_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12574_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n13195), 
            .I3(GND_net), .O(n17256));   // verilog/coms.v(126[12] 289[6])
    defparam i12574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12575_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n13195), 
            .I3(GND_net), .O(n17257));   // verilog/coms.v(126[12] 289[6])
    defparam i12575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12576_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n13195), 
            .I3(GND_net), .O(n17258));   // verilog/coms.v(126[12] 289[6])
    defparam i12576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12577_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n13195), 
            .I3(GND_net), .O(n17259));   // verilog/coms.v(126[12] 289[6])
    defparam i12577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12578_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n13195), 
            .I3(GND_net), .O(n17260));   // verilog/coms.v(126[12] 289[6])
    defparam i12578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12579_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n13195), 
            .I3(GND_net), .O(n17261));   // verilog/coms.v(126[12] 289[6])
    defparam i12579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12580_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n13195), 
            .I3(GND_net), .O(n17262));   // verilog/coms.v(126[12] 289[6])
    defparam i12580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12581_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n13195), 
            .I3(GND_net), .O(n17263));   // verilog/coms.v(126[12] 289[6])
    defparam i12581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12582_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n13195), 
            .I3(GND_net), .O(n17264));   // verilog/coms.v(126[12] 289[6])
    defparam i12582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12323_4_lut (.I0(n16746), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n16635), .O(n17005));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12323_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i22_3_lut_adj_1736 (.I0(bit_ctr[20]), .I1(n40178), .I2(n4385), 
            .I3(GND_net), .O(n33341));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1736.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2_adj_4630), 
            .I3(n5_adj_4925), .O(n35307));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1120_3_lut (.I0(n1647_adj_4526), .I1(n1714), .I2(n1679), 
            .I3(GND_net), .O(n1746));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1187_3_lut (.I0(n1746), .I1(n1813), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12583_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n13195), 
            .I3(GND_net), .O(n17265));   // verilog/coms.v(126[12] 289[6])
    defparam i12583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1194_3_lut (.I0(n1753), .I1(n1820), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12584_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n13195), 
            .I3(GND_net), .O(n17266));   // verilog/coms.v(126[12] 289[6])
    defparam i12584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34092_3_lut_3_lut (.I0(n533), .I1(n558), .I2(n511), .I3(GND_net), 
            .O(n649));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34092_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 unary_minus_28_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4328));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4327));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1524_3_lut (.I0(n2243), .I1(n2310), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2342));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35135_3_lut (.I0(n1653_adj_4532), .I1(n1720), .I2(n1679), 
            .I3(GND_net), .O(n1752));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1523_3_lut (.I0(n2242), .I1(n2309), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2341));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35136_3_lut (.I0(n1752), .I1(n1819), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1522_3_lut (.I0(n2241), .I1(n2308), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2340));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1191_3_lut (.I0(n1750), .I1(n1817), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35065_3_lut (.I0(n2150), .I1(n2217), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2249));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34845_3_lut (.I0(n2249), .I1(n2316), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2348));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35087_3_lut (.I0(n2151), .I1(n2218), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2250));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34843_3_lut (.I0(n2250), .I1(n2317), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2349));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1528_3_lut (.I0(n2247), .I1(n2314), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2346));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1533_3_lut (.I0(n2252), .I1(n2319), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2351));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1534_3_lut (.I0(n2253), .I1(n2320), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2352));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1532_3_lut (.I0(n2251), .I1(n2318), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2350));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1529_3_lut (.I0(n2248), .I1(n2315), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2347));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1535_3_lut (.I0(n2254), .I1(n2321), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2353));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1526_3_lut (.I0(n2245), .I1(n2312), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2344));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1527_3_lut (.I0(n2246), .I1(n2313), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2345));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1525_3_lut (.I0(n2244), .I1(n2311), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2343));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1539_3_lut (.I0(n2258), .I1(n2325), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2357_adj_4623));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1537_3_lut (.I0(n2256), .I1(n2323), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2355));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1536_3_lut (.I0(n2255), .I1(n2322), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2354));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1538_3_lut (.I0(n2257), .I1(n2324), .I2(n2273_adj_4629), 
            .I3(GND_net), .O(n2356));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1737 (.I0(n2356), .I1(n2358_adj_4622), .I2(GND_net), 
            .I3(GND_net), .O(n37700));
    defparam i1_2_lut_adj_1737.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n2354), .I1(n37700), .I2(n2355), .I3(n2357_adj_4623), 
            .O(n35597));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'ha080;
    SB_LUT4 i12_4_lut_adj_1739 (.I0(n2353), .I1(n2347), .I2(n2350), .I3(n2352), 
            .O(n28_adj_5010));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1740 (.I0(n2343), .I1(n2345), .I2(n2344), .I3(n35597), 
            .O(n26_adj_5012));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1740.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1190_3_lut (.I0(n1749), .I1(n1816), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1741 (.I0(n2351), .I1(n2346), .I2(n2349), .I3(n2348), 
            .O(n27_adj_5011));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1742 (.I0(n2340), .I1(n2341), .I2(n2339), .I3(n2342), 
            .O(n25_adj_5013));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1743 (.I0(n25_adj_5013), .I1(n27_adj_5011), .I2(n26_adj_5012), 
            .I3(n28_adj_5010), .O(n2372_adj_4620));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i15_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i13_3_lut (.I0(communication_counter[12]), .I1(n21_adj_4462), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2358_adj_4622));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4326));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(171[23:28])
    defparam unary_minus_28_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12585_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n13195), 
            .I3(GND_net), .O(n17267));   // verilog/coms.v(126[12] 289[6])
    defparam i12585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i4_3_lut (.I0(communication_counter[3]), .I1(n30_adj_4454), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3258));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12586_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n13195), 
            .I3(GND_net), .O(n17268));   // verilog/coms.v(126[12] 289[6])
    defparam i12586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12587_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n13195), 
            .I3(GND_net), .O(n17269));   // verilog/coms.v(126[12] 289[6])
    defparam i12587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4369));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1189_3_lut (.I0(n1748), .I1(n1815), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1744 (.I0(blink), .I1(n15_adj_4338), .I2(GND_net), 
            .I3(GND_net), .O(blink_N_255));
    defparam i1_2_lut_adj_1744.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i368_4_lut_4_lut (.I0(n533), .I1(n99), .I2(n2), .I3(n510), 
            .O(n648));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i368_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4370));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4371));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1467_3_lut (.I0(n2154), .I1(n2221), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2253));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1459_3_lut (.I0(n2146), .I1(n2213), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2245));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1457_3_lut (.I0(n2144), .I1(n2211), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2243));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1458_3_lut (.I0(n2145), .I1(n2212), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2244));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1456_3_lut (.I0(n2143), .I1(n2210), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2242));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1469_3_lut (.I0(n2156), .I1(n2223), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2255));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1468_3_lut (.I0(n2155), .I1(n2222), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2254));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1460_3_lut (.I0(n2147), .I1(n2214), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2246));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i1_1_lut (.I0(communication_counter[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_4996));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i2_1_lut (.I0(communication_counter[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_4995));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i3_1_lut (.I0(communication_counter[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_4994));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i4_1_lut (.I0(communication_counter[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_4993));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i5_1_lut (.I0(communication_counter[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_4992));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1461_3_lut (.I0(n2148), .I1(n2215), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2247));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i6_1_lut (.I0(communication_counter[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_4991));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1455_3_lut (.I0(n2142), .I1(n2209), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2241));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i7_1_lut (.I0(communication_counter[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_4990));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i8_1_lut (.I0(communication_counter[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_4989));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i9_1_lut (.I0(communication_counter[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4988));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i10_1_lut (.I0(communication_counter[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4987));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34848_3_lut (.I0(n2053), .I1(n2120), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2152));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34849_3_lut (.I0(n2152), .I1(n2219), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2251));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i11_1_lut (.I0(communication_counter[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4986));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1466_3_lut (.I0(n2153), .I1(n2220), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2252));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34854_3_lut (.I0(n2050), .I1(n2117), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2149));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i12_1_lut (.I0(communication_counter[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4985));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34855_3_lut (.I0(n2149), .I1(n2216), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2248));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i34855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i13_1_lut (.I0(communication_counter[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4984));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1471_3_lut (.I0(n2158), .I1(n2225), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2257));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1470_3_lut (.I0(n2157), .I1(n2224), .I2(n2174_adj_4638), 
            .I3(GND_net), .O(n2256));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1745 (.I0(n2256), .I1(n2257), .I2(n2258), .I3(GND_net), 
            .O(n35660));
    defparam i1_3_lut_adj_1745.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1746 (.I0(n2248), .I1(n2252), .I2(n2251), .I3(n2249), 
            .O(n26_adj_4524));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i11_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1747 (.I0(n2246), .I1(n2254), .I2(n35660), .I3(n2255), 
            .O(n19_adj_4621));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1747.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1748 (.I0(n2241), .I1(n2240), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4625));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_adj_1748.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1749 (.I0(n2242), .I1(n2244), .I2(n2243), .I3(n2245), 
            .O(n24_adj_4535));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i9_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1750 (.I0(n19_adj_4621), .I1(n26_adj_4524), .I2(n2247), 
            .I3(n2250), .O(n28_adj_4515));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1750.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1751 (.I0(n2253), .I1(n28_adj_4515), .I2(n24_adj_4535), 
            .I3(n16_adj_4625), .O(n2273_adj_4629));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i14_3_lut (.I0(communication_counter[13]), .I1(n20_adj_4463), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2258));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i14_1_lut (.I0(communication_counter[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4983));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4380));   // verilog/TinyFPGA_B.v(250[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i15_1_lut (.I0(communication_counter[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4982));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i16_1_lut (.I0(communication_counter[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4981));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i17_1_lut (.I0(communication_counter[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4980));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i18_1_lut (.I0(communication_counter[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4979));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i19_1_lut (.I0(communication_counter[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4978));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i20_1_lut (.I0(communication_counter[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4977));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i21_1_lut (.I0(communication_counter[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4976));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i22_1_lut (.I0(communication_counter[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4975));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i23_1_lut (.I0(communication_counter[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4974));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i24_1_lut (.I0(communication_counter[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4973));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i25_1_lut (.I0(communication_counter[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4972));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i26_1_lut (.I0(communication_counter[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4971));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i27_1_lut (.I0(communication_counter[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4970));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i28_1_lut (.I0(communication_counter[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4969));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i29_1_lut (.I0(communication_counter[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4968));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i30_1_lut (.I0(communication_counter[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4967));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2076_3_lut (.I0(n3051), .I1(n3118), .I2(n3065), .I3(GND_net), 
            .O(n3150));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2078_3_lut (.I0(n3053), .I1(n3120), .I2(n3065), .I3(GND_net), 
            .O(n3152));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2068_3_lut (.I0(n3043), .I1(n3110), .I2(n3065), .I3(GND_net), 
            .O(n3142));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2075_3_lut (.I0(n3050), .I1(n3117), .I2(n3065), .I3(GND_net), 
            .O(n3149));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2058_3_lut (.I0(n3033), .I1(n3100), .I2(n3065), .I3(GND_net), 
            .O(n3132));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2079_3_lut (.I0(n3054), .I1(n3121), .I2(n3065), .I3(GND_net), 
            .O(n3153));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2073_3_lut (.I0(n3048), .I1(n3115), .I2(n3065), .I3(GND_net), 
            .O(n3147));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2070_3_lut (.I0(n3045), .I1(n3112), .I2(n3065), .I3(GND_net), 
            .O(n3144));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2069_3_lut (.I0(n3044), .I1(n3111), .I2(n3065), .I3(GND_net), 
            .O(n3143));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2066_3_lut (.I0(n3041), .I1(n3108), .I2(n3065), .I3(GND_net), 
            .O(n3140));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2065_3_lut (.I0(n3040), .I1(n3107), .I2(n3065), .I3(GND_net), 
            .O(n3139));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2064_3_lut (.I0(n3039), .I1(n3106), .I2(n3065), .I3(GND_net), 
            .O(n3138));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i31_1_lut (.I0(communication_counter[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4966));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2062_3_lut (.I0(n3037), .I1(n3104), .I2(n3065), .I3(GND_net), 
            .O(n3136));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1127_3_lut (.I0(n1654), .I1(n1721), .I2(n1679), .I3(GND_net), 
            .O(n1753));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2063_3_lut (.I0(n3038), .I1(n3105), .I2(n3065), .I3(GND_net), 
            .O(n3137));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2061_3_lut (.I0(n3036), .I1(n3103), .I2(n3065), .I3(GND_net), 
            .O(n3135));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2060_3_lut (.I0(n3035), .I1(n3102), .I2(n3065), .I3(GND_net), 
            .O(n3134));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2059_3_lut (.I0(n3034), .I1(n3101), .I2(n3065), .I3(GND_net), 
            .O(n3133));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2071_3_lut (.I0(n3046), .I1(n3113), .I2(n3065), .I3(GND_net), 
            .O(n3145));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2077_3_lut (.I0(n3052), .I1(n3119), .I2(n3065), .I3(GND_net), 
            .O(n3151));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2072_3_lut (.I0(n3047), .I1(n3114), .I2(n3065), .I3(GND_net), 
            .O(n3146));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2074_3_lut (.I0(n3049), .I1(n3116), .I2(n3065), .I3(GND_net), 
            .O(n3148));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2081_3_lut (.I0(n3056), .I1(n3123), .I2(n3065), .I3(GND_net), 
            .O(n3155));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35140_3_lut (.I0(n1652_adj_4531), .I1(n1719), .I2(n1679), 
            .I3(GND_net), .O(n1751));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12279_3_lut (.I0(gearBoxRatio[0]), .I1(\data_in_frame[19] [0]), 
            .I2(n36885), .I3(GND_net), .O(n16961));   // verilog/coms.v(126[12] 289[6])
    defparam i12279_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12280_3_lut (.I0(Kp[0]), .I1(\data_in_frame[2] [0]), .I2(n36885), 
            .I3(GND_net), .O(n16962));   // verilog/coms.v(126[12] 289[6])
    defparam i12280_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12281_3_lut (.I0(Ki[0]), .I1(\data_in_frame[3] [0]), .I2(n36885), 
            .I3(GND_net), .O(n16963));   // verilog/coms.v(126[12] 289[6])
    defparam i12281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2067_3_lut (.I0(n3042), .I1(n3109), .I2(n3065), .I3(GND_net), 
            .O(n3141));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12282_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n16964));   // verilog/coms.v(126[12] 289[6])
    defparam i12282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2080_3_lut (.I0(n3055), .I1(n3122), .I2(n3065), .I3(GND_net), 
            .O(n3154));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12283_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n36885), .I3(GND_net), .O(n16965));   // verilog/coms.v(126[12] 289[6])
    defparam i12283_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12285_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[7] [0]), 
            .I2(n36885), .I3(GND_net), .O(n16967));   // verilog/coms.v(126[12] 289[6])
    defparam i12285_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2083_3_lut (.I0(n3058), .I1(n3125), .I2(n3065), .I3(GND_net), 
            .O(n3157));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2082_3_lut (.I0(n3057), .I1(n3124), .I2(n3065), .I3(GND_net), 
            .O(n3156));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1752 (.I0(n3156), .I1(n3157), .I2(n3158), .I3(GND_net), 
            .O(n35642));
    defparam i1_3_lut_adj_1752.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1753 (.I0(n3154), .I1(n3141), .I2(n35642), .I3(n3155), 
            .O(n30_adj_4949));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i6_4_lut_adj_1753.LUT_INIT = 16'heccc;
    SB_LUT4 i16_4_lut_adj_1754 (.I0(n3148), .I1(n3146), .I2(n3151), .I3(n3145), 
            .O(n40_adj_4947));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i16_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(n3133), .I1(n3134), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_4950));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1755 (.I0(n3135), .I1(n3137), .I2(n3136), .I3(n3138), 
            .O(n38_adj_4948));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i14_4_lut_adj_1755.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1756 (.I0(n3139), .I1(n40_adj_4947), .I2(n30_adj_4949), 
            .I3(n3140), .O(n44_adj_4943));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i20_4_lut_adj_1756.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1757 (.I0(n3143), .I1(n3144), .I2(n3147), .I3(n3153), 
            .O(n42_adj_4945));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i18_4_lut_adj_1757.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1758 (.I0(n3132), .I1(n38_adj_4948), .I2(n26_adj_4950), 
            .I3(n3131), .O(n43_adj_4944));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i19_4_lut_adj_1758.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1759 (.I0(n3149), .I1(n3142), .I2(n3152), .I3(n3150), 
            .O(n41_adj_4946));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i17_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n41_adj_4946), .I1(n43_adj_4944), .I2(n42_adj_4945), 
            .I3(n44_adj_4943), .O(n3164));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12286_3_lut (.I0(encoder0_position[0]), .I1(n2964), .I2(count_enable), 
            .I3(GND_net), .O(n16968));   // quad.v(35[10] 41[6])
    defparam i12286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1760 (.I0(\FRAME_MATCHER.i_31__N_2386 ), .I1(\FRAME_MATCHER.i_31__N_2390 ), 
            .I2(n737), .I3(n2855), .O(n6));   // verilog/coms.v(126[12] 289[6])
    defparam i2_4_lut_adj_1760.LUT_INIT = 16'h0ace;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n5), .I1(\FRAME_MATCHER.state [0]), .I2(n6), 
            .I3(n10283), .O(n36_adj_5007));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hc8fa;
    SB_LUT4 i12588_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n13195), 
            .I3(GND_net), .O(n17270));   // verilog/coms.v(126[12] 289[6])
    defparam i12588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12589_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n13195), 
            .I3(GND_net), .O(n17271));   // verilog/coms.v(126[12] 289[6])
    defparam i12589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n34657), .I1(n36_adj_5007), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n18962), .O(n33975));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hccdc;
    SB_LUT4 i12288_3_lut (.I0(encoder1_position[0]), .I1(n2914), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n16970));   // quad.v(35[10] 41[6])
    defparam i12288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12289_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n37155), 
            .I3(GND_net), .O(n16971));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12289_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12611_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n13195), .I3(GND_net), .O(n17293));   // verilog/coms.v(126[12] 289[6])
    defparam i12611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1763 (.I0(bit_ctr[25]), .I1(n40186), .I2(n4385), 
            .I3(GND_net), .O(n33359));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1763.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1124_3_lut (.I0(n1651_adj_4530), .I1(n1718), .I2(n1679), 
            .I3(GND_net), .O(n1750));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1123_3_lut (.I0(n1650_adj_4529), .I1(n1717), .I2(n1679), 
            .I3(GND_net), .O(n1749));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1764 (.I0(bit_ctr[24]), .I1(n40185), .I2(n4385), 
            .I3(GND_net), .O(n33357));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1764.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i367_4_lut_4_lut (.I0(n533), .I1(n98), .I2(n4_adj_4394), 
            .I3(n35307), .O(n35315));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i367_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i22_3_lut_adj_1765 (.I0(bit_ctr[23]), .I1(n40184), .I2(n4385), 
            .I3(GND_net), .O(n33355));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1765.LUT_INIT = 16'hacac;
    SB_LUT4 i12612_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n13195), .I3(GND_net), .O(n17294));   // verilog/coms.v(126[12] 289[6])
    defparam i12612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1766 (.I0(bit_ctr[22]), .I1(n40183), .I2(n4385), 
            .I3(GND_net), .O(n33353));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1766.LUT_INIT = 16'hacac;
    SB_LUT4 i12297_3_lut (.I0(tx_o), .I1(n3_adj_4952), .I2(r_SM_Main_adj_5053[2]), 
            .I3(GND_net), .O(n16979));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12297_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12590_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n13195), .I3(GND_net), .O(n17272));   // verilog/coms.v(126[12] 289[6])
    defparam i12590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1122_3_lut (.I0(n1649_adj_4528), .I1(n1716), .I2(n1679), 
            .I3(GND_net), .O(n1748));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1392_3_lut (.I0(n2047), .I1(n2114), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2146));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1391_3_lut (.I0(n2046), .I1(n2113), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2145));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1767 (.I0(bit_ctr[31]), .I1(n40192), .I2(n4385), 
            .I3(GND_net), .O(n33371));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1767.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut (.I0(n852), .I1(n6_adj_4410), .I2(n746), .I3(GND_net), 
            .O(n884));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i28617_2_lut_3_lut (.I0(n852), .I1(n6_adj_4410), .I2(n746), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i28617_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i35233_3_lut (.I0(n1553_adj_4533), .I1(n1620), .I2(n1580), 
            .I3(GND_net), .O(n1652_adj_4531));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34089_3_lut_3_lut (.I0(n671), .I1(n558), .I2(n650), .I3(GND_net), 
            .O(n785));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34089_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 rem_4_i1399_3_lut (.I0(n2054), .I1(n2121), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2153));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12217_4_lut (.I0(n26602), .I1(r_Clock_Count_adj_5054[5]), .I2(n316), 
            .I3(r_SM_Main_adj_5053[2]), .O(n16899));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12217_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i12223_4_lut (.I0(n26602), .I1(r_Clock_Count_adj_5054[3]), .I2(n318), 
            .I3(r_SM_Main_adj_5053[2]), .O(n16905));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12223_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 rem_4_i1390_3_lut (.I0(n2045), .I1(n2112), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2144));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i458_4_lut_4_lut (.I0(n671), .I1(n97), .I2(n6_adj_4475), 
            .I3(n35315), .O(n35317));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i458_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1389_3_lut (.I0(n2044), .I1(n2111), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2143));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12299_4_lut (.I0(r_SM_Main_adj_5053[2]), .I1(n29), .I2(n26612), 
            .I3(r_SM_Main_adj_5053[0]), .O(n16981));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12299_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i3_2_lut_adj_1768 (.I0(color_23__N_164[3]), .I1(color_23__N_164[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4964));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i3_2_lut_adj_1768.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(color_23__N_164[4]), .I1(color_23__N_164[6]), 
            .I2(color_23__N_164[2]), .I3(color_23__N_164[0]), .O(n13_adj_4963));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(color_23__N_164[7]), .I1(n13_adj_4963), 
            .I2(n11_adj_4964), .I3(color_23__N_164[1]), .O(n15_adj_4338));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i460_4_lut_4_lut (.I0(n671), .I1(n99), .I2(n2_adj_4559), 
            .I3(n649), .O(n784));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i460_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i1_2_lut_adj_1771 (.I0(color_23__N_164[1]), .I1(blink), .I2(GND_net), 
            .I3(GND_net), .O(n37558));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_2_lut_adj_1771.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(color_23__N_164[7]), .I1(n13_adj_4963), 
            .I2(n11_adj_4964), .I3(n37558), .O(n16695));   // verilog/TinyFPGA_B.v(76[6:36])
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 i12880_3_lut (.I0(color[4]), .I1(n16695), .I2(n15_adj_4338), 
            .I3(GND_net), .O(n17562));   // verilog/TinyFPGA_B.v(73[8] 96[4])
    defparam i12880_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12300_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1169), .I3(GND_net), .O(n16982));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1388_3_lut (.I0(n2043), .I1(n2110), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2142));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1396_3_lut (.I0(n2051), .I1(n2118), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2150));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1397_3_lut (.I0(n2052), .I1(n2119), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2151));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1394_3_lut (.I0(n2049), .I1(n2116), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2148));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1401_3_lut (.I0(n2056), .I1(n2123), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2155));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1393_3_lut (.I0(n2048), .I1(n2115), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2147));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1400_3_lut (.I0(n2055), .I1(n2122), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2154));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1403_3_lut (.I0(n2058), .I1(n2125), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2157));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1402_3_lut (.I0(n2057), .I1(n2124), .I2(n2075_adj_4653), 
            .I3(GND_net), .O(n2156));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1773 (.I0(n2156), .I1(n2157), .I2(n2158), .I3(GND_net), 
            .O(n35585));
    defparam i1_3_lut_adj_1773.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1774 (.I0(n2154), .I1(n2147), .I2(n35585), .I3(n2155), 
            .O(n18_adj_4961));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i4_4_lut_adj_1774.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut_adj_1775 (.I0(n2148), .I1(n2151), .I2(n2149), .I3(n2150), 
            .O(n24_adj_4954));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i10_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1776 (.I0(n2142), .I1(n2143), .I2(n2141), .I3(n2144), 
            .O(n22_adj_4956));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i8_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1777 (.I0(n2145), .I1(n24_adj_4954), .I2(n18_adj_4961), 
            .I3(n2146), .O(n26_adj_4953));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i12_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1778 (.I0(n2152), .I1(n26_adj_4953), .I2(n22_adj_4956), 
            .I3(n2153), .O(n2174_adj_4638));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i13_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i15_3_lut (.I0(communication_counter[14]), .I1(n19_adj_4464), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2158));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12591_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n13195), .I3(GND_net), .O(n17273));   // verilog/coms.v(126[12] 289[6])
    defparam i12591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12304_3_lut (.I0(setpoint[0]), .I1(n4292), .I2(n36839), .I3(GND_net), 
            .O(n16986));   // verilog/coms.v(126[12] 289[6])
    defparam i12304_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12211_4_lut (.I0(n26602), .I1(r_Clock_Count_adj_5054[7]), .I2(n314), 
            .I3(r_SM_Main_adj_5053[2]), .O(n16893));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12211_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i12205_4_lut (.I0(n30_adj_4346), .I1(r_Clock_Count[1]), .I2(n225), 
            .I3(n3_adj_5009), .O(n16887));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12205_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i12208_4_lut (.I0(n26602), .I1(r_Clock_Count_adj_5054[8]), .I2(n313), 
            .I3(r_SM_Main_adj_5053[2]), .O(n16890));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12208_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i12199_4_lut (.I0(n30_adj_4346), .I1(r_Clock_Count[3]), .I2(n223), 
            .I3(n3_adj_5009), .O(n16881));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12199_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i35138_3_lut (.I0(n1751), .I1(n1818), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i35138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i28_3_lut (.I0(communication_counter[27]), .I1(n6_adj_4511), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n855));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1188_3_lut (.I0(n1747), .I1(n1814), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i29_3_lut (.I0(communication_counter[28]), .I1(n5_adj_4512), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n749));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i30_3_lut (.I0(communication_counter[29]), .I1(n4_adj_4513), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n748));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i652_3_lut (.I0(n955), .I1(n1022), .I2(n986), .I3(GND_net), 
            .O(n1054));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i719_3_lut (.I0(n1054), .I1(n1121), .I2(n1085), .I3(GND_net), 
            .O(n1153));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i786_3_lut (.I0(n1153), .I1(n1220), .I2(n1184), .I3(GND_net), 
            .O(n1252));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i853_3_lut (.I0(n1252), .I1(n1319), .I2(n1283), .I3(GND_net), 
            .O(n1351));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i920_3_lut (.I0(n1351), .I1(n1418_adj_4537), .I2(n1382), 
            .I3(GND_net), .O(n1450));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i987_3_lut (.I0(n1450), .I1(n1517), .I2(n1481), .I3(GND_net), 
            .O(n1549));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1054_3_lut (.I0(n1549), .I1(n1616), .I2(n1580), .I3(GND_net), 
            .O(n1648_adj_4527));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i459_4_lut_4_lut (.I0(n671), .I1(n98), .I2(n4_adj_4476), 
            .I3(n648), .O(n783));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i459_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i550_4_lut_4_lut (.I0(n806), .I1(n99), .I2(n2_adj_4342), 
            .I3(n785), .O(n917));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i550_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4640));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i12308_3_lut (.I0(quadB_debounced_adj_4373), .I1(reg_B_adj_5064[0]), 
            .I2(n36606), .I3(GND_net), .O(n16990));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4595));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1779 (.I0(control_mode[0]), .I1(n15508), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_4321));   // verilog/TinyFPGA_B.v(228[5:22])
    defparam i1_2_lut_3_lut_adj_1779.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4594));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1780 (.I0(control_mode[0]), .I1(n15508), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(228[5:22])
    defparam i1_2_lut_3_lut_adj_1780.LUT_INIT = 16'hefef;
    SB_LUT4 div_46_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4593));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4592));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4591));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1060_3_lut (.I0(n1555), .I1(n1622), .I2(n1580), .I3(GND_net), 
            .O(n1654));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4590));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1059_rep_25_3_lut (.I0(n1554_adj_4534), .I1(n1621), .I2(n1580), 
            .I3(GND_net), .O(n1653_adj_4532));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1059_rep_25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4589));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4588));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1057_3_lut (.I0(n1552), .I1(n1619), .I2(n1580), .I3(GND_net), 
            .O(n1651_adj_4530));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1056_3_lut (.I0(n1551), .I1(n1618), .I2(n1580), .I3(GND_net), 
            .O(n1650_adj_4529));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4587));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4586));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1055_3_lut (.I0(n1550), .I1(n1617), .I2(n1580), .I3(GND_net), 
            .O(n1649_adj_4528));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4585));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4584));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4583));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4582));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4581));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4580));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4579));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1781 (.I0(n1856), .I1(n1857), .I2(n1858), .I3(GND_net), 
            .O(n35596));
    defparam i1_3_lut_adj_1781.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i1121_3_lut (.I0(n1648_adj_4527), .I1(n1715), .I2(n1679), 
            .I3(GND_net), .O(n1747));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4578));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n1854), .I1(n1853), .I2(n35596), .I3(n1855), 
            .O(n12_adj_4353));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'heccc;
    SB_LUT4 rem_4_mux_3_i23_3_lut (.I0(communication_counter[22]), .I1(n11_adj_4506), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1358));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i993_3_lut (.I0(n1456), .I1(n1523), .I2(n1481), .I3(GND_net), 
            .O(n1555));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4577));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i992_3_lut (.I0(n1455), .I1(n1522), .I2(n1481), .I3(GND_net), 
            .O(n1554_adj_4534));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4576));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i991_rep_29_3_lut (.I0(n1454), .I1(n1521), .I2(n1481), 
            .I3(GND_net), .O(n1553_adj_4533));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i991_rep_29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4575));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i990_3_lut (.I0(n1453), .I1(n1520), .I2(n1481), .I3(GND_net), 
            .O(n1552));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4574));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4573));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i989_3_lut (.I0(n1452), .I1(n1519), .I2(n1481), .I3(GND_net), 
            .O(n1551));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4572));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i988_3_lut (.I0(n1451), .I1(n1518), .I2(n1481), .I3(GND_net), 
            .O(n1550));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4619));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12187_4_lut (.I0(n30_adj_4346), .I1(r_Clock_Count[7]), .I2(n219), 
            .I3(n3_adj_5009), .O(n16869));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12187_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4618));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1783 (.I0(n1849), .I1(n1847), .I2(n1848), .I3(n1851), 
            .O(n18_adj_4352));
    defparam i7_4_lut_adj_1783.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4617));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4616));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4615));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i927_3_lut (.I0(n1358), .I1(n1425), .I2(n1382), .I3(GND_net), 
            .O(n1457));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4614));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4613));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i926_3_lut (.I0(n1357), .I1(n1424), .I2(n1382), .I3(GND_net), 
            .O(n1456));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4612));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34083_3_lut_3_lut (.I0(n806), .I1(n558), .I2(n651), .I3(GND_net), 
            .O(n918));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34083_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 rem_4_i925_3_lut (.I0(n1356), .I1(n1423), .I2(n1382), .I3(GND_net), 
            .O(n1455));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4611));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4610));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i924_3_lut (.I0(n1355), .I1(n1422), .I2(n1382), .I3(GND_net), 
            .O(n1454));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4609));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i923_3_lut (.I0(n1354), .I1(n1421), .I2(n1382), .I3(GND_net), 
            .O(n1453));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4608));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i548_4_lut_4_lut (.I0(n806), .I1(n97), .I2(n6_adj_4323), 
            .I3(n783), .O(n915));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i548_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i549_4_lut_4_lut (.I0(n806), .I1(n98), .I2(n4_adj_4325), 
            .I3(n784), .O(n916));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i549_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i922_3_lut (.I0(n1353), .I1(n1420_adj_4539), .I2(n1382), 
            .I3(GND_net), .O(n1452));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i921_3_lut (.I0(n1352), .I1(n1419_adj_4538), .I2(n1382), 
            .I3(GND_net), .O(n1451));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4607));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4606));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4605));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4604));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4603));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12190_4_lut (.I0(n30_adj_4346), .I1(r_Clock_Count[6]), .I2(n220), 
            .I3(n3_adj_5009), .O(n16872));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12190_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i12896_3_lut (.I0(setpoint[5]), .I1(n4297), .I2(n36839), .I3(GND_net), 
            .O(n17578));   // verilog/coms.v(126[12] 289[6])
    defparam i12896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4602));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i547_4_lut_4_lut (.I0(n806), .I1(n96), .I2(n8), .I3(n35317), 
            .O(n914));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i547_4_lut_4_lut.LUT_INIT = 16'h14eb;
    SB_LUT4 i12895_3_lut (.I0(setpoint[4]), .I1(n4296), .I2(n36839), .I3(GND_net), 
            .O(n17577));   // verilog/coms.v(126[12] 289[6])
    defparam i12895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4601));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4600));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4599));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12894_3_lut (.I0(setpoint[3]), .I1(n4295), .I2(n36839), .I3(GND_net), 
            .O(n17576));   // verilog/coms.v(126[12] 289[6])
    defparam i12894_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12893_3_lut (.I0(setpoint[2]), .I1(n4294), .I2(n36839), .I3(GND_net), 
            .O(n17575));   // verilog/coms.v(126[12] 289[6])
    defparam i12893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12892_3_lut (.I0(setpoint[1]), .I1(n4293), .I2(n36839), .I3(GND_net), 
            .O(n17574));   // verilog/coms.v(126[12] 289[6])
    defparam i12892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4598));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4597));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12891_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1169), .I3(GND_net), .O(n17573));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12905_3_lut (.I0(setpoint[14]), .I1(n4306), .I2(n36839), 
            .I3(GND_net), .O(n17587));   // verilog/coms.v(126[12] 289[6])
    defparam i12905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4596));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    coms setpoint_23__I_0 (.\data_in_frame[1] ({\data_in_frame[1] }), .\data_in_frame[17] ({\data_in_frame[17] }), 
         .clk32MHz(clk32MHz), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .GND_net(GND_net), .\data_in_frame[5] ({\data_in_frame[5] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .rx_data({rx_data}), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n17581(n17581), .setpoint({setpoint}), .n17582(n17582), .n17583(n17583), 
         .n17584(n17584), .n17585(n17585), .n17586(n17586), .n17587(n17587), 
         .n17574(n17574), .n17575(n17575), .n17576(n17576), .n17577(n17577), 
         .n17578(n17578), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .n17595(n17595), .n17596(n17596), .n17593(n17593), .n17594(n17594), 
         .n17591(n17591), .n17592(n17592), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n17588(n17588), .n17589(n17589), .n17590(n17590), .n17579(n17579), 
         .n17580(n17580), .n17495(n17495), .PWMLimit({PWMLimit}), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n17496(n17496), .n17497(n17497), .n17498(n17498), .n17499(n17499), 
         .n17500(n17500), .n17501(n17501), .n17487(n17487), .n17488(n17488), 
         .n17489(n17489), .n17490(n17490), .n17491(n17491), .n17492(n17492), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .n43272(n43272), .\data_in_frame[19] ({\data_in_frame[19] }), 
         .\data_in_frame[18] ({\data_in_frame[18] }), .n17493(n17493), .n17494(n17494), 
         .n17479(n17479), .n17480(n17480), .n17481(n17481), .n17482(n17482), 
         .n17483(n17483), .n17484(n17484), .n17485(n17485), .n17486(n17486), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .n17303(n17303), 
         .control_mode({control_mode}), .n17302(n17302), .n17301(n17301), 
         .n17300(n17300), .n17299(n17299), .n17298(n17298), .n17297(n17297), 
         .n17295(n17295), .n17294(n17294), .n17293(n17293), .n17292(n17292), 
         .n17291(n17291), .n17290(n17290), .n17289(n17289), .n17288(n17288), 
         .n17287(n17287), .n17286(n17286), .n17285(n17285), .n17284(n17284), 
         .n17283(n17283), .n17282(n17282), .n17281(n17281), .n17280(n17280), 
         .n17279(n17279), .n17278(n17278), .rx_data_ready(rx_data_ready), 
         .n17277(n17277), .n17276(n17276), .n17275(n17275), .n17274(n17274), 
         .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), .n36839(n36839), 
         .n4300(n4300), .n17273(n17273), .n17272(n17272), .n17271(n17271), 
         .n17270(n17270), .\data_in_frame[8] ({\data_in_frame[8] }), .n17269(n17269), 
         .n17268(n17268), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .n17267(n17267), .n17266(n17266), .n17265(n17265), .n17264(n17264), 
         .n17263(n17263), .n17262(n17262), .n17261(n17261), .n17260(n17260), 
         .n17259(n17259), .n17258(n17258), .n17257(n17257), .n17256(n17256), 
         .n17255(n17255), .n34657(n34657), .n18962(n18962), .n63(n63), 
         .n17254(n17254), .n17253(n17253), .n17252(n17252), .n17251(n17251), 
         .n17250(n17250), .n17249(n17249), .n17248(n17248), .n17247(n17247), 
         .n17246(n17246), .n17245(n17245), .n17244(n17244), .n17243(n17243), 
         .n17242(n17242), .n17241(n17241), .n17240(n17240), .n17239(n17239), 
         .n17238(n17238), .n17237(n17237), .n17236(n17236), .n17235(n17235), 
         .n17234(n17234), .n17233(n17233), .n17232(n17232), .n17231(n17231), 
         .n17230(n17230), .n17229(n17229), .n17228(n17228), .n17227(n17227), 
         .n17226(n17226), .n17225(n17225), .n17224(n17224), .n17223(n17223), 
         .n17222(n17222), .n17221(n17221), .n17220(n17220), .n17219(n17219), 
         .n17218(n17218), .n17217(n17217), .n17216(n17216), .n17215(n17215), 
         .n17214(n17214), .n17213(n17213), .n17212(n17212), .n17211(n17211), 
         .n17210(n17210), .n17209(n17209), .n17208(n17208), .n17207(n17207), 
         .n17206(n17206), .n17205(n17205), .n17204(n17204), .n17203(n17203), 
         .n17202(n17202), .n17201(n17201), .n17200(n17200), .n17199(n17199), 
         .n17198(n17198), .n17197(n17197), .n17196(n17196), .n17195(n17195), 
         .n17194(n17194), .n17193(n17193), .n17192(n17192), .n17191(n17191), 
         .n17190(n17190), .n17189(n17189), .n17188(n17188), .n17187(n17187), 
         .n17186(n17186), .n17185(n17185), .n17184(n17184), .n17183(n17183), 
         .n17182(n17182), .n17181(n17181), .n17180(n17180), .n17179(n17179), 
         .n17178(n17178), .n17177(n17177), .n17176(n17176), .n17175(n17175), 
         .n17174(n17174), .n17173(n17173), .n17172(n17172), .n17171(n17171), 
         .n17170(n17170), .n17169(n17169), .n17165(n17165), .n17164(n17164), 
         .\data_in[3] ({\data_in[3] }), .n17163(n17163), .n17162(n17162), 
         .n17161(n17161), .n17160(n17160), .n17159(n17159), .n17158(n17158), 
         .n17157(n17157), .n17155(n17155), .\data_in[2][6] (\data_in[2] [6]), 
         .n17154(n17154), .\data_in[2][5] (\data_in[2] [5]), .n17153(n17153), 
         .\data_in[2][4] (\data_in[2] [4]), .\data_in[2][3] (\data_in[2] [3]), 
         .n17151(n17151), .\data_in[2][2] (\data_in[2] [2]), .\data_in[2][1] (\data_in[2] [1]), 
         .n17149(n17149), .\data_in[2][0] (\data_in[2] [0]), .n17147(n17147), 
         .\data_in[1][6] (\data_in[1] [6]), .n13195(n13195), .\data_in[0] ({Open_0, 
         Open_1, Open_2, Open_3, Open_4, \data_in[0] [2], Open_5, 
         Open_6}), .n17146(n17146), .\data_in[1][5] (\data_in[1] [5]), 
         .n737(n737), .\data_in[1][3] (\data_in[1] [3]), .\data_in[0][5] (\data_in[0] [5]), 
         .\data_in[1][2] (\data_in[1] [2]), .\data_in[0][1] (\data_in[0] [1]), 
         .n17145(n17145), .\data_in[1][4] (\data_in[1] [4]), .n17144(n17144), 
         .n17143(n17143), .\data_in[0][0] (\data_in[0] [0]), .\data_in[1][1] (\data_in[1] [1]), 
         .\data_in[0][4] (\data_in[0] [4]), .\data_in[0][3] (\data_in[0] [3]), 
         .\data_in[0][6] (\data_in[0] [6]), .\data_in[1][0] (\data_in[1] [0]), 
         .n17142(n17142), .n17141(n17141), .n17139(n17139), .n17138(n17138), 
         .\FRAME_MATCHER.i_31__N_2390 (\FRAME_MATCHER.i_31__N_2390 ), .n2855(n2855), 
         .n10283(n10283), .n17137(n17137), .n17136(n17136), .n17135(n17135), 
         .\FRAME_MATCHER.i_31__N_2386 (\FRAME_MATCHER.i_31__N_2386 ), .n122(n122), 
         .n17134(n17134), .n17133(n17133), .\Ki[7] (Ki[7]), .n17132(n17132), 
         .\Ki[6] (Ki[6]), .n17131(n17131), .\Ki[5] (Ki[5]), .n17130(n17130), 
         .\Ki[4] (Ki[4]), .n17129(n17129), .\Ki[3] (Ki[3]), .n8849(n8849), 
         .n17128(n17128), .\Ki[2] (Ki[2]), .n17127(n17127), .\Ki[1] (Ki[1]), 
         .n17126(n17126), .\Kp[7] (Kp[7]), .n17125(n17125), .\Kp[6] (Kp[6]), 
         .n17124(n17124), .\Kp[5] (Kp[5]), .n17123(n17123), .\Kp[4] (Kp[4]), 
         .n17122(n17122), .\Kp[3] (Kp[3]), .n17121(n17121), .\Kp[2] (Kp[2]), 
         .n17120(n17120), .\Kp[1] (Kp[1]), .n17119(n17119), .gearBoxRatio({gearBoxRatio}), 
         .n17118(n17118), .n17117(n17117), .n17116(n17116), .n4(n4_adj_5006), 
         .\FRAME_MATCHER.state_31__N_2426[2] (\FRAME_MATCHER.state_31__N_2426 [2]), 
         .n7(n7_adj_4477), .n17115(n17115), .n17114(n17114), .n17113(n17113), 
         .n17112(n17112), .n17111(n17111), .n17110(n17110), .n17109(n17109), 
         .n17108(n17108), .n17107(n17107), .n17106(n17106), .n17105(n17105), 
         .n17104(n17104), .n17103(n17103), .n17102(n17102), .n17101(n17101), 
         .n17100(n17100), .n17099(n17099), .n17098(n17098), .n17097(n17097), 
         .n17096(n17096), .IntegralLimit({IntegralLimit}), .n17095(n17095), 
         .n17094(n17094), .n17093(n17093), .n17092(n17092), .n17091(n17091), 
         .n17090(n17090), .n17089(n17089), .n17088(n17088), .n17087(n17087), 
         .n17086(n17086), .n17085(n17085), .n17084(n17084), .n17083(n17083), 
         .n17082(n17082), .n17081(n17081), .n17080(n17080), .n17079(n17079), 
         .n17078(n17078), .n17077(n17077), .n17076(n17076), .n17075(n17075), 
         .n17074(n17074), .n36885(n36885), .n4299(n4299), .n4298(n4298), 
         .n4309(n4309), .n4308(n4308), .n4307(n4307), .n4311(n4311), 
         .LED_c(LED_c), .n4310(n4310), .n4313(n4313), .n4312(n4312), 
         .n4315(n4315), .n4314(n4314), .n16832(n16832), .n16986(n16986), 
         .n33975(n33975), .n16967(n16967), .n16965(n16965), .n16964(n16964), 
         .n16963(n16963), .\Ki[0] (Ki[0]), .n16962(n16962), .\Kp[0] (Kp[0]), 
         .n16961(n16961), .n4292(n4292), .n4297(n4297), .n4296(n4296), 
         .n4295(n4295), .n4294(n4294), .n4293(n4293), .n4306(n4306), 
         .n4305(n4305), .n4304(n4304), .n4303(n4303), .n4302(n4302), 
         .n4301(n4301), .n5(n5), .n318(n318), .\r_Clock_Count[3] (r_Clock_Count_adj_5054[3]), 
         .n16918(n16918), .r_Bit_Index({r_Bit_Index_adj_5055}), .n16915(n16915), 
         .n16911(n16911), .\r_Clock_Count[1] (r_Clock_Count_adj_5054[1]), 
         .n16890(n16890), .\r_Clock_Count[8] (r_Clock_Count_adj_5054[8]), 
         .n16893(n16893), .\r_Clock_Count[7] (r_Clock_Count_adj_5054[7]), 
         .n16905(n16905), .n16899(n16899), .\r_Clock_Count[5] (r_Clock_Count_adj_5054[5]), 
         .n17029(n17029), .n17566(n17566), .r_SM_Main({r_SM_Main_adj_5053}), 
         .n26602(n26602), .n320(n320), .VCC_net(VCC_net), .n4613(n4613), 
         .n26612(n26612), .n16641(n16641), .n16772(n16772), .tx_o(tx_o), 
         .tx_enable(tx_enable), .n313(n313), .n314(n314), .n16981(n16981), 
         .n16979(n16979), .n316(n316), .n3(n3_adj_4952), .n29(n29), 
         .n16872(n16872), .\r_Clock_Count[6] (r_Clock_Count[6]), .n16869(n16869), 
         .\r_Clock_Count[7]_adj_3 (r_Clock_Count[7]), .n16881(n16881), .\r_Clock_Count[3]_adj_4 (r_Clock_Count[3]), 
         .n16887(n16887), .\r_Clock_Count[1]_adj_5 (r_Clock_Count[1]), .n17005(n17005), 
         .r_Bit_Index_adj_13({r_Bit_Index}), .n17002(n17002), .n17550(n17550), 
         .r_Rx_Data(r_Rx_Data), .PIN_13_N_105(PIN_13_N_105), .n219(n219), 
         .n220(n220), .n30(n30_adj_4346), .n223(n223), .n3_adj_9(n3_adj_5009), 
         .n225(n225), .n15459(n15459), .n4_adj_10(n4_adj_4379), .n16746(n16746), 
         .n16635(n16635), .n17012(n17012), .n17011(n17011), .n17010(n17010), 
         .n17009(n17009), .n17008(n17008), .n17007(n17007), .n17006(n17006), 
         .n4591(n4591), .n24014(n24014), .n4_adj_11(n4_adj_4375), .n4_adj_12(n4), 
         .n15454(n15454)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(202[8] 223[4])
    SB_LUT4 i12324_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n24014), 
            .I3(n15454), .O(n17006));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12324_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i12904_3_lut (.I0(setpoint[13]), .I1(n4305), .I2(n36839), 
            .I3(GND_net), .O(n17586));   // verilog/coms.v(126[12] 289[6])
    defparam i12904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12903_3_lut (.I0(setpoint[12]), .I1(n4304), .I2(n36839), 
            .I3(GND_net), .O(n17585));   // verilog/coms.v(126[12] 289[6])
    defparam i12903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12325_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n24014), 
            .I3(n15459), .O(n17007));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12325_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 div_46_i638_3_lut_3_lut (.I0(n938), .I1(n5804), .I2(n918), 
            .I3(GND_net), .O(n1047));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i638_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12902_3_lut (.I0(setpoint[11]), .I1(n4303), .I2(n36839), 
            .I3(GND_net), .O(n17584));   // verilog/coms.v(126[12] 289[6])
    defparam i12902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i639_3_lut_3_lut (.I0(n938), .I1(n5805), .I2(n652), 
            .I3(GND_net), .O(n1048));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i639_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12326_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4375), 
            .I3(n15454), .O(n17008));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12326_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12901_3_lut (.I0(setpoint[10]), .I1(n4302), .I2(n36839), 
            .I3(GND_net), .O(n17583));   // verilog/coms.v(126[12] 289[6])
    defparam i12901_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12327_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4375), 
            .I3(n15459), .O(n17009));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12327_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12328_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4), .I3(n15454), 
            .O(n17010));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12328_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12900_3_lut (.I0(setpoint[9]), .I1(n4301), .I2(n36839), .I3(GND_net), 
            .O(n17582));   // verilog/coms.v(126[12] 289[6])
    defparam i12900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12329_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4), .I3(n15459), 
            .O(n17011));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12329_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12330_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4379), 
            .I3(n15454), .O(n17012));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12330_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12335_4_lut (.I0(n16754), .I1(state[1]), .I2(state_3__N_362[1]), 
            .I3(n16530), .O(n17017));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12335_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i12149_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n37092), .I3(GND_net), .O(n16831));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i636_3_lut_3_lut (.I0(n938), .I1(n5802), .I2(n916), 
            .I3(GND_net), .O(n1045));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i636_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12150_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n36885), .I3(GND_net), .O(n16832));   // verilog/coms.v(126[12] 289[6])
    defparam i12150_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34074_2_lut (.I0(start), .I1(n24907), .I2(GND_net), .I3(GND_net), 
            .O(n40203));   // verilog/neopixel.v(35[12] 117[6])
    defparam i34074_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31_4_lut (.I0(n40203), .I1(n40201), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n33387));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 div_46_i635_3_lut_3_lut (.I0(n938), .I1(n5801), .I2(n915), 
            .I3(GND_net), .O(n1044));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i635_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i634_3_lut_3_lut (.I0(n938), .I1(n5800), .I2(n914), 
            .I3(GND_net), .O(n1043));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i634_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i24_3_lut (.I0(communication_counter[23]), .I1(n10_adj_4507), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1258));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i859_3_lut (.I0(n1258), .I1(n1325), .I2(n1283), .I3(GND_net), 
            .O(n1357));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i25_3_lut (.I0(communication_counter[24]), .I1(n9_adj_4508), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1158));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i791_3_lut (.I0(n1158), .I1(n1225), .I2(n1184), .I3(GND_net), 
            .O(n1257));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i858_3_lut (.I0(n1257), .I1(n1324), .I2(n1283), .I3(GND_net), 
            .O(n1356));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[0]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_106[0]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i723_3_lut (.I0(n1058), .I1(n1125), .I2(n1085), .I3(GND_net), 
            .O(n1157));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i790_3_lut (.I0(n1157), .I1(n1224), .I2(n1184), .I3(GND_net), 
            .O(n1256));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i857_3_lut (.I0(n1256), .I1(n1323), .I2(n1283), .I3(GND_net), 
            .O(n1355));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[1]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_46_i637_3_lut_3_lut (.I0(n938), .I1(n5803), .I2(n917), 
            .I3(GND_net), .O(n1046));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i637_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_70_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_106[1]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i722_3_lut (.I0(n1057), .I1(n1124), .I2(n1085), .I3(GND_net), 
            .O(n1156));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i789_3_lut (.I0(n1156), .I1(n1223), .I2(n1184), .I3(GND_net), 
            .O(n1255));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i856_3_lut (.I0(n1255), .I1(n1322), .I2(n1283), .I3(GND_net), 
            .O(n1354));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[2]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_106[2]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i721_3_lut (.I0(n1056), .I1(n1123), .I2(n1085), .I3(GND_net), 
            .O(n1155));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i788_3_lut (.I0(n1155), .I1(n1222), .I2(n1184), .I3(GND_net), 
            .O(n1254));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i855_3_lut (.I0(n1254), .I1(n1321), .I2(n1283), .I3(GND_net), 
            .O(n1353));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4322), .I3(n15), .O(motor_state_23__N_106[3]));   // verilog/TinyFPGA_B.v(229[5] 232[10])
    defparam mux_71_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_106[3]), 
            .I2(n15_adj_4321), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(228[5] 232[10])
    defparam mux_70_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i720_3_lut (.I0(n1055), .I1(n1122), .I2(n1085), .I3(GND_net), 
            .O(n1154));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i787_3_lut (.I0(n1154), .I1(n1221), .I2(n1184), .I3(GND_net), 
            .O(n1253));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i854_3_lut (.I0(n1253), .I1(n1320), .I2(n1283), .I3(GND_net), 
            .O(n1352));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n6075), 
            .I3(n2724), .O(n41_adj_4915));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n6076), 
            .I3(n2724), .O(n39_adj_4914));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4358), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n670));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n6073), 
            .I3(n2724), .O(n45_adj_4917));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n6074), 
            .I3(n2724), .O(n43_adj_4916));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n6077), 
            .I3(n2724), .O(n37_adj_4913));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i21_4_lut (.I0(n2712_adj_4420), .I1(n90), 
            .I2(n6085), .I3(n2724), .O(n21_adj_4903));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n6084), 
            .I3(n2724), .O(n23_adj_4904));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i25_4_lut (.I0(n2710_adj_4419), .I1(n88), 
            .I2(n6083), .I3(n2724), .O(n25_adj_4906));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i17_4_lut (.I0(n2714_adj_4421), .I1(n92), 
            .I2(n6087), .I3(n2724), .O(n17_adj_4901));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n6086), 
            .I3(n2724), .O(n19_adj_4902));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n6092), 
            .I3(n2724), .O(n7_adj_4892));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i29_4_lut (.I0(n2708_adj_4418), .I1(n86), 
            .I2(n6081), .I3(n2724), .O(n29_adj_4908));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n6080), 
            .I3(n2724), .O(n31_adj_4910));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i9_4_lut (.I0(n2718_adj_4423), .I1(n96), 
            .I2(n6091), .I3(n2724), .O(n9_adj_4894));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4627));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n6078), 
            .I3(n2724), .O(n35_adj_4912));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n6090), 
            .I3(n2724), .O(n11_adj_4896));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i13_4_lut (.I0(n2716_adj_4422), .I1(n94), 
            .I2(n6089), .I3(n2724), .O(n13_adj_4898));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n6082), 
            .I3(n2724), .O(n27_adj_4907));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n6088), 
            .I3(n2724), .O(n15_adj_4899));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n6079), 
            .I3(n2724), .O(n33_adj_4911));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33987_4_lut (.I0(n27_adj_4907), .I1(n15_adj_4899), .I2(n13_adj_4898), 
            .I3(n11_adj_4896), .O(n40751));
    defparam i33987_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4911), 
            .I3(GND_net), .O(n12_adj_4897));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i33965_2_lut (.I0(n33_adj_4911), .I1(n15_adj_4899), .I2(GND_net), 
            .I3(GND_net), .O(n40729));
    defparam i33965_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4898), 
            .I3(GND_net), .O(n10_adj_4895));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i30_3_lut (.I0(n12_adj_4897), .I1(n83), 
            .I2(n35_adj_4912), .I3(GND_net), .O(n30_adj_4909));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1828_3_lut (.I0(n2720_adj_4424), .I1(n6093), .I2(n2724), 
            .I3(GND_net), .O(n2798));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33653_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n40415));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33653_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i34035_3_lut (.I0(n7_adj_4892), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n40799));
    defparam i34035_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i34646_4_lut (.I0(n13_adj_4898), .I1(n11_adj_4896), .I2(n9_adj_4894), 
            .I3(n40799), .O(n41410));
    defparam i34646_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34634_4_lut (.I0(n19_adj_4902), .I1(n17_adj_4901), .I2(n15_adj_4899), 
            .I3(n41410), .O(n41398));
    defparam i34634_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35359_4_lut (.I0(n25_adj_4906), .I1(n23_adj_4904), .I2(n21_adj_4903), 
            .I3(n41398), .O(n42123));
    defparam i35359_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34932_4_lut (.I0(n31_adj_4910), .I1(n29_adj_4908), .I2(n27_adj_4907), 
            .I3(n42123), .O(n41696));
    defparam i34932_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35454_4_lut (.I0(n37_adj_4913), .I1(n35_adj_4912), .I2(n33_adj_4911), 
            .I3(n41696), .O(n42218));
    defparam i35454_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4916), 
            .I3(GND_net), .O(n16_adj_4900));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4892), 
            .I3(GND_net), .O(n6_adj_4891));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i35022_3_lut (.I0(n6_adj_4891), .I1(n90), .I2(n21_adj_4903), 
            .I3(GND_net), .O(n41786));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35022_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35023_3_lut (.I0(n41786), .I1(n89), .I2(n23_adj_4904), .I3(GND_net), 
            .O(n41787));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35023_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34013_4_lut (.I0(n21_adj_4903), .I1(n19_adj_4902), .I2(n17_adj_4901), 
            .I3(n9_adj_4894), .O(n40777));
    defparam i34013_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33927_2_lut (.I0(n43_adj_4916), .I1(n19_adj_4902), .I2(GND_net), 
            .I3(GND_net), .O(n40691));
    defparam i33927_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4901), 
            .I3(GND_net), .O(n8_adj_4893));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_LessThan_1830_i24_3_lut (.I0(n16_adj_4900), .I1(n78), 
            .I2(n45_adj_4917), .I3(GND_net), .O(n24_adj_4905));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33935_4_lut (.I0(n43_adj_4916), .I1(n25_adj_4906), .I2(n23_adj_4904), 
            .I3(n40777), .O(n40699));
    defparam i33935_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35133_4_lut (.I0(n24_adj_4905), .I1(n8_adj_4893), .I2(n45_adj_4917), 
            .I3(n40691), .O(n41897));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35133_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34451_3_lut (.I0(n41787), .I1(n88), .I2(n25_adj_4906), .I3(GND_net), 
            .O(n41215));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34451_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1829_3_lut (.I0(n669), .I1(n6094), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i4_4_lut (.I0(n670), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4890));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35020_3_lut (.I0(n4_adj_4890), .I1(n87), .I2(n27_adj_4907), 
            .I3(GND_net), .O(n41784));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35020_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35021_3_lut (.I0(n41784), .I1(n86), .I2(n29_adj_4908), .I3(GND_net), 
            .O(n41785));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35021_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33973_4_lut (.I0(n33_adj_4911), .I1(n31_adj_4910), .I2(n29_adj_4908), 
            .I3(n40751), .O(n40737));
    defparam i33973_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35363_4_lut (.I0(n30_adj_4909), .I1(n10_adj_4895), .I2(n35_adj_4912), 
            .I3(n40729), .O(n42127));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35363_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34453_3_lut (.I0(n41785), .I1(n85), .I2(n31_adj_4910), .I3(GND_net), 
            .O(n41217));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34453_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35534_4_lut (.I0(n41217), .I1(n42127), .I2(n35_adj_4912), 
            .I3(n40737), .O(n42298));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35534_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35535_3_lut (.I0(n42298), .I1(n82), .I2(n37_adj_4913), .I3(GND_net), 
            .O(n42299));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35535_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35488_3_lut (.I0(n42299), .I1(n81), .I2(n39_adj_4914), .I3(GND_net), 
            .O(n42252));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35488_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33945_4_lut (.I0(n43_adj_4916), .I1(n41_adj_4915), .I2(n39_adj_4914), 
            .I3(n42218), .O(n40709));
    defparam i33945_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35446_4_lut (.I0(n41215), .I1(n41897), .I2(n45_adj_4917), 
            .I3(n40699), .O(n42210));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35446_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34459_3_lut (.I0(n42252), .I1(n80), .I2(n41_adj_4915), .I3(GND_net), 
            .O(n41223));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34459_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1807_3_lut (.I0(n2699), .I1(n6072), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35448_4_lut (.I0(n41223), .I1(n42210), .I2(n45_adj_4917), 
            .I3(n40709), .O(n42212));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35448_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35449_3_lut (.I0(n42212), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35449_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_46_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4887));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4885));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4889));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4888));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i25_2_lut (.I0(n2710_adj_4419), .I1(n89), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4882));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4883));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i21_2_lut (.I0(n2712_adj_4420), .I1(n91), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4880));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4881));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n669));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4879));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i9_2_lut (.I0(n2718_adj_4423), .I1(n97), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4871));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4873));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i13_2_lut (.I0(n2716_adj_4422), .I1(n95), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4875));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4877));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i17_2_lut (.I0(n2714_adj_4421), .I1(n93), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4878));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i29_2_lut (.I0(n2708_adj_4418), .I1(n87), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4884));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34118_4_lut (.I0(n29_adj_4884), .I1(n17_adj_4878), .I2(n15_adj_4877), 
            .I3(n13_adj_4875), .O(n40882));
    defparam i34118_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34197_4_lut (.I0(n11_adj_4873), .I1(n9_adj_4871), .I2(n2719), 
            .I3(n98), .O(n40961));
    defparam i34197_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34758_4_lut (.I0(n17_adj_4878), .I1(n15_adj_4877), .I2(n13_adj_4875), 
            .I3(n40961), .O(n41522));
    defparam i34758_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34752_4_lut (.I0(n23_adj_4881), .I1(n21_adj_4880), .I2(n19_adj_4879), 
            .I3(n41522), .O(n41516));
    defparam i34752_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34127_4_lut (.I0(n29_adj_4884), .I1(n27_adj_4883), .I2(n25_adj_4882), 
            .I3(n41516), .O(n40891));
    defparam i34127_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1777_i6_4_lut (.I0(n669), .I1(n99), .I2(n2720_adj_4424), 
            .I3(n558), .O(n6_adj_4869));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35028_3_lut (.I0(n6_adj_4869), .I1(n87), .I2(n29_adj_4884), 
            .I3(GND_net), .O(n41792));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35028_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1777_i32_3_lut (.I0(n14_adj_4876), .I1(n83), 
            .I2(n37_adj_4889), .I3(GND_net), .O(n32_adj_4886));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35029_3_lut (.I0(n41792), .I1(n86), .I2(n31_adj_4885), .I3(GND_net), 
            .O(n41793));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35029_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34097_4_lut (.I0(n35_adj_4888), .I1(n33_adj_4887), .I2(n31_adj_4885), 
            .I3(n40882), .O(n40861));
    defparam i34097_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35347_4_lut (.I0(n32_adj_4886), .I1(n12_adj_4874), .I2(n37_adj_4889), 
            .I3(n40854), .O(n42111));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35347_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34439_3_lut (.I0(n41793), .I1(n85), .I2(n33_adj_4887), .I3(GND_net), 
            .O(n41203));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34439_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35030_3_lut (.I0(n8_adj_4870), .I1(n90), .I2(n23_adj_4881), 
            .I3(GND_net), .O(n41794));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35030_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35031_3_lut (.I0(n41794), .I1(n89), .I2(n25_adj_4882), .I3(GND_net), 
            .O(n41795));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35031_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34744_4_lut (.I0(n25_adj_4882), .I1(n23_adj_4881), .I2(n21_adj_4880), 
            .I3(n40227), .O(n41508));
    defparam i34744_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35131_3_lut (.I0(n10_adj_4872), .I1(n91), .I2(n21_adj_4880), 
            .I3(GND_net), .O(n41895));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35131_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34437_3_lut (.I0(n41795), .I1(n88), .I2(n27_adj_4883), .I3(GND_net), 
            .O(n41201));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34437_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35199_4_lut (.I0(n35_adj_4888), .I1(n33_adj_4887), .I2(n31_adj_4885), 
            .I3(n40891), .O(n41963));
    defparam i35199_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35532_4_lut (.I0(n41203), .I1(n42111), .I2(n37_adj_4889), 
            .I3(n40861), .O(n42296));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35532_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35225_4_lut (.I0(n41201), .I1(n41895), .I2(n27_adj_4883), 
            .I3(n41508), .O(n41989));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35225_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35569_4_lut (.I0(n41989), .I1(n42296), .I2(n37_adj_4889), 
            .I3(n41963), .O(n42333));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35569_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35570_3_lut (.I0(n42333), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n42334));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35570_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35468_3_lut (.I0(n42334), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n42232));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35468_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35419_3_lut (.I0(n42232), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n42183));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35419_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35420_3_lut (.I0(n42183), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n42184));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35420_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1992_4_lut (.I0(n42184), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1992_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 i8_4_lut_adj_1784 (.I0(n1846), .I1(n1844), .I2(n1850), .I3(n1852), 
            .O(n19_adj_4351));
    defparam i8_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1722_i45_2_lut (.I0(n2619), .I1(n80), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4868));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i41_2_lut (.I0(n2621), .I1(n82), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4865));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i43_2_lut (.I0(n2620), .I1(n81), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4866));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4393), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n668));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4860));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4862));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i724_3_lut_3_lut (.I0(n1067), .I1(n5813), .I2(n1048), 
            .I3(GND_net), .O(n1174));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i724_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4857));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4858));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4855));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4856));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4864));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4845));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i725_3_lut_3_lut (.I0(n1067), .I1(n5814), .I2(n653), 
            .I3(GND_net), .O(n1175));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i725_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4656));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4849));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4851));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4852));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4859));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33535_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n40297));
    defparam i33535_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4863));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4658));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4847));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4854));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4667));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33513_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n40275));
    defparam i33513_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4669));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut (.I0(n855), .I1(n884), .I2(n956), .I3(n958), 
            .O(n35536));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfff6;
    SB_LUT4 i33511_4_lut (.I0(n31_adj_4859), .I1(n19_adj_4852), .I2(n17_adj_4851), 
            .I3(n15_adj_4849), .O(n40273));
    defparam i33511_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1722_i34_3_lut (.I0(n16_adj_4850), .I1(n83), 
            .I2(n39_adj_4864), .I3(GND_net), .O(n34_adj_4861));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34253_4_lut (.I0(n13_adj_4847), .I1(n11_adj_4845), .I2(n2637), 
            .I3(n98), .O(n41017));
    defparam i34253_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34782_4_lut (.I0(n19_adj_4852), .I1(n17_adj_4851), .I2(n15_adj_4849), 
            .I3(n41017), .O(n41546));
    defparam i34782_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34778_4_lut (.I0(n25_adj_4856), .I1(n23_adj_4855), .I2(n21_adj_4854), 
            .I3(n41546), .O(n41542));
    defparam i34778_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33515_4_lut (.I0(n31_adj_4859), .I1(n29_adj_4858), .I2(n27_adj_4857), 
            .I3(n41542), .O(n40277));
    defparam i33515_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35008_4_lut (.I0(n37_adj_4863), .I1(n35_adj_4862), .I2(n33_adj_4860), 
            .I3(n40277), .O(n41772));
    defparam i35008_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35241_3_lut (.I0(n10_adj_4844), .I1(n90), .I2(n25_adj_4856), 
            .I3(GND_net), .O(n42005));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35241_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35242_3_lut (.I0(n42005), .I1(n89), .I2(n27_adj_4857), .I3(GND_net), 
            .O(n42006));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35242_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i887_3_lut_3_lut (.I0(n1316), .I1(n5831), .I2(n1296), 
            .I3(GND_net), .O(n1416));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i887_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34235_4_lut (.I0(n27_adj_4857), .I1(n25_adj_4856), .I2(n23_adj_4855), 
            .I3(n40293), .O(n40999));
    defparam i34235_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1722_i20_3_lut (.I0(n12_adj_4846), .I1(n91), 
            .I2(n23_adj_4855), .I3(GND_net), .O(n20_adj_4853));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35122_3_lut (.I0(n42006), .I1(n88), .I2(n29_adj_4858), .I3(GND_net), 
            .O(n41886));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35122_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1722_i8_4_lut (.I0(n668), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4843));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35239_3_lut (.I0(n8_adj_4843), .I1(n87), .I2(n31_adj_4859), 
            .I3(GND_net), .O(n42003));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35239_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35240_3_lut (.I0(n42003), .I1(n86), .I2(n33_adj_4860), .I3(GND_net), 
            .O(n42004));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35240_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33499_4_lut (.I0(n37_adj_4863), .I1(n35_adj_4862), .I2(n33_adj_4860), 
            .I3(n40273), .O(n40261));
    defparam i33499_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35479_4_lut (.I0(n34_adj_4861), .I1(n14_adj_4848), .I2(n39_adj_4864), 
            .I3(n40255), .O(n42243));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35479_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35124_3_lut (.I0(n42004), .I1(n85), .I2(n35_adj_4862), .I3(GND_net), 
            .O(n41888));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35124_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35555_4_lut (.I0(n41888), .I1(n42243), .I2(n39_adj_4864), 
            .I3(n40261), .O(n42319));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35555_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35556_3_lut (.I0(n42319), .I1(n82), .I2(n41_adj_4865), .I3(GND_net), 
            .O(n42320));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35556_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35523_3_lut (.I0(n42320), .I1(n81), .I2(n43_adj_4866), .I3(GND_net), 
            .O(n42287));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35523_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i994_3_lut (.I0(n1457), .I1(n1524), .I2(n1481), .I3(GND_net), 
            .O(n1556));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35481_4_lut (.I0(n43_adj_4866), .I1(n41_adj_4865), .I2(n39_adj_4864), 
            .I3(n41772), .O(n42245));
    defparam i35481_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i722_3_lut_3_lut (.I0(n1067), .I1(n5811), .I2(n1046), 
            .I3(GND_net), .O(n1172));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i722_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35127_4_lut (.I0(n41886), .I1(n20_adj_4853), .I2(n29_adj_4858), 
            .I3(n40999), .O(n41891));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35127_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_46_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4679));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35505_3_lut (.I0(n42287), .I1(n80), .I2(n45_adj_4868), .I3(GND_net), 
            .O(n44_adj_4867));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35505_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35129_4_lut (.I0(n44_adj_4867), .I1(n41891), .I2(n45_adj_4868), 
            .I3(n42245), .O(n41893));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35129_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n41893), .I1(n15549), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'hceef;
    SB_LUT4 i33477_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n40239));
    defparam i33477_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4681));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34144_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n40908));
    defparam i34144_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4696));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4692));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34129_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n40893));
    defparam i34129_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4840));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4694));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4842));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4838));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4706));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4357), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n667));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34081_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n40845));
    defparam i34081_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4841));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4708));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34093_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n40857));
    defparam i34093_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4835));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4836));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4710));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i721_3_lut_3_lut (.I0(n1067), .I1(n5810), .I2(n1045), 
            .I3(GND_net), .O(n1171));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i721_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4723));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4823));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4825));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34025_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n40789));
    defparam i34025_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4725));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34037_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n40801));
    defparam i34037_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4832));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4833));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4834));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4727));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4740));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4827));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4829));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33975_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n40739));
    defparam i33975_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4830));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4837));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33570_4_lut (.I0(n33_adj_4837), .I1(n21_adj_4830), .I2(n19_adj_4829), 
            .I3(n17_adj_4827), .O(n40332));
    defparam i33570_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34309_4_lut (.I0(n15_adj_4825), .I1(n13_adj_4823), .I2(n2552), 
            .I3(n98), .O(n41073));
    defparam i34309_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 div_46_i720_3_lut_3_lut (.I0(n1067), .I1(n5809), .I2(n1044), 
            .I3(GND_net), .O(n1170));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i720_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34806_4_lut (.I0(n21_adj_4830), .I1(n19_adj_4829), .I2(n17_adj_4827), 
            .I3(n41073), .O(n41570));
    defparam i34806_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34802_4_lut (.I0(n27_adj_4834), .I1(n25_adj_4833), .I2(n23_adj_4832), 
            .I3(n41570), .O(n41566));
    defparam i34802_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33577_4_lut (.I0(n33_adj_4837), .I1(n31_adj_4836), .I2(n29_adj_4835), 
            .I3(n41566), .O(n40339));
    defparam i33577_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_i886_3_lut_3_lut (.I0(n1316), .I1(n5830), .I2(n1295), 
            .I3(GND_net), .O(n1415));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i886_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1665_i10_4_lut (.I0(n667), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4821));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35247_3_lut (.I0(n10_adj_4821), .I1(n87), .I2(n33_adj_4837), 
            .I3(GND_net), .O(n42011));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35247_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4742));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35248_3_lut (.I0(n42011), .I1(n86), .I2(n35_adj_4838), .I3(GND_net), 
            .O(n42012));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35248_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i36_3_lut (.I0(n18_adj_4828), .I1(n83), 
            .I2(n41_adj_4842), .I3(GND_net), .O(n36_adj_4839));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33560_4_lut (.I0(n39_adj_4841), .I1(n37_adj_4840), .I2(n35_adj_4838), 
            .I3(n40332), .O(n40322));
    defparam i33560_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35477_4_lut (.I0(n36_adj_4839), .I1(n16_adj_4826), .I2(n41_adj_4842), 
            .I3(n40318), .O(n42241));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35477_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35118_3_lut (.I0(n42012), .I1(n85), .I2(n37_adj_4840), .I3(GND_net), 
            .O(n41882));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35118_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i22_3_lut (.I0(n14_adj_4824), .I1(n91), 
            .I2(n25_adj_4833), .I3(GND_net), .O(n22_adj_4831));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35475_4_lut (.I0(n22_adj_4831), .I1(n12_adj_4822), .I2(n25_adj_4833), 
            .I3(n40361), .O(n42239));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35475_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35476_3_lut (.I0(n42239), .I1(n90), .I2(n27_adj_4834), .I3(GND_net), 
            .O(n42240));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35476_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35394_3_lut (.I0(n42240), .I1(n89), .I2(n29_adj_4835), .I3(GND_net), 
            .O(n42158));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35394_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i1061_3_lut (.I0(n1556), .I1(n1623), .I2(n1580), .I3(GND_net), 
            .O(n1655));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35016_4_lut (.I0(n39_adj_4841), .I1(n37_adj_4840), .I2(n35_adj_4838), 
            .I3(n40339), .O(n41780));
    defparam i35016_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35553_4_lut (.I0(n41882), .I1(n42241), .I2(n41_adj_4842), 
            .I3(n40322), .O(n42317));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35553_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35318_3_lut (.I0(n42158), .I1(n88), .I2(n31_adj_4836), .I3(GND_net), 
            .O(n42082));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35318_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4744));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35573_4_lut (.I0(n42082), .I1(n42317), .I2(n41_adj_4842), 
            .I3(n41780), .O(n42337));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35573_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35574_3_lut (.I0(n42337), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n42338));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35574_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35572_3_lut (.I0(n42338), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n42336));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35572_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n42336), .I1(n15546), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hceef;
    SB_LUT4 i33991_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n40755));
    defparam i33991_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4760));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33923_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n40687));
    defparam i33923_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4818));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4762));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4816));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4764));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4820));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33937_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n40701));
    defparam i33937_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4819));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4778));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33806_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n40570));
    defparam i33806_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4780));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4782));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4810));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4811));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4812));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33717_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n40479));
    defparam i33717_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4392), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n666));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4784));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4801));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4800));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4803));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33694_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n40456));
    defparam i33694_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4802));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4804));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4813));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4814));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33634_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n40396));
    defparam i33634_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4806));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i719_3_lut_3_lut (.I0(n1067), .I1(n5808), .I2(n1043), 
            .I3(GND_net), .O(n1169_adj_4409));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4805));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4807));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4808));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4815));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33649_4_lut (.I0(n35_adj_4815), .I1(n23_adj_4808), .I2(n21_adj_4807), 
            .I3(n19_adj_4805), .O(n40411));
    defparam i33649_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34388_4_lut (.I0(n17_adj_4803), .I1(n15_adj_4801), .I2(n2464), 
            .I3(n98), .O(n41152));
    defparam i34388_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34820_4_lut (.I0(n23_adj_4808), .I1(n21_adj_4807), .I2(n19_adj_4805), 
            .I3(n41152), .O(n41584));
    defparam i34820_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34816_4_lut (.I0(n29_adj_4812), .I1(n27_adj_4811), .I2(n25_adj_4810), 
            .I3(n41584), .O(n41580));
    defparam i34816_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33651_4_lut (.I0(n35_adj_4815), .I1(n33_adj_4814), .I2(n31_adj_4813), 
            .I3(n41580), .O(n40413));
    defparam i33651_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1606_i12_4_lut (.I0(n666), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_4799));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35253_3_lut (.I0(n12_adj_4799), .I1(n87), .I2(n35_adj_4815), 
            .I3(GND_net), .O(n42017));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35253_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4822));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i38_3_lut (.I0(n20_adj_4806), .I1(n83), 
            .I2(n43_adj_4820), .I3(GND_net), .O(n38_adj_4817));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35254_3_lut (.I0(n42017), .I1(n86), .I2(n37_adj_4816), .I3(GND_net), 
            .O(n42018));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35254_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33638_4_lut (.I0(n41_adj_4819), .I1(n39_adj_4818), .I2(n37_adj_4816), 
            .I3(n40411), .O(n40400));
    defparam i33638_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35251_4_lut (.I0(n38_adj_4817), .I1(n18_adj_4804), .I2(n43_adj_4820), 
            .I3(n40396), .O(n42015));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35251_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33599_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n40361));
    defparam i33599_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i35112_3_lut (.I0(n42018), .I1(n85), .I2(n39_adj_4818), .I3(GND_net), 
            .O(n41876));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35112_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4824));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i24_3_lut (.I0(n16_adj_4802), .I1(n91), 
            .I2(n27_adj_4811), .I3(GND_net), .O(n24_adj_4809));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35473_4_lut (.I0(n24_adj_4809), .I1(n14_adj_4800), .I2(n27_adj_4811), 
            .I3(n40456), .O(n42237));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35473_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35474_3_lut (.I0(n42237), .I1(n90), .I2(n29_adj_4812), .I3(GND_net), 
            .O(n42238));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35474_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35396_3_lut (.I0(n42238), .I1(n89), .I2(n31_adj_4813), .I3(GND_net), 
            .O(n42160));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35396_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35046_4_lut (.I0(n41_adj_4819), .I1(n39_adj_4818), .I2(n37_adj_4816), 
            .I3(n40413), .O(n41810));
    defparam i35046_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35458_4_lut (.I0(n41876), .I1(n42015), .I2(n43_adj_4820), 
            .I3(n40400), .O(n42222));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35458_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35316_3_lut (.I0(n42160), .I1(n88), .I2(n33_adj_4814), .I3(GND_net), 
            .O(n42080));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35316_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35561_4_lut (.I0(n42080), .I1(n42222), .I2(n43_adj_4820), 
            .I3(n41810), .O(n42325));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35561_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_46_i723_3_lut_3_lut (.I0(n1067), .I1(n5812), .I2(n1047), 
            .I3(GND_net), .O(n1173));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i723_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35562_3_lut (.I0(n42325), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n42326));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35562_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n42326), .I1(n15543), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4826));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33556_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n40318));
    defparam i33556_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4828));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4796));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4798));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4794));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4632));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n665));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4846));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4788));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4789));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4790));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4844));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i1128_3_lut (.I0(n1655), .I1(n1722), .I2(n1679), .I3(GND_net), 
            .O(n1754_adj_4494));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4797));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4848));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33493_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n40255));
    defparam i33493_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4850));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4779));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4781));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33531_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n40293));
    defparam i33531_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4783));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4785));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4786));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718_adj_4423), 
            .I3(GND_net), .O(n8_adj_4870));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4874));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4791));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4792));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4793));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33743_4_lut (.I0(n37_adj_4793), .I1(n25_adj_4786), .I2(n23_adj_4785), 
            .I3(n21_adj_4783), .O(n40505));
    defparam i33743_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34502_4_lut (.I0(n19_adj_4781), .I1(n17_adj_4779), .I2(n2373), 
            .I3(n98), .O(n41266));
    defparam i34502_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i34876_4_lut (.I0(n25_adj_4786), .I1(n23_adj_4785), .I2(n21_adj_4783), 
            .I3(n41266), .O(n41640));
    defparam i34876_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34870_4_lut (.I0(n31_adj_4790), .I1(n29_adj_4789), .I2(n27_adj_4788), 
            .I3(n41640), .O(n41634));
    defparam i34870_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33745_4_lut (.I0(n37_adj_4793), .I1(n35_adj_4792), .I2(n33_adj_4791), 
            .I3(n41634), .O(n40507));
    defparam i33745_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1545_i14_4_lut (.I0(n665), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4777));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35257_3_lut (.I0(n14_adj_4777), .I1(n87), .I2(n37_adj_4793), 
            .I3(GND_net), .O(n42021));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35257_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35258_3_lut (.I0(n42021), .I1(n86), .I2(n39_adj_4794), .I3(GND_net), 
            .O(n42022));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35258_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1545_i40_3_lut (.I0(n22_adj_4784), .I1(n83), 
            .I2(n45_adj_4798), .I3(GND_net), .O(n40_adj_4795));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33725_4_lut (.I0(n43_adj_4797), .I1(n41_adj_4796), .I2(n39_adj_4794), 
            .I3(n40505), .O(n40487));
    defparam i33725_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34856_4_lut (.I0(n40_adj_4795), .I1(n20_adj_4782), .I2(n45_adj_4798), 
            .I3(n40479), .O(n41620));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34856_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35108_3_lut (.I0(n42022), .I1(n85), .I2(n41_adj_4796), .I3(GND_net), 
            .O(n41872));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35108_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1545_i26_3_lut (.I0(n18_adj_4780), .I1(n91), 
            .I2(n29_adj_4789), .I3(GND_net), .O(n26_adj_4787));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33640_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n40402));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33640_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i34090_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714_adj_4421), 
            .I3(n93), .O(n40854));
    defparam i34090_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i35339_4_lut (.I0(n26_adj_4787), .I1(n16_adj_4778), .I2(n29_adj_4789), 
            .I3(n40570), .O(n42103));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35339_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35340_3_lut (.I0(n42103), .I1(n90), .I2(n31_adj_4790), .I3(GND_net), 
            .O(n42104));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35340_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35232_3_lut (.I0(n42104), .I1(n89), .I2(n33_adj_4791), .I3(GND_net), 
            .O(n41996));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35232_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35098_4_lut (.I0(n43_adj_4797), .I1(n41_adj_4796), .I2(n39_adj_4794), 
            .I3(n40507), .O(n41862));
    defparam i35098_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35312_4_lut (.I0(n41872), .I1(n41620), .I2(n45_adj_4798), 
            .I3(n40487), .O(n42076));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35312_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34435_3_lut (.I0(n41996), .I1(n88), .I2(n35_adj_4792), .I3(GND_net), 
            .O(n41199));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34435_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35314_4_lut (.I0(n41199), .I1(n42076), .I2(n45_adj_4798), 
            .I3(n41862), .O(n42078));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35314_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n42078), .I1(n15535), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4876));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4872));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33465_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n40227));
    defparam i33465_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4773));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4776));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4775));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4774));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n664));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4770));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4771));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4772));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4761));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4763));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4765));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4766));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4767));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4769));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4759));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33939_4_lut (.I0(n23_adj_4765), .I1(n21_adj_4763), .I2(n19_adj_4761), 
            .I3(n17_adj_4759), .O(n40703));
    defparam i33939_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33929_4_lut (.I0(n29_adj_4769), .I1(n27_adj_4767), .I2(n25_adj_4766), 
            .I3(n40703), .O(n40693));
    defparam i33929_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35171_4_lut (.I0(n35_adj_4772), .I1(n33_adj_4771), .I2(n31_adj_4770), 
            .I3(n40693), .O(n41935));
    defparam i35171_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1482_i16_4_lut (.I0(n664), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4758));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35034_3_lut (.I0(n16_adj_4758), .I1(n87), .I2(n39_adj_4774), 
            .I3(GND_net), .O(n41798));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35034_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35035_3_lut (.I0(n41798), .I1(n86), .I2(n41_adj_4775), .I3(GND_net), 
            .O(n41799));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35035_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34526_4_lut (.I0(n41_adj_4775), .I1(n39_adj_4774), .I2(n27_adj_4767), 
            .I3(n40701), .O(n41290));
    defparam i34526_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35105_3_lut (.I0(n22_adj_4764), .I1(n93), .I2(n27_adj_4767), 
            .I3(GND_net), .O(n41869));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35105_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34427_3_lut (.I0(n41799), .I1(n85), .I2(n43_adj_4776), .I3(GND_net), 
            .O(n41191));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34427_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i888_3_lut_3_lut (.I0(n1316), .I1(n5832), .I2(n1297), 
            .I3(GND_net), .O(n1417));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i888_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1482_i28_3_lut (.I0(n20_adj_4762), .I1(n91), 
            .I2(n31_adj_4770), .I3(GND_net), .O(n28_adj_4768));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i885_3_lut_3_lut (.I0(n1316), .I1(n5829), .I2(n1294), 
            .I3(GND_net), .O(n1414));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i885_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35417_4_lut (.I0(n28_adj_4768), .I1(n18_adj_4760), .I2(n31_adj_4770), 
            .I3(n40687), .O(n42181));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35417_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35418_3_lut (.I0(n42181), .I1(n90), .I2(n33_adj_4771), .I3(GND_net), 
            .O(n42182));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35418_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35244_3_lut (.I0(n42182), .I1(n89), .I2(n35_adj_4772), .I3(GND_net), 
            .O(n42008));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35244_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34528_4_lut (.I0(n41_adj_4775), .I1(n39_adj_4774), .I2(n37_adj_4773), 
            .I3(n41935), .O(n41292));
    defparam i34528_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35235_4_lut (.I0(n41191), .I1(n41869), .I2(n43_adj_4776), 
            .I3(n41290), .O(n41999));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35235_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34425_3_lut (.I0(n42008), .I1(n88), .I2(n37_adj_4773), .I3(GND_net), 
            .O(n41189));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34425_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35491_4_lut (.I0(n41189), .I1(n41999), .I2(n43_adj_4776), 
            .I3(n41292), .O(n42255));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35491_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35492_3_lut (.I0(n42255), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n42256));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35492_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n42256), .I1(n15530), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4754));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4757));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4756));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_mux_3_i31_3_lut (.I0(communication_counter[30]), .I1(n3_adj_4514), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n852));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4755));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4748));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4750));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n663));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4751));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4752));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4753));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4747));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4741));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4743));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4745));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4739));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33999_4_lut (.I0(n25_adj_4745), .I1(n23_adj_4743), .I2(n21_adj_4741), 
            .I3(n19_adj_4739), .O(n40763));
    defparam i33999_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33983_4_lut (.I0(n31_adj_4750), .I1(n29_adj_4748), .I2(n27_adj_4747), 
            .I3(n40763), .O(n40747));
    defparam i33983_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35181_4_lut (.I0(n37_adj_4753), .I1(n35_adj_4752), .I2(n33_adj_4751), 
            .I3(n40747), .O(n41945));
    defparam i35181_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1417_i18_4_lut (.I0(n663), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4738));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35038_3_lut (.I0(n18_adj_4738), .I1(n87), .I2(n41_adj_4755), 
            .I3(GND_net), .O(n41802));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35038_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35039_3_lut (.I0(n41802), .I1(n86), .I2(n43_adj_4756), .I3(GND_net), 
            .O(n41803));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35039_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34572_4_lut (.I0(n43_adj_4756), .I1(n41_adj_4755), .I2(n29_adj_4748), 
            .I3(n40755), .O(n41336));
    defparam i34572_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1417_i26_3_lut (.I0(n24_adj_4744), .I1(n93), 
            .I2(n29_adj_4748), .I3(GND_net), .O(n26_adj_4746));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34421_3_lut (.I0(n41803), .I1(n85), .I2(n45_adj_4757), .I3(GND_net), 
            .O(n41185));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34421_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1417_i30_3_lut (.I0(n22_adj_4742), .I1(n91), 
            .I2(n33_adj_4751), .I3(GND_net), .O(n30_adj_4749));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35415_4_lut (.I0(n30_adj_4749), .I1(n20_adj_4740), .I2(n33_adj_4751), 
            .I3(n40739), .O(n42179));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35415_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35416_3_lut (.I0(n42179), .I1(n90), .I2(n35_adj_4752), .I3(GND_net), 
            .O(n42180));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35416_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35261_3_lut (.I0(n42180), .I1(n89), .I2(n37_adj_4753), .I3(GND_net), 
            .O(n42025));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35261_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34578_4_lut (.I0(n43_adj_4756), .I1(n41_adj_4755), .I2(n39_adj_4754), 
            .I3(n41945), .O(n41342));
    defparam i34578_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35102_4_lut (.I0(n41185), .I1(n26_adj_4746), .I2(n45_adj_4757), 
            .I3(n41336), .O(n41866));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35102_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34419_3_lut (.I0(n42025), .I1(n88), .I2(n39_adj_4754), .I3(GND_net), 
            .O(n41183));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34419_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35104_4_lut (.I0(n41183), .I1(n41866), .I2(n45_adj_4757), 
            .I3(n41342), .O(n41868));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35104_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n41868), .I1(n15576), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4737));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4736));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4735));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4734));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n662));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4730));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4731));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4733));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12884_3_lut_4_lut (.I0(r_SM_Main_adj_5053[2]), .I1(r_SM_Main_adj_5053[0]), 
            .I2(n26612), .I3(r_SM_Main_adj_5053[1]), .O(n17566));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12884_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 div_46_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4724));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4726));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4728));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4722));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34043_4_lut (.I0(n27_adj_4728), .I1(n25_adj_4726), .I2(n23_adj_4724), 
            .I3(n21_adj_4722), .O(n40807));
    defparam i34043_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34029_4_lut (.I0(n33_adj_4733), .I1(n31_adj_4731), .I2(n29_adj_4730), 
            .I3(n40807), .O(n40793));
    defparam i34029_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1350_i20_4_lut (.I0(n662), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4721));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1350_i28_3_lut (.I0(n26_adj_4727), .I1(n93), 
            .I2(n31_adj_4731), .I3(GND_net), .O(n28_adj_4729));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1350_i32_3_lut (.I0(n24_adj_4725), .I1(n91), 
            .I2(n35_adj_4734), .I3(GND_net), .O(n32_adj_4732));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35409_4_lut (.I0(n32_adj_4732), .I1(n22_adj_4723), .I2(n35_adj_4734), 
            .I3(n40789), .O(n42173));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35409_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35410_3_lut (.I0(n42173), .I1(n90), .I2(n37_adj_4735), .I3(GND_net), 
            .O(n42174));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35410_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35283_3_lut (.I0(n42174), .I1(n89), .I2(n39_adj_4736), .I3(GND_net), 
            .O(n42047));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35283_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35189_4_lut (.I0(n39_adj_4736), .I1(n37_adj_4735), .I2(n35_adj_4734), 
            .I3(n40793), .O(n41953));
    defparam i35189_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35411_4_lut (.I0(n28_adj_4729), .I1(n20_adj_4721), .I2(n31_adj_4731), 
            .I3(n40801), .O(n42175));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35411_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34409_3_lut (.I0(n42047), .I1(n88), .I2(n41_adj_4737), .I3(GND_net), 
            .O(n41173));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34409_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35464_4_lut (.I0(n41173), .I1(n42175), .I2(n41_adj_4737), 
            .I3(n41953), .O(n42228));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35464_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35465_3_lut (.I0(n42228), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n42229));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35465_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35424_3_lut (.I0(n42229), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n42188));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35424_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n42188), .I1(n15573), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4720));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4719));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4718));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4717));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4378), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n661));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4713));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4714));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4716));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4707));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4709));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4711));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4705));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34095_4_lut (.I0(n29_adj_4711), .I1(n27_adj_4709), .I2(n25_adj_4707), 
            .I3(n23_adj_4705), .O(n40859));
    defparam i34095_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34085_4_lut (.I0(n35_adj_4716), .I1(n33_adj_4714), .I2(n31_adj_4713), 
            .I3(n40859), .O(n40849));
    defparam i34085_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1281_i22_4_lut (.I0(n661), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4704));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1281_i30_3_lut (.I0(n28_adj_4710), .I1(n93), 
            .I2(n33_adj_4714), .I3(GND_net), .O(n30_adj_4712));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1281_i34_3_lut (.I0(n26_adj_4708), .I1(n91), 
            .I2(n37_adj_4717), .I3(GND_net), .O(n34_adj_4715));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35407_4_lut (.I0(n34_adj_4715), .I1(n24_adj_4706), .I2(n37_adj_4717), 
            .I3(n40845), .O(n42171));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35407_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35408_3_lut (.I0(n42171), .I1(n90), .I2(n39_adj_4718), .I3(GND_net), 
            .O(n42172));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35408_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35285_3_lut (.I0(n42172), .I1(n89), .I2(n41_adj_4719), .I3(GND_net), 
            .O(n42049));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35285_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35197_4_lut (.I0(n41_adj_4719), .I1(n39_adj_4718), .I2(n37_adj_4717), 
            .I3(n40849), .O(n41961));
    defparam i35197_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35397_4_lut (.I0(n30_adj_4712), .I1(n22_adj_4704), .I2(n33_adj_4714), 
            .I3(n40857), .O(n42161));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35397_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34405_3_lut (.I0(n42049), .I1(n88), .I2(n43_adj_4720), .I3(GND_net), 
            .O(n41169));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34405_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35483_4_lut (.I0(n41169), .I1(n42161), .I2(n43_adj_4720), 
            .I3(n41961), .O(n42247));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35483_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35484_3_lut (.I0(n42247), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n42248));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35484_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n42248), .I1(n15526), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4700));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4320), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n660));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i808_3_lut_3_lut (.I0(n1193), .I1(n5823), .I2(n1175), 
            .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i808_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4699));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4703));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4702));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4693));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4695));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4697));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4691));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34151_4_lut (.I0(n31_adj_4697), .I1(n29_adj_4695), .I2(n27_adj_4693), 
            .I3(n25_adj_4691), .O(n40915));
    defparam i34151_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1210_i36_3_lut (.I0(n28_adj_4694), .I1(n91), 
            .I2(n39_adj_4703), .I3(GND_net), .O(n36_adj_4701));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1210_i24_4_lut (.I0(n660), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4690));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1210_i32_3_lut (.I0(n30_adj_4696), .I1(n93), 
            .I2(n35_adj_4700), .I3(GND_net), .O(n32_adj_4698));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34133_4_lut (.I0(n37_adj_4702), .I1(n35_adj_4700), .I2(n33_adj_4699), 
            .I3(n40915), .O(n40897));
    defparam i34133_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35405_4_lut (.I0(n36_adj_4701), .I1(n26_adj_4692), .I2(n39_adj_4703), 
            .I3(n40893), .O(n42169));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35405_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35092_4_lut (.I0(n32_adj_4698), .I1(n24_adj_4690), .I2(n35_adj_4700), 
            .I3(n40908), .O(n41856));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35092_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35530_4_lut (.I0(n41856), .I1(n42169), .I2(n39_adj_4703), 
            .I3(n40897), .O(n42294));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35530_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35531_3_lut (.I0(n42294), .I1(n90), .I2(n1865), .I3(GND_net), 
            .O(n42295));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35531_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35494_3_lut (.I0(n42295), .I1(n89), .I2(n1864), .I3(GND_net), 
            .O(n42258));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35494_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35094_3_lut (.I0(n42258), .I1(n88), .I2(n1863), .I3(GND_net), 
            .O(n41858));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35094_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n41858), .I1(n15570), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hceef;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n17519(n17519), .encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .n17520(n17520), .n17521(n17521), .n17522(n17522), 
            .n17523(n17523), .n17524(n17524), .n17515(n17515), .n17516(n17516), 
            .n17517(n17517), .n17518(n17518), .n17513(n17513), .n17514(n17514), 
            .n17511(n17511), .n17512(n17512), .n17509(n17509), .n17510(n17510), 
            .n17507(n17507), .n17508(n17508), .n17505(n17505), .n17506(n17506), 
            .n17502(n17502), .n17503(n17503), .n17504(n17504), .data_o({quadA_debounced, 
            quadB_debounced}), .n2940({n2941, n2942, n2943, n2944, 
            n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
            n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, 
            n2961, n2962, n2963, n2964}), .GND_net(GND_net), .count_enable(count_enable), 
            .n16968(n16968), .n17551(n17551), .reg_B({reg_B}), .n37155(n37155), 
            .PIN_2_c_0(PIN_2_c_0), .PIN_1_c_1(PIN_1_c_1), .n16971(n16971)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(254[15] 259[4])
    SB_LUT4 div_46_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4685));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i36257_1_lut_2_lut (.I0(n3362), .I1(n10082), .I2(GND_net), 
            .I3(GND_net), .O(n43021));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i36257_1_lut_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_46_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4684));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i809_3_lut_3_lut (.I0(n1193), .I1(n5824), .I2(n654), 
            .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i809_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4377), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n659));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4688));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4680));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4682));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4683));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4687));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4678));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33497_4_lut (.I0(n33_adj_4683), .I1(n31_adj_4682), .I2(n29_adj_4680), 
            .I3(n27_adj_4678), .O(n40259));
    defparam i33497_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1137_i38_3_lut (.I0(n30_adj_4681), .I1(n91), 
            .I2(n41_adj_4688), .I3(GND_net), .O(n38_adj_4686));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1137_i26_4_lut (.I0(n659), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26_adj_4677));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35304_3_lut (.I0(n26_adj_4677), .I1(n95), .I2(n33_adj_4683), 
            .I3(GND_net), .O(n42068));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35304_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10_4_lut_adj_1794 (.I0(n19_adj_4351), .I1(n1845), .I2(n18_adj_4352), 
            .I3(n12_adj_4353), .O(n1877));
    defparam i10_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1196_3_lut (.I0(n1755_adj_4495), .I1(n1822), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35305_3_lut (.I0(n42068), .I1(n94), .I2(n35_adj_4684), .I3(GND_net), 
            .O(n42069));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35305_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33483_4_lut (.I0(n39_adj_4687), .I1(n37_adj_4685), .I2(n35_adj_4684), 
            .I3(n40259), .O(n40245));
    defparam i33483_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_i805_3_lut_3_lut (.I0(n1193), .I1(n5820), .I2(n1172), 
            .I3(GND_net), .O(n1295));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i805_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35471_4_lut (.I0(n38_adj_4686), .I1(n28_adj_4679), .I2(n41_adj_4688), 
            .I3(n40239), .O(n42235));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35471_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35089_3_lut (.I0(n42069), .I1(n93), .I2(n37_adj_4685), .I3(GND_net), 
            .O(n41853));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35089_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35567_4_lut (.I0(n41853), .I1(n42235), .I2(n41_adj_4688), 
            .I3(n40245), .O(n42331));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35567_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35568_3_lut (.I0(n42331), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n42332));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35568_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35548_3_lut (.I0(n42332), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n42312));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35548_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n42312), .I1(n15522), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4673));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4672));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n658));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4676));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n15491), 
            .O(n249));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 div_46_i804_3_lut_3_lut (.I0(n1193), .I1(n5819), .I2(n1171), 
            .I3(GND_net), .O(n1294));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i804_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut (.I0(n98), .I1(n97), .I2(n96), .I3(n15498), 
            .O(n15491));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4668));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4671));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1796 (.I0(n97), .I1(n96), .I2(n15498), 
            .I3(GND_net), .O(n15555));
    defparam i1_2_lut_3_lut_adj_1796.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4670));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1797 (.I0(n95), .I1(n94), .I2(n93), .I3(n15504), 
            .O(n15498));
    defparam i1_2_lut_4_lut_adj_1797.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4675));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1798 (.I0(n94), .I1(n93), .I2(n15504), 
            .I3(GND_net), .O(n15501));
    defparam i1_2_lut_3_lut_adj_1798.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4666));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33523_4_lut (.I0(n35_adj_4671), .I1(n33_adj_4670), .I2(n31_adj_4668), 
            .I3(n29_adj_4666), .O(n40285));
    defparam i33523_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_i884_3_lut_3_lut (.I0(n1316), .I1(n5828), .I2(n1293), 
            .I3(GND_net), .O(n1413));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i884_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1062_i40_3_lut (.I0(n32_adj_4669), .I1(n91), 
            .I2(n43_adj_4676), .I3(GND_net), .O(n40_adj_4674));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1062_i28_4_lut (.I0(n658), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28_adj_4665));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35266_3_lut (.I0(n28_adj_4665), .I1(n95), .I2(n35_adj_4671), 
            .I3(GND_net), .O(n42030));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35266_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35267_3_lut (.I0(n42030), .I1(n94), .I2(n37_adj_4672), .I3(GND_net), 
            .O(n42031));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35267_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i883_3_lut_3_lut (.I0(n1316), .I1(n5827), .I2(n1292), 
            .I3(GND_net), .O(n1412));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i883_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33517_4_lut (.I0(n41_adj_4675), .I1(n39_adj_4673), .I2(n37_adj_4672), 
            .I3(n40285), .O(n40279));
    defparam i33517_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35264_4_lut (.I0(n40_adj_4674), .I1(n30_adj_4667), .I2(n43_adj_4676), 
            .I3(n40275), .O(n42028));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35264_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35083_3_lut (.I0(n42031), .I1(n93), .I2(n39_adj_4673), .I3(GND_net), 
            .O(n41847));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35083_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35460_4_lut (.I0(n41847), .I1(n42028), .I2(n43_adj_4676), 
            .I3(n40279), .O(n42224));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35460_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_46_i806_3_lut_3_lut (.I0(n1193), .I1(n5821), .I2(n1173), 
            .I3(GND_net), .O(n1296));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i806_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33597_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n40359));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33597_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i35461_3_lut (.I0(n42224), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n42225));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35461_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n42225), .I1(n15567), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hceef;
    SB_LUT4 i1_2_lut_4_lut_adj_1800 (.I0(n92), .I1(n91), .I2(n90), .I3(n15517), 
            .O(n15504));
    defparam i1_2_lut_4_lut_adj_1800.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4661));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4660));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1801 (.I0(n91), .I1(n90), .I2(n15517), 
            .I3(GND_net), .O(n15561));
    defparam i1_2_lut_3_lut_adj_1801.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i803_3_lut_3_lut (.I0(n1193), .I1(n5818), .I2(n1170), 
            .I3(GND_net), .O(n1293));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i803_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4345), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n657));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1802 (.I0(n89), .I1(n88), .I2(n87), .I3(n15570), 
            .O(n15517));
    defparam i1_2_lut_4_lut_adj_1802.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4664));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1803 (.I0(n88), .I1(n87), .I2(n15570), 
            .I3(GND_net), .O(n15567));
    defparam i1_2_lut_3_lut_adj_1803.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i802_3_lut_3_lut (.I0(n1193), .I1(n5817), .I2(n1169_adj_4409), 
            .I3(GND_net), .O(n1292));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i802_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i807_3_lut_3_lut (.I0(n1193), .I1(n5822), .I2(n1174), 
            .I3(GND_net), .O(n1297));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i807_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1804 (.I0(n86), .I1(n85), .I2(n84), .I3(n15576), 
            .O(n15570));
    defparam i1_2_lut_4_lut_adj_1804.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4636));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4657));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4659));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1805 (.I0(n85), .I1(n84), .I2(n15576), 
            .I3(GND_net), .O(n15526));
    defparam i1_2_lut_3_lut_adj_1805.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1806 (.I0(n83), .I1(n82), .I2(n81), .I3(n15543), 
            .O(n15576));
    defparam i1_2_lut_4_lut_adj_1806.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33624_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n40386));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i33624_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4663));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1807 (.I0(n82), .I1(n81), .I2(n15543), 
            .I3(GND_net), .O(n15530));
    defparam i1_2_lut_3_lut_adj_1807.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4655));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33554_4_lut (.I0(n37_adj_4659), .I1(n35), .I2(n33_adj_4657), 
            .I3(n31_adj_4655), .O(n40316));
    defparam i33554_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_985_i42_3_lut (.I0(n34_adj_4658), .I1(n91), 
            .I2(n45_adj_4664), .I3(GND_net), .O(n42_adj_4662));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_985_i30_4_lut (.I0(n657), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30_adj_4654));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35270_3_lut (.I0(n30_adj_4654), .I1(n95), .I2(n37_adj_4659), 
            .I3(GND_net), .O(n42034));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35270_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35271_3_lut (.I0(n42034), .I1(n94), .I2(n39_adj_4660), .I3(GND_net), 
            .O(n42035));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35271_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33537_4_lut (.I0(n43_adj_4663), .I1(n41_adj_4661), .I2(n39_adj_4660), 
            .I3(n40316), .O(n40299));
    defparam i33537_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34838_4_lut (.I0(n42_adj_4662), .I1(n32_adj_4656), .I2(n45_adj_4664), 
            .I3(n40297), .O(n41602));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34838_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35081_3_lut (.I0(n42035), .I1(n93), .I2(n41_adj_4661), .I3(GND_net), 
            .O(n41845));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35081_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35302_4_lut (.I0(n41845), .I1(n41602), .I2(n45_adj_4664), 
            .I3(n40299), .O(n42066));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35302_4_lut.LUT_INIT = 16'hccca;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n2890({n2891, n2892, n2893, 
            n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
            n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, 
            n2910, n2911, n2912, n2913, n2914}), .encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .n17542(n17542), .clk32MHz(clk32MHz), .n17543(n17543), 
            .n17544(n17544), .n17545(n17545), .n17546(n17546), .n17547(n17547), 
            .n17548(n17548), .n17534(n17534), .n17535(n17535), .n17536(n17536), 
            .n17537(n17537), .n17538(n17538), .n17539(n17539), .n17540(n17540), 
            .n17541(n17541), .n17530(n17530), .n17531(n17531), .n17532(n17532), 
            .n17533(n17533), .n17526(n17526), .n17527(n17527), .n17528(n17528), 
            .n17529(n17529), .data_o({quadA_debounced_adj_4372, quadB_debounced_adj_4373}), 
            .count_enable(count_enable_adj_4374), .n16970(n16970), .n17597(n17597), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B_adj_5064}), .PIN_7_c_1(PIN_7_c_1), 
            .n36606(n36606), .n16990(n16990)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(262[15] 267[4])
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n42066), .I1(n15517), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hceef;
    motorControl control (.VCC_net(VCC_net), .GND_net(GND_net), .\Ki[4] (Ki[4]), 
            .\Kp[3] (Kp[3]), .\Kp[6] (Kp[6]), .\Kp[0] (Kp[0]), .setpoint({setpoint}), 
            .\Kp[4] (Kp[4]), .\Kp[2] (Kp[2]), .\Kp[1] (Kp[1]), .\Kp[5] (Kp[5]), 
            .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Ki[5] (Ki[5]), .\Ki[2] (Ki[2]), 
            .\Ki[3] (Ki[3]), .PWMLimit({PWMLimit}), .\Ki[6] (Ki[6]), .IntegralLimit({IntegralLimit}), 
            .\Ki[7] (Ki[7]), .duty({duty}), .clk32MHz(clk32MHz), .\Kp[7] (Kp[7]), 
            .motor_state({motor_state}), .n25(n25), .n43079(n43079)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(234[16] 247[4])
    SB_LUT4 i1_2_lut_4_lut_adj_1809 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n15543));
    defparam i1_2_lut_4_lut_adj_1809.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1810 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n15546));
    defparam i1_2_lut_3_lut_adj_1810.LUT_INIT = 16'hf7f7;
    \pwm(32000000,20000,32000000,23,1)  PWM (.PIN_19_c_0(PIN_19_c_0), .CLK_c(CLK_c), 
            .\half_duty_new[0] (half_duty_new[0]), .n17573(n17573), .\half_duty[0][7] (\half_duty[0] [7]), 
            .n17567(n17567), .\half_duty[0][1] (\half_duty[0] [1]), .n17568(n17568), 
            .\half_duty[0][2] (\half_duty[0] [2]), .n17569(n17569), .\half_duty[0][3] (\half_duty[0] [3]), 
            .n17570(n17570), .\half_duty[0][4] (\half_duty[0] [4]), .n17572(n17572), 
            .\half_duty[0][6] (\half_duty[0] [6]), .n1169(n1169), .GND_net(GND_net), 
            .VCC_net(VCC_net), .\half_duty_new[1] (half_duty_new[1]), .\half_duty[0][0] (\half_duty[0] [0]), 
            .\half_duty_new[2] (half_duty_new[2]), .\half_duty_new[3] (half_duty_new[3]), 
            .\half_duty_new[4] (half_duty_new[4]), .\half_duty_new[6] (half_duty_new[6]), 
            .\half_duty_new[7] (half_duty_new[7]), .n16982(n16982), .pwm_setpoint({pwm_setpoint})) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(153[43] 159[3])
    SB_LUT4 div_46_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4652));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4649));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4651));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22825_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n511), .I3(n558), 
            .O(n4_adj_4394));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22825_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_46_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4650));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4344), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n656));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22849_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n650), .I3(n558), 
            .O(n4_adj_4476));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22849_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_46_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20187_4_lut (.I0(n954), .I1(n953), .I2(n35536), .I3(n955), 
            .O(n986));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam i20187_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 div_46_LessThan_906_i32_4_lut (.I0(n656), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32_adj_4647));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35276_3_lut (.I0(n32_adj_4647), .I1(n95), .I2(n39_adj_4650), 
            .I3(GND_net), .O(n42040));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35276_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35277_3_lut (.I0(n42040), .I1(n94), .I2(n41_adj_4651), .I3(GND_net), 
            .O(n42041));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35277_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34279_4_lut (.I0(n41_adj_4651), .I1(n39_adj_4650), .I2(n37_adj_4649), 
            .I3(n40346), .O(n41043));
    defparam i34279_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 rem_4_i1195_3_lut (.I0(n1754_adj_4494), .I1(n1821), .I2(n1778_adj_4500), 
            .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(76[6:33])
    defparam rem_4_i1195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34836_3_lut (.I0(n34_adj_4648), .I1(n96), .I2(n37_adj_4649), 
            .I3(GND_net), .O(n41600));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i34836_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35077_3_lut (.I0(n42041), .I1(n93), .I2(n43_adj_4652), .I3(GND_net), 
            .O(n41841));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35077_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35274_4_lut (.I0(n41841), .I1(n41600), .I2(n43_adj_4652), 
            .I3(n41043), .O(n42038));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35274_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35275_3_lut (.I0(n42038), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n42039));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i35275_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n42039), .I1(n15564), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hceef;
    SB_LUT4 i22881_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n651), .I3(n558), 
            .O(n4_adj_4325));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam i22881_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_46_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4646));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4642));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4644));   // verilog/TinyFPGA_B.v(250[21:53])
    defparam div_46_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (VCC_net, timer, \neo_pixel_transmitter.done , clk32MHz, 
            bit_ctr, n40170, GND_net, n11, n33373, n33375, n33361, 
            n33363, n33365, n33367, n33369, n33335, n33377, n33379, 
            n33381, n33383, n33385, n33323, n33371, n33353, n33355, 
            n33357, n33359, n33341, n33343, n33347, n33349, n33351, 
            n33331, n33333, n33329, n33327, n33317, n33319, n33321, 
            \neo_pixel_transmitter.t0 , n40197, n19, n40169, n40168, 
            n40196, n40181, n40180, n40195, n40179, \state_3__N_362[1] , 
            \state[1] , n1163, \state[0] , n4385, n40176, \one_wire_N_513[10] , 
            \one_wire_N_513[8] , \one_wire_N_513[5] , \one_wire_N_513[11] , 
            \one_wire_N_513[7] , \one_wire_N_513[9] , \one_wire_N_513[6] , 
            start, n15464, n35361, n24867, n33325, n17072, n17071, 
            n17070, n17069, n17068, n17067, n17066, n17065, n17064, 
            n17063, n17062, n17061, n17060, n17059, n17058, n17057, 
            n17056, n17055, n35481, n40194, n17054, n17053, n24907, 
            n17052, n17051, n17050, n17049, n17048, n17047, n17046, 
            n37092, n17045, n17044, n17043, n17042, n40175, n16530, 
            n16754, PIN_8_c, n36917, n40172, n40192, n40191, n40190, 
            n40189, n40188, n40187, n40186, n40193, n40185, n40171, 
            n40184, n40199, n33387, n16831, n17017, n40183, n40177, 
            n40198, n40182, n40178, n40174, n40173, n24853, \color[2] , 
            \color[3] , \color[4] , \color[1] ) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input VCC_net;
    output [31:0]timer;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output [31:0]bit_ctr;
    output n40170;
    input GND_net;
    input n11;
    input n33373;
    input n33375;
    input n33361;
    input n33363;
    input n33365;
    input n33367;
    input n33369;
    input n33335;
    input n33377;
    input n33379;
    input n33381;
    input n33383;
    input n33385;
    input n33323;
    input n33371;
    input n33353;
    input n33355;
    input n33357;
    input n33359;
    input n33341;
    input n33343;
    input n33347;
    input n33349;
    input n33351;
    input n33331;
    input n33333;
    input n33329;
    input n33327;
    input n33317;
    input n33319;
    input n33321;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output n40197;
    input n19;
    output n40169;
    output n40168;
    output n40196;
    output n40181;
    output n40180;
    output n40195;
    output n40179;
    output \state_3__N_362[1] ;
    output \state[1] ;
    output n1163;
    output \state[0] ;
    output n4385;
    output n40176;
    output \one_wire_N_513[10] ;
    output \one_wire_N_513[8] ;
    output \one_wire_N_513[5] ;
    output \one_wire_N_513[11] ;
    output \one_wire_N_513[7] ;
    output \one_wire_N_513[9] ;
    output \one_wire_N_513[6] ;
    output start;
    output n15464;
    output n35361;
    output n24867;
    input n33325;
    input n17072;
    input n17071;
    input n17070;
    input n17069;
    input n17068;
    input n17067;
    input n17066;
    input n17065;
    input n17064;
    input n17063;
    input n17062;
    input n17061;
    input n17060;
    input n17059;
    input n17058;
    input n17057;
    input n17056;
    input n17055;
    input n35481;
    output n40194;
    input n17054;
    input n17053;
    output n24907;
    input n17052;
    input n17051;
    input n17050;
    input n17049;
    input n17048;
    input n17047;
    input n17046;
    output n37092;
    input n17045;
    input n17044;
    input n17043;
    input n17042;
    output n40175;
    output n16530;
    output n16754;
    output PIN_8_c;
    input n36917;
    output n40172;
    output n40192;
    output n40191;
    output n40190;
    output n40189;
    output n40188;
    output n40187;
    output n40186;
    output n40193;
    output n40185;
    output n40171;
    output n40184;
    output n40199;
    input n33387;
    input n16831;
    input n17017;
    output n40183;
    output n40177;
    output n40198;
    output n40182;
    output n40178;
    output n40174;
    output n40173;
    output n24853;
    input \color[2] ;
    input \color[3] ;
    input \color[4] ;
    input \color[1] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n29284, n2492, n2522, n29285, n2592, n2493, n29283;
    wire [31:0]n1;
    
    wire n28071, \neo_pixel_transmitter.done_N_570 , n37238, n2593, 
        n2494, n29282, n2594, n2495, n29281, n2595, n2496, n29280, 
        n28246, n1107, n1136, n28247, n2596, n2497, n29279, n1207, 
        n1108, n28245, n2597, n2498, n29278, n2598, n2499, n29277, 
        n2599, n2500, n29276, n1208, n1109, n43073, n28244, n2600, 
        n2501, n29275, n1209, n27894, n2601, n2502, n29274, n2602, 
        n2503, n29273, n2603, n2504, n29272, n2604, n2505, n29271, 
        n2605, n2506, n29270, n2606, n2507, n29269, n27882, n27895, 
        n2607, n2508, n29268, n2608, n2509, n43072, n29267, n1301, 
        n1202, n1235, n28237, n2609, n1302, n1203, n28236, n1303, 
        n1204, n28235, n1304, n1205, n28234, n2489, n2390, n2423, 
        n29266, n2490, n2391, n29265, n1305, n1206, n28233, n1306, 
        n28232, n2491, n2392, n29264, n2393, n29263, n43074, n27893, 
        n1307, n28231, n2394, n29262, n27883, n1308, n28230, n27892, 
        n1309, n2395, n29261, n2396, n29260, n2397, n29259, n2398, 
        n29258, n2399, n29257, n2400, n29256, n2401, n29255, n2402, 
        n29254, n2403, n29253, n1334, n43085, n1806, n1803, n1798, 
        n1805, n24, n1808, n1804, n1802, n1807, n22, n27881, 
        n2404, n29252, n2405, n29251, n1800, n1799, n1797, n1801, 
        n23, n1796, n1809, n21, n2406, n29250, n27891, n2407, 
        n29249, n1829, n1928, n43086, n2408, n29248, n2409, n43075, 
        n29247, n2291, n2324, n29246, n2292, n29245, n2293, n29244, 
        n2294, n29243, n2295, n29242, n2296, n29241, n2297, n29240, 
        n2298, n29239, n2299, n29238, n2300, n29237, n2301, n29236, 
        n2302, n29235, n2303, n29234, n27890, n2304, n29233, n2305, 
        n29232, n2306, n29231, n27880, n2307, n29230, n2308, n29229, 
        n2309, n43076, n29228, n3182, n3083, n3116, n29434, n3183, 
        n3084, n29433, n3184, n3085, n29432, n2192, n2225, n29227, 
        n2193, n29226, n3185, n3086, n29431, n2194, n29225, n3186, 
        n3087, n29430, n2195, n29224, n2196, n29223, n3187, n3088, 
        n29429, n2907, n2909, n33_adj_4186, n2900, n2891, n2897, 
        n2888, n41, n2906, n2887, n2892, n38, n2896, n2885, 
        n2905, n2902, n43, n27, n33_adj_4187, n2899, n2890, n2898, 
        n2908, n40, n2889, n2901, n46, n2886, n2894, n2895, 
        n2903, n39, n2904, n2893, n47, n32, n31, n35, n37, 
        n2918, n1433, n43082, n3188, n3089, n29428, n2197, n29222, 
        n3189, n3090, n29427, n2198, n29221, n2199, n29220, n3190, 
        n3091, n29426, n3191, n3092, n29425, n2200, n29219, n3192, 
        n3093, n29424, n2201, n29218, n2202, n29217, n3193, n3094, 
        n29423, n2203, n29216, n3194, n3095, n29422, n2204, n29215, 
        n27889, n2205, n29214, n3195, n3096, n29421, n2206, n29213, 
        n3196, n3097, n29420, n2207, n29212;
    wire [31:0]n133;
    
    wire n28681, n28680, n2208, n29211, n3197, n3098, n29419, 
        n28679, n3198, n3099, n29418, n28678, n28677, n2209, n43078, 
        n29210, n3199, n3100, n29417, n2093, n2126, n29209, n28676, 
        n2094, n29208, n3200, n3101, n29416, n3201, n3102, n29415, 
        n3202, n3103, n29414, n2095, n29207, n3203, n3104, n29413, 
        n2096, n29206, n3204, n3105, n29412, n2097, n29205, n3205, 
        n3106, n29411, n2098, n29204, n3206, n3107, n29410, n2099, 
        n29203, n3207, n3108, n29409, n3208, n3109, n43077, n29408, 
        n2100, n29202, n3209, n2101, n29201, n28675, n28674, n28673, 
        n2102, n29200, n28672, n2984, n3017, n29407, n2985, n29406, 
        n28671, n28670, n28669, n2103, n29199, n28668, n28667, 
        n2104, n29198, n28666, n2105, n29197, n28665, n2106, n29196, 
        n28664, n2986, n29405, n28663, n1499, n1400, n27999, n1500, 
        n1401, n27998, n28662, n28661, n30, n48, n46_adj_4188, 
        n47_adj_4189, n45, n44, n43_adj_4190, n54, n49, n15466, 
        n4357, n28660, n28659, n28658, n28657, n28656, n1501, 
        n1402, n27997, n28655, n28654, n28653;
    wire [31:0]one_wire_N_513;
    
    wire n30086, n28652, n28651, n2987, n29404, n2107, n29195, 
        n2988, n29403, n2108, n29194, n2989, n29402, n27888, n1502, 
        n1403, n27996, n24891, n4, n10, n15538, n14, n15335, 
        n43081, n2109, n43080, n29193, n2990, n29401, n24268, 
        n1105, n1103, n12, n1106, n1104, n1895, n1902, n1899, 
        n1897, n26, n1907, n1909, n19_adj_4191, n1908, n1900, 
        n16, n1904, n1901, n1906, n1898, n24_adj_4192, n1905, 
        n1903, n28, n1896, n14_adj_4193, n9, n2027, n43084, n34616, 
        n5, n21_adj_4194, n23_adj_4195, n22_adj_4196, n24_adj_4197, 
        n36, n25, n27_adj_4198, n26_adj_4199, n28_adj_4200, n37_adj_4201, 
        n29, n30_adj_4202, n35378, n30241, n34664, n116, n24_adj_4203, 
        n34, n22_adj_4204, n38_adj_4205, n36_adj_4206, n37_adj_4207, 
        n35_adj_4208, n10_adj_4209, n12_adj_4210, n16_adj_4211, n2991, 
        n29400, n1994, n29192, n1995, n29191, n1503, n1404, n27995, 
        n2992, n29399, n1996, n29190, n2993, n29398, n1997, n29189, 
        n2994, n29397, n1998, n29188, n2995, n29396, n1504, n1405, 
        n27994, n1999, n29187, n2996, n29395, n1505, n1406, n27993, 
        n2997, n29394, n2000, n29186, n2998, n29393, n2001, n29185, 
        n2002, n29184, n2003, n29183, n2999, n29392, n2004, n29182, 
        n3000, n29391, n2005, n29181, n3001, n29390, n2006, n29180, 
        n3002, n29389, n2007, n29179, n28110, n3003, n29388, n2008, 
        n29178, n28109, n3004, n29387, n2009, n29177, n3005, n29386, 
        n29176, n29175, n1506, n1407, n27992, n28108, n3006, n29385, 
        n29174, n3007, n29384, n27879, n29173, n29172, n3008, 
        n29383, n29171, n29170, n3009, n29382, n28107, n1507, 
        n1408, n27991, n18, n28_adj_4212, n26_adj_4213, n27_adj_4214, 
        n25_adj_4215, n35367, n35983, n35798, n29169, n28106, n1508, 
        n1409, n27990, n29168, n29381, n29380, n27887, n29167, 
        n29379, n28105, n29166, n29378, n29165, n29377, n28104, 
        n29164, n29376, n1509, n29375, n29163, n29162, n28103, 
        n29374, n29161, n28102, n29160, n29373, n29159, n29372, 
        n29158, n29371, n29370, n29157, n29369, n29156, n29155, 
        n29368, n29154, n29367, n29153, n29366, n29152, n28101, 
        n28100, n29151, n29365, n29150, n29364, n29149, n29363, 
        n43088, n29148, n28099;
    wire [3:0]state_3__N_362;
    
    wire n28098, \neo_pixel_transmitter.done_N_576 , n16544, n27886, 
        n28097, n29362, n28096, n29361, n1697, n1730, n29147, 
        n1698, n29146, n29360, n1699, n29145, n27908, n29359, 
        n1700, n29144, n28095, n29358, n1701, n29143, n28094, 
        n27907, n43087, n29357, n1702, n29142, n1703, n29141, 
        n2786, n2819, n29356, n1704, n29140, n28093, n2787, n29355, 
        n1705, n29139, n27906, n2788, n29354, n1706, n29138, n27905, 
        n2789, n29353, n2790, n29352, n1707, n29137, n27904, n1708, 
        n29136, n27903, n2791, n29351, n1709, n43090, n29135, 
        n27902, n2792, n29350, n27878, n27901, n28092, n2793, 
        n29349, n1598, n1631, n29134, n1599, n29133, n27885, n28091, 
        n2794, n29348, n2795, n29347, n1600, n29132, n2796, n29346, 
        n1601, n29131, n1602, n29130, n2797, n29345, n1603, n29129, 
        n2798, n29344, n1604, n29128, n2799, n29343, n1605, n29127, 
        n2800, n29342, n1606, n29126, n1607, n29125, n28090, n2801, 
        n29341, n2802, n29340, n1608, n29124, n1609, n43092, n29123, 
        n28089, n2803, n29339, n1532, n29122, n2804, n29338, n29121, 
        n27900, n2805, n29337, n29120, n2806, n29336, n27884, 
        n29119, n2807, n29335, n2808, n29334, n29118, n28088, 
        n28087, n2809, n43091, n29333, n29117, n28086, n29116, 
        n29115, n2687, n2720, n29332, n29114, n2688, n29331, n29113, 
        n43093, n29112, n2689, n29330, n2690, n29329, n2691, n29328, 
        n2692, n29327, n2693, n29326, n2694, n29325, n2695, n29324, 
        n2696, n29323, n2697, n29322, n28085, n2698, n29321, n28084, 
        n28083, n2699, n29320, n2700, n29319, n2701, n29318, n2702, 
        n29317, n2703, n29316, n2704, n29315, n2705, n29314, n2706, 
        n29313, n2707, n29312, n2708, n29311, n27899, n2709, n43094, 
        n29310, n2588, n2621, n29309, n2589, n29308, n2590, n29307, 
        n2591, n29306, n29305, n28082, n29304, n29303, n29302, 
        n28081;
    wire [31:0]n971;
    
    wire n905, n28312, n906, n28311, n35441, n28310, n16683, n28309, 
        n14144, n28308, n4_adj_4228, n1037, n28307, n1005, n28306, 
        n1006, n28305, n29301, n1007, n28304, n1008, n28303, n1009, 
        n43096, n28302, n29300, n28080, n29299, n29298, n27898, 
        n29297, n29296, n29295, n28079, n29294, n35321, n14146, 
        n807, n838, n29293, n27897, n29292, n28078, n27896, n29291, 
        n28077, n29290, n28076, n28075, n29289, n28074, n28073, 
        n43095, n29288, n24913, n35437, n28072, n4_adj_4239, n29287, 
        n29286, n28250, n28249, n28248, n24695, n24707, n16_adj_4240, 
        n17_adj_4241, n40_adj_4242, n44_adj_4243, n42, n43_adj_4244, 
        n41_adj_4245, n38_adj_4246, n46_adj_4247, n50, n37_adj_4248, 
        n18_adj_4249, n24689, n30_adj_4250, n28_adj_4251, n29_adj_4252, 
        n27_adj_4253, n28_adj_4254, n32_adj_4255, n30_adj_4256, n31_adj_4257, 
        n29_adj_4258, n42_adj_4259, n46_adj_4260, n44_adj_4261, n45_adj_4262, 
        n43_adj_4263, n40_adj_4264, n48_adj_4265, n52, n39_adj_4266, 
        n22_adj_4267, n30_adj_4268, n34_adj_4269, n32_adj_4270, n33_adj_4271, 
        n31_adj_4272, n31213, n38080, n38082, n6_adj_4273, n60, 
        n608, n708, n35339, n36_adj_4274, n25_adj_4275, n34_adj_4276, 
        n40_adj_4277, n38_adj_4278, n39_adj_4279, n37_adj_4280, n28_adj_4281, 
        n38_adj_4282, n24823, n36_adj_4283, n42_adj_4284, n40_adj_4285, 
        n41_adj_4286, n39_adj_4287, n12_adj_4288, n18_adj_4289, n19_adj_4290, 
        n20_adj_4291, n13_adj_4292, n18_adj_4293, n22_adj_4294, n40_adj_4295, 
        n38_adj_4296, n39_adj_4297, n37_adj_4298, n34_adj_4299, n42_adj_4300, 
        n46_adj_4301, n33_adj_4302, n17_adj_4303, n21_adj_4304, n20_adj_4305, 
        n24_adj_4306, n35457, n24733, n35483, n103, n34539, n24813, 
        n20_adj_4307, n19_adj_4308, n21_adj_4309, n18_adj_4310, n30_adj_4311, 
        n28_adj_4312, n29_adj_4313, n27_adj_4314, n24877, n1166, n4_adj_4315, 
        n2_adj_4316, n4_adj_4317, n41093, n7_adj_4318, n38035;
    
    SB_CARRY mod_5_add_1741_20 (.CI(n29284), .I0(n2492), .I1(n2522), .CO(n29285));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n29283), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n28071));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n37238), .D(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_19 (.CI(n29283), .I0(n2493), .I1(n2522), .CO(n29284));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n29282), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n29282), .I0(n2494), .I1(n2522), .CO(n29283));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n29281), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n29281), .I0(n2495), .I1(n2522), .CO(n29282));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n29280), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n29280), .I0(n2496), .I1(n2522), .CO(n29281));
    SB_CARRY mod_5_add_803_5 (.CI(n28246), .I0(n1107), .I1(n1136), .CO(n28247));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n29279), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n29279), .I0(n2497), .I1(n2522), .CO(n29280));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28245), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n29278), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n29278), .I0(n2498), .I1(n2522), .CO(n29279));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n29277), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n29277), .I0(n2499), .I1(n2522), .CO(n29278));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n29276), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n28245), .I0(n1108), .I1(n1136), .CO(n28246));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n43073), 
            .I3(n28244), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_12 (.CI(n29276), .I0(n2500), .I1(n2522), .CO(n29277));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n29275), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_3 (.CI(n28244), .I0(n1109), .I1(n43073), .CO(n28245));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n43073), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_19_lut (.I0(n11), .I1(bit_ctr[17]), .I2(GND_net), .I3(n27894), 
            .O(n40170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n43073), 
            .CO(n28244));
    SB_CARRY mod_5_add_1741_11 (.CI(n29275), .I0(n2501), .I1(n2522), .CO(n29276));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n29274), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n29274), .I0(n2502), .I1(n2522), .CO(n29275));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n29273), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n29273), .I0(n2503), .I1(n2522), .CO(n29274));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n29272), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n33373));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n33375));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .D(n33361));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n33363));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n33365));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n33367));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n33369));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n33335));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n33377));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n33379));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n33381));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .D(n33383));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n33385));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .D(n33323));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n33371));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n33353));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n33355));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n33357));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n33359));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n33341));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n33343));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n33347));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n33349));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n33351));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .D(n33331));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n33333));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n33329));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n33327));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(VCC_net), 
            .D(n33317));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(VCC_net), 
            .D(n33319));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(VCC_net), 
            .D(n33321));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1741_8 (.CI(n29272), .I0(n2504), .I1(n2522), .CO(n29273));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n29271), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_7 (.CI(n29271), .I0(n2505), .I1(n2522), .CO(n29272));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n29270), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n29270), .I0(n2506), .I1(n2522), .CO(n29271));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n29269), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n29269), .I0(n2507), .I1(n2522), .CO(n29270));
    SB_LUT4 add_21_7_lut (.I0(n19), .I1(bit_ctr[5]), .I2(GND_net), .I3(n27882), 
            .O(n40197)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_19 (.CI(n27894), .I0(bit_ctr[17]), .I1(GND_net), .CO(n27895));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n29268), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n29268), .I0(n2508), .I1(n2522), .CO(n29269));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n43072), 
            .I3(n29267), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_3 (.CI(n29267), .I0(n2509), .I1(n43072), .CO(n29268));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28237), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n43072), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n43072), 
            .CO(n29267));
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28236), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28236), .I0(n1203), .I1(n1235), .CO(n28237));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28235), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n28235), .I0(n1204), .I1(n1235), .CO(n28236));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28234), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n28234), .I0(n1205), .I1(n1235), .CO(n28235));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n29266), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n29265), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28233), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n28233), .I0(n1206), .I1(n1235), .CO(n28234));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28232), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n29265), .I0(n2391), .I1(n2423), .CO(n29266));
    SB_CARRY mod_5_add_870_5 (.CI(n28232), .I0(n1207), .I1(n1235), .CO(n28233));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n29264), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n29264), .I0(n2392), .I1(n2423), .CO(n29265));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n29263), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i36312_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43074));
    defparam i36312_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_18_lut (.I0(n11), .I1(bit_ctr[16]), .I2(GND_net), .I3(n27893), 
            .O(n40169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28231), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n29263), .I0(n2393), .I1(n2423), .CO(n29264));
    SB_CARRY mod_5_add_870_4 (.CI(n28231), .I0(n1208), .I1(n1235), .CO(n28232));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n29262), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_7 (.CI(n27882), .I0(bit_ctr[5]), .I1(GND_net), .CO(n27883));
    SB_CARRY add_21_18 (.CI(n27893), .I0(bit_ctr[16]), .I1(GND_net), .CO(n27894));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n43074), 
            .I3(n28230), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_17_lut (.I0(n11), .I1(bit_ctr[15]), .I2(GND_net), .I3(n27892), 
            .O(n40168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_870_3 (.CI(n28230), .I0(n1209), .I1(n43074), .CO(n28231));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n43074), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n43074), 
            .CO(n28230));
    SB_CARRY mod_5_add_1674_18 (.CI(n29262), .I0(n2394), .I1(n2423), .CO(n29263));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n29261), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n29261), .I0(n2395), .I1(n2423), .CO(n29262));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n29260), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n29260), .I0(n2396), .I1(n2423), .CO(n29261));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n29259), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_17 (.CI(n27892), .I0(bit_ctr[15]), .I1(GND_net), .CO(n27893));
    SB_CARRY mod_5_add_1674_15 (.CI(n29259), .I0(n2397), .I1(n2423), .CO(n29260));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n29258), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n29258), .I0(n2398), .I1(n2423), .CO(n29259));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n29257), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n29257), .I0(n2399), .I1(n2423), .CO(n29258));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n29256), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n29256), .I0(n2400), .I1(n2423), .CO(n29257));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n29255), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n29255), .I0(n2401), .I1(n2423), .CO(n29256));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n29254), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n29254), .I0(n2402), .I1(n2423), .CO(n29255));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n29253), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n29253), .I0(n2403), .I1(n2423), .CO(n29254));
    SB_LUT4 i36323_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43085));
    defparam i36323_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_6_lut (.I0(n19), .I1(bit_ctr[4]), .I2(GND_net), .I3(n27881), 
            .O(n40196)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n29252), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n29252), .I0(n2404), .I1(n2423), .CO(n29253));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n29251), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n29251), .I0(n2405), .I1(n2423), .CO(n29252));
    SB_LUT4 i9_4_lut (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n21));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n29250), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n29250), .I0(n2406), .I1(n2423), .CO(n29251));
    SB_LUT4 add_21_16_lut (.I0(n19), .I1(bit_ctr[14]), .I2(GND_net), .I3(n27891), 
            .O(n40181)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n29249), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut (.I0(n21), .I1(n23), .I2(n22), .I3(n24), .O(n1829));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_5 (.CI(n29249), .I0(n2407), .I1(n2423), .CO(n29250));
    SB_LUT4 i36324_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43086));
    defparam i36324_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n29248), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n29248), .I0(n2408), .I1(n2423), .CO(n29249));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n43075), 
            .I3(n29247), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n29247), .I0(n2409), .I1(n43075), .CO(n29248));
    SB_CARRY add_21_16 (.CI(n27891), .I0(bit_ctr[14]), .I1(GND_net), .CO(n27892));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n43075), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n43075), 
            .CO(n29247));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n29246), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n29245), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n29245), .I0(n2292), .I1(n2324), .CO(n29246));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n29244), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n29244), .I0(n2293), .I1(n2324), .CO(n29245));
    SB_CARRY add_21_6 (.CI(n27881), .I0(bit_ctr[4]), .I1(GND_net), .CO(n27882));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n29243), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n29243), .I0(n2294), .I1(n2324), .CO(n29244));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n29242), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n29242), .I0(n2295), .I1(n2324), .CO(n29243));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n29241), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n29241), .I0(n2296), .I1(n2324), .CO(n29242));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n29240), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n29240), .I0(n2297), .I1(n2324), .CO(n29241));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n29239), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n29239), .I0(n2298), .I1(n2324), .CO(n29240));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n29238), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n29238), .I0(n2299), .I1(n2324), .CO(n29239));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n29237), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n29237), .I0(n2300), .I1(n2324), .CO(n29238));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n29236), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n29236), .I0(n2301), .I1(n2324), .CO(n29237));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n29235), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n29235), .I0(n2302), .I1(n2324), .CO(n29236));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n29234), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n29234), .I0(n2303), .I1(n2324), .CO(n29235));
    SB_LUT4 add_21_15_lut (.I0(n19), .I1(bit_ctr[13]), .I2(GND_net), .I3(n27890), 
            .O(n40180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n29233), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n29233), .I0(n2304), .I1(n2324), .CO(n29234));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n29232), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n29232), .I0(n2305), .I1(n2324), .CO(n29233));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n29231), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_5_lut (.I0(n19), .I1(bit_ctr[3]), .I2(GND_net), .I3(n27880), 
            .O(n40195)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1607_6 (.CI(n29231), .I0(n2306), .I1(n2324), .CO(n29232));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n29230), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n29230), .I0(n2307), .I1(n2324), .CO(n29231));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n29229), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n29229), .I0(n2308), .I1(n2324), .CO(n29230));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n43076), 
            .I3(n29228), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n29228), .I0(n2309), .I1(n43076), .CO(n29229));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n43076), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n29434), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n29433), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n29433), .I0(n3084), .I1(n3116), .CO(n29434));
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n43076), 
            .CO(n29228));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n29432), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n29227), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n29432), .I0(n3085), .I1(n3116), .CO(n29433));
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n29226), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n29431), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n29226), .I0(n2193), .I1(n2225), .CO(n29227));
    SB_CARRY mod_5_add_2143_26 (.CI(n29431), .I0(n3086), .I1(n3116), .CO(n29432));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n29225), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n29430), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n29225), .I0(n2194), .I1(n2225), .CO(n29226));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n29224), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n29430), .I0(n3087), .I1(n3116), .CO(n29431));
    SB_CARRY mod_5_add_1540_17 (.CI(n29224), .I0(n2195), .I1(n2225), .CO(n29225));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n29223), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n29429), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n29223), .I0(n2196), .I1(n2225), .CO(n29224));
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4186));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1460 (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), 
            .I3(GND_net), .O(n27));
    defparam i7_3_lut_adj_1460.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1461 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4187));
    defparam i13_4_lut_adj_1461.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n41), .I1(n33_adj_4186), .I2(n2889), .I3(n2901), 
            .O(n46));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_24 (.CI(n29429), .I0(n3088), .I1(n3116), .CO(n29430));
    SB_LUT4 i14_4_lut (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43), .I1(n2904), .I2(n38), .I3(n2893), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1462 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35));
    defparam i15_4_lut_adj_1462.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n33_adj_4187), .I1(n27), .I2(n2404), .I3(n2401), 
            .O(n37));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39), .I2(n46), .I3(n40), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n35), .I2(n31), .I3(n32), .O(n2423));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36320_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43082));
    defparam i36320_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n29428), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n29222), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n29428), .I0(n3089), .I1(n3116), .CO(n29429));
    SB_CARRY mod_5_add_1540_15 (.CI(n29222), .I0(n2197), .I1(n2225), .CO(n29223));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n29427), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n29221), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_15 (.CI(n27890), .I0(bit_ctr[13]), .I1(GND_net), .CO(n27891));
    SB_CARRY mod_5_add_1540_14 (.CI(n29221), .I0(n2198), .I1(n2225), .CO(n29222));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n29220), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n29427), .I0(n3090), .I1(n3116), .CO(n29428));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n29426), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n29426), .I0(n3091), .I1(n3116), .CO(n29427));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n29425), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n29220), .I0(n2199), .I1(n2225), .CO(n29221));
    SB_CARRY mod_5_add_2143_20 (.CI(n29425), .I0(n3092), .I1(n3116), .CO(n29426));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n29219), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n29219), .I0(n2200), .I1(n2225), .CO(n29220));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n29424), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n29424), .I0(n3093), .I1(n3116), .CO(n29425));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n29218), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n29218), .I0(n2201), .I1(n2225), .CO(n29219));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n29217), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n29217), .I0(n2202), .I1(n2225), .CO(n29218));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n29423), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n29216), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n29423), .I0(n3094), .I1(n3116), .CO(n29424));
    SB_CARRY mod_5_add_1540_9 (.CI(n29216), .I0(n2203), .I1(n2225), .CO(n29217));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n29422), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n29215), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n29215), .I0(n2204), .I1(n2225), .CO(n29216));
    SB_LUT4 add_21_14_lut (.I0(n19), .I1(bit_ctr[12]), .I2(GND_net), .I3(n27889), 
            .O(n40179)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n29214), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n29422), .I0(n3095), .I1(n3116), .CO(n29423));
    SB_CARRY mod_5_add_1540_7 (.CI(n29214), .I0(n2205), .I1(n2225), .CO(n29215));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n29421), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n29213), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n29421), .I0(n3096), .I1(n3116), .CO(n29422));
    SB_CARRY mod_5_add_1540_6 (.CI(n29213), .I0(n2206), .I1(n2225), .CO(n29214));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n29420), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n29212), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n28681), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_5 (.CI(n29212), .I0(n2207), .I1(n2225), .CO(n29213));
    SB_LUT4 timer_1177_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n28680), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_15 (.CI(n29420), .I0(n3097), .I1(n3116), .CO(n29421));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n29211), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1177_add_4_32 (.CI(n28680), .I0(GND_net), .I1(timer[30]), 
            .CO(n28681));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n29419), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n28679), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_31 (.CI(n28679), .I0(GND_net), .I1(timer[29]), 
            .CO(n28680));
    SB_CARRY mod_5_add_2143_14 (.CI(n29419), .I0(n3098), .I1(n3116), .CO(n29420));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n29418), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n28678), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_13 (.CI(n29418), .I0(n3099), .I1(n3116), .CO(n29419));
    SB_CARRY mod_5_add_1540_4 (.CI(n29211), .I0(n2208), .I1(n2225), .CO(n29212));
    SB_CARRY timer_1177_add_4_30 (.CI(n28678), .I0(GND_net), .I1(timer[28]), 
            .CO(n28679));
    SB_LUT4 timer_1177_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n28677), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n43078), 
            .I3(n29210), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n29210), .I0(n2209), .I1(n43078), .CO(n29211));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n43078), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n29417), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1177_add_4_29 (.CI(n28677), .I0(GND_net), .I1(timer[27]), 
            .CO(n28678));
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n43078), 
            .CO(n29210));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n29209), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n28676), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n29208), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n29417), .I0(n3100), .I1(n3116), .CO(n29418));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n29416), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n29208), .I0(n2094), .I1(n2126), .CO(n29209));
    SB_CARRY mod_5_add_2143_11 (.CI(n29416), .I0(n3101), .I1(n3116), .CO(n29417));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n29415), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n29415), .I0(n3102), .I1(n3116), .CO(n29416));
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n29414), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n29207), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n29414), .I0(n3103), .I1(n3116), .CO(n29415));
    SB_CARRY mod_5_add_1473_17 (.CI(n29207), .I0(n2095), .I1(n2126), .CO(n29208));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n29413), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n29206), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n29413), .I0(n3104), .I1(n3116), .CO(n29414));
    SB_CARRY mod_5_add_1473_16 (.CI(n29206), .I0(n2096), .I1(n2126), .CO(n29207));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n29412), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n29205), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n29412), .I0(n3105), .I1(n3116), .CO(n29413));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n29411), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n29205), .I0(n2097), .I1(n2126), .CO(n29206));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n29204), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n29204), .I0(n2098), .I1(n2126), .CO(n29205));
    SB_CARRY mod_5_add_2143_6 (.CI(n29411), .I0(n3106), .I1(n3116), .CO(n29412));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n29410), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n29410), .I0(n3107), .I1(n3116), .CO(n29411));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n29203), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n29409), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n29409), .I0(n3108), .I1(n3116), .CO(n29410));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n43077), 
            .I3(n29408), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_13 (.CI(n29203), .I0(n2099), .I1(n2126), .CO(n29204));
    SB_CARRY timer_1177_add_4_28 (.CI(n28676), .I0(GND_net), .I1(timer[26]), 
            .CO(n28677));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n29202), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_3 (.CI(n29408), .I0(n3109), .I1(n43077), .CO(n29409));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n43077), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_12 (.CI(n29202), .I0(n2100), .I1(n2126), .CO(n29203));
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n43077), 
            .CO(n29408));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n29201), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n28675), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_11 (.CI(n29201), .I0(n2101), .I1(n2126), .CO(n29202));
    SB_CARRY timer_1177_add_4_27 (.CI(n28675), .I0(GND_net), .I1(timer[25]), 
            .CO(n28676));
    SB_LUT4 timer_1177_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n28674), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_26 (.CI(n28674), .I0(GND_net), .I1(timer[24]), 
            .CO(n28675));
    SB_LUT4 timer_1177_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n28673), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_25 (.CI(n28673), .I0(GND_net), .I1(timer[23]), 
            .CO(n28674));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n29200), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n28672), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_24 (.CI(n28672), .I0(GND_net), .I1(timer[22]), 
            .CO(n28673));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n29407), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n29406), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n29200), .I0(n2102), .I1(n2126), .CO(n29201));
    SB_LUT4 timer_1177_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n28671), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_23 (.CI(n28671), .I0(GND_net), .I1(timer[21]), 
            .CO(n28672));
    SB_LUT4 timer_1177_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n28670), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_22 (.CI(n28670), .I0(GND_net), .I1(timer[20]), 
            .CO(n28671));
    SB_LUT4 timer_1177_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n28669), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n29199), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n29406), .I0(n2985), .I1(n3017), .CO(n29407));
    SB_CARRY mod_5_add_1473_9 (.CI(n29199), .I0(n2103), .I1(n2126), .CO(n29200));
    SB_CARRY timer_1177_add_4_21 (.CI(n28669), .I0(GND_net), .I1(timer[19]), 
            .CO(n28670));
    SB_LUT4 timer_1177_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n28668), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_20 (.CI(n28668), .I0(GND_net), .I1(timer[18]), 
            .CO(n28669));
    SB_LUT4 timer_1177_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n28667), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n29198), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n29198), .I0(n2104), .I1(n2126), .CO(n29199));
    SB_CARRY timer_1177_add_4_19 (.CI(n28667), .I0(GND_net), .I1(timer[17]), 
            .CO(n28668));
    SB_LUT4 timer_1177_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n28666), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_18 (.CI(n28666), .I0(GND_net), .I1(timer[16]), 
            .CO(n28667));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n29197), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n28665), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_7 (.CI(n29197), .I0(n2105), .I1(n2126), .CO(n29198));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n29196), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1177_add_4_17 (.CI(n28665), .I0(GND_net), .I1(timer[15]), 
            .CO(n28666));
    SB_LUT4 timer_1177_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n28664), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_16 (.CI(n28664), .I0(GND_net), .I1(timer[14]), 
            .CO(n28665));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n29405), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n28663), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n27999), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1177_add_4_15 (.CI(n28663), .I0(GND_net), .I1(timer[13]), 
            .CO(n28664));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n27998), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n28662), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_14 (.CI(n28662), .I0(GND_net), .I1(timer[12]), 
            .CO(n28663));
    SB_LUT4 timer_1177_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n28661), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1463 (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46_adj_4188));
    defparam i18_4_lut_adj_1463.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1464 (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47_adj_4189));
    defparam i19_4_lut_adj_1464.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1465 (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut_adj_1465.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1466 (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i16_4_lut_adj_1466.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1467 (.I0(bit_ctr[3]), .I1(n30), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43_adj_4190));
    defparam i15_4_lut_adj_1467.LUT_INIT = 16'hfefc;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47_adj_4189), .I2(n46_adj_4188), 
            .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1468 (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut_adj_1468.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43_adj_4190), .I3(n44), 
            .O(\state_3__N_362[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2039_3_lut (.I0(n15466), .I1(\state_3__N_362[1] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n4357));
    defparam i2039_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14_4_lut_adj_1469 (.I0(n1163), .I1(n4357), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n4385));
    defparam i14_4_lut_adj_1469.LUT_INIT = 16'hcfca;
    SB_CARRY timer_1177_add_4_13 (.CI(n28661), .I0(GND_net), .I1(timer[11]), 
            .CO(n28662));
    SB_CARRY mod_5_add_1004_11 (.CI(n27998), .I0(n1401), .I1(n1433), .CO(n27999));
    SB_DFF timer_1177__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 timer_1177_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n28660), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_12 (.CI(n28660), .I0(GND_net), .I1(timer[10]), 
            .CO(n28661));
    SB_LUT4 timer_1177_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n28659), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_11 (.CI(n28659), .I0(GND_net), .I1(timer[9]), 
            .CO(n28660));
    SB_LUT4 timer_1177_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n28658), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_10 (.CI(n28658), .I0(GND_net), .I1(timer[8]), 
            .CO(n28659));
    SB_LUT4 timer_1177_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n28657), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_9 (.CI(n28657), .I0(GND_net), .I1(timer[7]), 
            .CO(n28658));
    SB_LUT4 timer_1177_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n28656), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_26 (.CI(n29405), .I0(n2986), .I1(n3017), .CO(n29406));
    SB_CARRY timer_1177_add_4_8 (.CI(n28656), .I0(GND_net), .I1(timer[6]), 
            .CO(n28657));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n27997), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n28655), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_7 (.CI(n28655), .I0(GND_net), .I1(timer[5]), 
            .CO(n28656));
    SB_LUT4 timer_1177_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n28654), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_6 (.CI(n28654), .I0(GND_net), .I1(timer[4]), 
            .CO(n28655));
    SB_LUT4 timer_1177_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n28653), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1177_add_4_5 (.CI(n28653), .I0(GND_net), .I1(timer[3]), 
            .CO(n28654));
    SB_LUT4 i2_3_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[4]), .I2(one_wire_N_513[2]), 
            .I3(GND_net), .O(n30086));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_CARRY mod_5_add_1004_10 (.CI(n27997), .I0(n1402), .I1(n1433), .CO(n27998));
    SB_LUT4 timer_1177_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n28652), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_14 (.CI(n27889), .I0(bit_ctr[12]), .I1(GND_net), .CO(n27890));
    SB_CARRY timer_1177_add_4_4 (.CI(n28652), .I0(GND_net), .I1(timer[2]), 
            .CO(n28653));
    SB_LUT4 timer_1177_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n28651), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n29404), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n29196), .I0(n2106), .I1(n2126), .CO(n29197));
    SB_CARRY timer_1177_add_4_3 (.CI(n28651), .I0(GND_net), .I1(timer[1]), 
            .CO(n28652));
    SB_CARRY mod_5_add_2076_25 (.CI(n29404), .I0(n2987), .I1(n3017), .CO(n29405));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n29195), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1177_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1177_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n29403), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n29195), .I0(n2107), .I1(n2126), .CO(n29196));
    SB_CARRY timer_1177_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n28651));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n29194), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n29403), .I0(n2988), .I1(n3017), .CO(n29404));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n29402), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_13_lut (.I0(n19), .I1(bit_ctr[11]), .I2(GND_net), .I3(n27888), 
            .O(n40176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n27996), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut (.I0(n24891), .I1(one_wire_N_513[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1470 (.I0(\one_wire_N_513[10] ), .I1(\one_wire_N_513[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/neopixel.v(62[15:42])
    defparam i2_2_lut_adj_1470.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(\one_wire_N_513[5] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[7] ), .I3(n15538), .O(n14));   // verilog/neopixel.v(62[15:42])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(\one_wire_N_513[9] ), .I1(n14), .I2(n10), .I3(\one_wire_N_513[6] ), 
            .O(n15335));   // verilog/neopixel.v(62[15:42])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_326_i8_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n15464));
    defparam equal_326_i8_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i28665_2_lut (.I0(\state[1] ), .I1(n15466), .I2(GND_net), 
            .I3(GND_net), .O(n35361));
    defparam i28665_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20209_2_lut (.I0(n30086), .I1(n15335), .I2(GND_net), .I3(GND_net), 
            .O(n24867));
    defparam i20209_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i36311_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43073));
    defparam i36311_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36319_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43081));
    defparam i36319_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_23 (.CI(n29402), .I0(n2989), .I1(n3017), .CO(n29403));
    SB_CARRY mod_5_add_1473_4 (.CI(n29194), .I0(n2108), .I1(n2126), .CO(n29195));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n43080), 
            .I3(n29193), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n29193), .I0(n2109), .I1(n43080), .CO(n29194));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n29401), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .D(n33325));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n17072));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n17071));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n17070));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n17069));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n17068));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n17067));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n17066));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n17065));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n17064));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n17063));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n17062));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n17061));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n17060));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n17059));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n17058));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n17057));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n17056));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n17055));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2076_22 (.CI(n29401), .I0(n2990), .I1(n3017), .CO(n29402));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n43080), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_5 (.CI(n27880), .I0(bit_ctr[3]), .I1(GND_net), .CO(n27881));
    SB_LUT4 i19613_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n24268));
    defparam i19613_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n24268), .I3(n1108), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1471 (.I0(n1107), .I1(n12), .I2(n1106), .I3(n1104), 
            .O(n1136));
    defparam i6_4_lut_adj_1471.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1472 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26));
    defparam i11_4_lut_adj_1472.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), .I3(GND_net), 
            .O(n19_adj_4191));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16));
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1474 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4192));
    defparam i9_4_lut_adj_1474.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1475 (.I0(n19_adj_4191), .I1(n26), .I2(n1905), 
            .I3(n1903), .O(n28));
    defparam i13_4_lut_adj_1475.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1476 (.I0(n1896), .I1(n28), .I2(n24_adj_4192), 
            .I3(n16), .O(n1928));
    defparam i14_4_lut_adj_1476.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1477 (.I0(n1205), .I1(n1208), .I2(n1202), .I3(n1206), 
            .O(n14_adj_4193));
    defparam i6_4_lut_adj_1477.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[23]), .I1(n1207), .I2(n1209), .I3(GND_net), 
            .O(n9));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1004_9 (.CI(n27996), .I0(n1403), .I1(n1433), .CO(n27997));
    SB_LUT4 i36322_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43084));
    defparam i36322_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n34616));
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n5));
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'heeee;
    SB_LUT4 i16_4_lut_adj_1480 (.I0(n21_adj_4194), .I1(n23_adj_4195), .I2(n22_adj_4196), 
            .I3(n24_adj_4197), .O(n36));   // verilog/neopixel.v(62[15:42])
    defparam i16_4_lut_adj_1480.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1481 (.I0(n25), .I1(n27_adj_4198), .I2(n26_adj_4199), 
            .I3(n28_adj_4200), .O(n37_adj_4201));   // verilog/neopixel.v(62[15:42])
    defparam i17_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1482 (.I0(n37_adj_4201), .I1(n29), .I2(n36), 
            .I3(n30_adj_4202), .O(n15538));   // verilog/neopixel.v(62[15:42])
    defparam i19_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 i28679_2_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[2]), 
            .I2(GND_net), .I3(GND_net), .O(n35378));
    defparam i28679_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20232_2_lut (.I0(n30241), .I1(one_wire_N_513[3]), .I2(GND_net), 
            .I3(GND_net), .O(n24891));
    defparam i20232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(one_wire_N_513[4]), .I1(n34664), .I2(n24891), 
            .I3(n35378), .O(n116));
    defparam i1_4_lut.LUT_INIT = 16'h45cd;
    SB_LUT4 i36295_3_lut (.I0(n35481), .I1(n116), .I2(n15538), .I3(GND_net), 
            .O(n37238));
    defparam i36295_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut (.I0(n2503), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4203));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1483 (.I0(n2496), .I1(n2502), .I2(n2491), .I3(n2490), 
            .O(n34));
    defparam i13_4_lut_adj_1483.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1484 (.I0(n2489), .I1(bit_ctr[10]), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4204));
    defparam i1_3_lut_adj_1484.LUT_INIT = 16'heaea;
    SB_LUT4 i17_4_lut_adj_1485 (.I0(n2492), .I1(n34), .I2(n24_adj_4203), 
            .I3(n2494), .O(n38_adj_4205));
    defparam i17_4_lut_adj_1485.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1486 (.I0(n2501), .I1(n2499), .I2(n2495), .I3(n2505), 
            .O(n36_adj_4206));
    defparam i15_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1487 (.I0(n2497), .I1(n2506), .I2(n2493), .I3(n22_adj_4204), 
            .O(n37_adj_4207));
    defparam i16_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1488 (.I0(n2507), .I1(n2498), .I2(n2500), .I3(n2508), 
            .O(n35_adj_4208));
    defparam i14_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1489 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4209));
    defparam i1_2_lut_adj_1489.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12_adj_4210));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1490 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4209), 
            .O(n16_adj_4211));
    defparam i7_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1491 (.I0(n1307), .I1(n16_adj_4211), .I2(n12_adj_4210), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n29400), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n43080), 
            .CO(n29193));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n29192), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n29400), .I0(n2991), .I1(n3017), .CO(n29401));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n29191), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n27995), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n29191), .I0(n1995), .I1(n2027), .CO(n29192));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n29399), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n29190), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n29399), .I0(n2992), .I1(n3017), .CO(n29400));
    SB_CARRY mod_5_add_1406_16 (.CI(n29190), .I0(n1996), .I1(n2027), .CO(n29191));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n29398), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n29189), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n29398), .I0(n2993), .I1(n3017), .CO(n29399));
    SB_LUT4 i20_4_lut_adj_1492 (.I0(n35_adj_4208), .I1(n37_adj_4207), .I2(n36_adj_4206), 
            .I3(n38_adj_4205), .O(n2522));
    defparam i20_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n29397), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n29189), .I0(n1997), .I1(n2027), .CO(n29190));
    SB_CARRY mod_5_add_1004_8 (.CI(n27995), .I0(n1404), .I1(n1433), .CO(n27996));
    SB_CARRY mod_5_add_2076_18 (.CI(n29397), .I0(n2994), .I1(n3017), .CO(n29398));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n29188), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n29396), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n29188), .I0(n1998), .I1(n2027), .CO(n29189));
    SB_CARRY mod_5_add_2076_17 (.CI(n29396), .I0(n2995), .I1(n3017), .CO(n29397));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n27994), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n27994), .I0(n1405), .I1(n1433), .CO(n27995));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n29187), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n29395), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n29187), .I0(n1999), .I1(n2027), .CO(n29188));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n27993), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n29395), .I0(n2996), .I1(n3017), .CO(n29396));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n29394), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n29186), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n29394), .I0(n2997), .I1(n3017), .CO(n29395));
    SB_CARRY mod_5_add_1004_6 (.CI(n27993), .I0(n1406), .I1(n1433), .CO(n27994));
    SB_CARRY mod_5_add_1406_12 (.CI(n29186), .I0(n2000), .I1(n2027), .CO(n29187));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n29393), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n29185), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n29185), .I0(n2001), .I1(n2027), .CO(n29186));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n29184), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n29393), .I0(n2998), .I1(n3017), .CO(n29394));
    SB_CARRY mod_5_add_1406_10 (.CI(n29184), .I0(n2002), .I1(n2027), .CO(n29185));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n29183), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n29392), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n29183), .I0(n2003), .I1(n2027), .CO(n29184));
    SB_CARRY mod_5_add_2076_13 (.CI(n29392), .I0(n2999), .I1(n3017), .CO(n29393));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n29182), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_13 (.CI(n27888), .I0(bit_ctr[11]), .I1(GND_net), .CO(n27889));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n29391), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n29182), .I0(n2004), .I1(n2027), .CO(n29183));
    SB_CARRY mod_5_add_2076_12 (.CI(n29391), .I0(n3000), .I1(n3017), .CO(n29392));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n29181), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n29390), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n29181), .I0(n2005), .I1(n2027), .CO(n29182));
    SB_CARRY mod_5_add_2076_11 (.CI(n29390), .I0(n3001), .I1(n3017), .CO(n29391));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n29180), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n29389), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n29180), .I0(n2006), .I1(n2027), .CO(n29181));
    SB_CARRY mod_5_add_2076_10 (.CI(n29389), .I0(n3002), .I1(n3017), .CO(n29390));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n29179), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28110), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n29388), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n29388), .I0(n3003), .I1(n3017), .CO(n29389));
    SB_CARRY mod_5_add_1406_5 (.CI(n29179), .I0(n2007), .I1(n2027), .CO(n29180));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n29178), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28109), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n29387), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n29178), .I0(n2008), .I1(n2027), .CO(n29179));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n43084), 
            .I3(n29177), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_8 (.CI(n29387), .I0(n3004), .I1(n3017), .CO(n29388));
    SB_CARRY mod_5_add_1406_3 (.CI(n29177), .I0(n2009), .I1(n43084), .CO(n29178));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n43084), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n29386), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n43084), 
            .CO(n29177));
    SB_CARRY mod_5_add_2076_7 (.CI(n29386), .I0(n3005), .I1(n3017), .CO(n29387));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n29176), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n29175), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n28109), .I0(n1302), .I1(n1334), .CO(n28110));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n27992), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28108), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n28108), .I0(n1303), .I1(n1334), .CO(n28109));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n29385), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n29175), .I0(n1896), .I1(n1928), .CO(n29176));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n29174), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n29385), .I0(n3006), .I1(n3017), .CO(n29386));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n29384), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n29174), .I0(n1897), .I1(n1928), .CO(n29175));
    SB_LUT4 add_21_4_lut (.I0(n19), .I1(bit_ctr[2]), .I2(GND_net), .I3(n27879), 
            .O(n40194)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n29173), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n27992), .I0(n1407), .I1(n1433), .CO(n27993));
    SB_CARRY mod_5_add_1339_14 (.CI(n29173), .I0(n1898), .I1(n1928), .CO(n29174));
    SB_CARRY mod_5_add_2076_5 (.CI(n29384), .I0(n3007), .I1(n3017), .CO(n29385));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n29172), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n29172), .I0(n1899), .I1(n1928), .CO(n29173));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n29383), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n29171), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n29383), .I0(n3008), .I1(n3017), .CO(n29384));
    SB_CARRY mod_5_add_1339_12 (.CI(n29171), .I0(n1900), .I1(n1928), .CO(n29172));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n29170), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1493 (.I0(n9), .I1(n14_adj_4193), .I2(n1203), 
            .I3(n1204), .O(n1235));
    defparam i7_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i36310_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43072));
    defparam i36310_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n43081), 
            .I3(n29382), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n17054));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1339_11 (.CI(n29170), .I0(n1901), .I1(n1928), .CO(n29171));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28107), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n27991), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_3 (.CI(n29382), .I0(n3009), .I1(n43081), .CO(n29383));
    SB_CARRY mod_5_add_937_8 (.CI(n28107), .I0(n1304), .I1(n1334), .CO(n28108));
    SB_LUT4 i2_2_lut_adj_1494 (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i2_2_lut_adj_1494.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1495 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28_adj_4212));
    defparam i12_4_lut_adj_1495.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1496 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26_adj_4213));
    defparam i10_4_lut_adj_1496.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1497 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4214));
    defparam i11_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1498 (.I0(bit_ctr[15]), .I1(n18), .I2(n2006), 
            .I3(n2009), .O(n25_adj_4215));
    defparam i9_4_lut_adj_1498.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1499 (.I0(n25_adj_4215), .I1(n27_adj_4214), .I2(n26_adj_4213), 
            .I3(n28_adj_4212), .O(n2027));
    defparam i15_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n17053));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i28747_4_lut (.I0(n15335), .I1(n30086), .I2(n4), .I3(\state[0] ), 
            .O(n24907));
    defparam i28747_4_lut.LUT_INIT = 16'hfaee;
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n17052));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n17051));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n17050));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n17049));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n17048));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i3_4_lut (.I0(n5), .I1(\state[1] ), .I2(n15335), .I3(n35367), 
            .O(n35983));
    defparam i3_4_lut.LUT_INIT = 16'heeef;
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n17047));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n17046));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i2_4_lut (.I0(\state[1] ), .I1(n35983), .I2(start), .I3(n35798), 
            .O(n37092));
    defparam i2_4_lut.LUT_INIT = 16'h8c00;
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n17045));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n17044));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n17043));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n17042));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n29169), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n27991), .I0(n1408), .I1(n1433), .CO(n27992));
    SB_CARRY mod_5_add_1339_10 (.CI(n29169), .I0(n1902), .I1(n1928), .CO(n29170));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n43081), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28106), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n28106), .I0(n1305), .I1(n1334), .CO(n28107));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n43082), 
            .I3(n27990), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n29168), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_3 (.CI(n27990), .I0(n1409), .I1(n43082), .CO(n27991));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n43081), 
            .CO(n29382));
    SB_CARRY mod_5_add_1339_9 (.CI(n29168), .I0(n1903), .I1(n1928), .CO(n29169));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n29381), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i36318_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43080));
    defparam i36318_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n29380), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n29380), .I0(n2886), .I1(n2918), .CO(n29381));
    SB_LUT4 add_21_12_lut (.I0(n19), .I1(bit_ctr[10]), .I2(GND_net), .I3(n27887), 
            .O(n40175)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n29167), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n29379), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n29167), .I0(n1904), .I1(n1928), .CO(n29168));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28105), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n29166), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n28105), .I0(n1306), .I1(n1334), .CO(n28106));
    SB_CARRY mod_5_add_2009_25 (.CI(n29379), .I0(n2887), .I1(n2918), .CO(n29380));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n29378), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n29166), .I0(n1905), .I1(n1928), .CO(n29167));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n29165), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n29378), .I0(n2888), .I1(n2918), .CO(n29379));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n29377), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28104), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n29165), .I0(n1906), .I1(n1928), .CO(n29166));
    SB_CARRY mod_5_add_937_5 (.CI(n28104), .I0(n1307), .I1(n1334), .CO(n28105));
    SB_CARRY mod_5_add_2009_23 (.CI(n29377), .I0(n2889), .I1(n2918), .CO(n29378));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n29164), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n29376), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n29164), .I0(n1907), .I1(n1928), .CO(n29165));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n43082), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_22 (.CI(n29376), .I0(n2890), .I1(n2918), .CO(n29377));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n29375), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n29163), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n29163), .I0(n1908), .I1(n1928), .CO(n29164));
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n43082), 
            .CO(n27990));
    SB_CARRY add_21_12 (.CI(n27887), .I0(bit_ctr[10]), .I1(GND_net), .CO(n27888));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n43086), 
            .I3(n29162), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_21 (.CI(n29375), .I0(n2891), .I1(n2918), .CO(n29376));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28103), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n29374), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n29374), .I0(n2892), .I1(n2918), .CO(n29375));
    SB_CARRY mod_5_add_1339_3 (.CI(n29162), .I0(n1909), .I1(n43086), .CO(n29163));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n43086), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n43086), 
            .CO(n29162));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n29161), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n28103), .I0(n1308), .I1(n1334), .CO(n28104));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n43085), 
            .I3(n28102), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n29160), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n29373), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n29160), .I0(n1797), .I1(n1829), .CO(n29161));
    SB_CARRY mod_5_add_2009_19 (.CI(n29373), .I0(n2893), .I1(n2918), .CO(n29374));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n29159), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n29372), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n29159), .I0(n1798), .I1(n1829), .CO(n29160));
    SB_CARRY mod_5_add_2009_18 (.CI(n29372), .I0(n2894), .I1(n2918), .CO(n29373));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n29158), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_3 (.CI(n28102), .I0(n1309), .I1(n43085), .CO(n28103));
    SB_CARRY mod_5_add_1272_13 (.CI(n29158), .I0(n1799), .I1(n1829), .CO(n29159));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n29371), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_4 (.CI(n27879), .I0(bit_ctr[2]), .I1(GND_net), .CO(n27880));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n43085), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_17 (.CI(n29371), .I0(n2895), .I1(n2918), .CO(n29372));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n29370), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n29370), .I0(n2896), .I1(n2918), .CO(n29371));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n29157), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n29157), .I0(n1800), .I1(n1829), .CO(n29158));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n29369), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n29156), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n29156), .I0(n1801), .I1(n1829), .CO(n29157));
    SB_CARRY mod_5_add_2009_15 (.CI(n29369), .I0(n2897), .I1(n2918), .CO(n29370));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n29155), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n29155), .I0(n1802), .I1(n1829), .CO(n29156));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n29368), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n29154), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n29368), .I0(n2898), .I1(n2918), .CO(n29369));
    SB_CARRY mod_5_add_1272_9 (.CI(n29154), .I0(n1803), .I1(n1829), .CO(n29155));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n29367), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n29153), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n29367), .I0(n2899), .I1(n2918), .CO(n29368));
    SB_CARRY mod_5_add_1272_8 (.CI(n29153), .I0(n1804), .I1(n1829), .CO(n29154));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n29366), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n29152), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n43085), 
            .CO(n28102));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_513[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n28101), .O(n22_adj_4196)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_513[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n28100), .O(n23_adj_4195)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1272_7 (.CI(n29152), .I0(n1805), .I1(n1829), .CO(n29153));
    SB_CARRY sub_14_add_2_32 (.CI(n28100), .I0(timer[30]), .I1(n1[30]), 
            .CO(n28101));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n29151), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n29366), .I0(n2900), .I1(n2918), .CO(n29367));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n29365), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n29365), .I0(n2901), .I1(n2918), .CO(n29366));
    SB_CARRY mod_5_add_1272_6 (.CI(n29151), .I0(n1806), .I1(n1829), .CO(n29152));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n29150), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n29364), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n29150), .I0(n1807), .I1(n1829), .CO(n29151));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n29149), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n29364), .I0(n2902), .I1(n2918), .CO(n29365));
    SB_CARRY mod_5_add_1272_4 (.CI(n29149), .I0(n1808), .I1(n1829), .CO(n29150));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n29363), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n29363), .I0(n2903), .I1(n2918), .CO(n29364));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n43088), 
            .I3(n29148), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_513[19]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n28099), .O(n28_adj_4200)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n28099), .I0(timer[29]), .I1(n1[29]), 
            .CO(n28100));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n16530), .D(state_3__N_362[0]), 
            .S(n16754));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_513[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n28098), .O(n26_adj_4199)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n28098), .I0(timer[28]), .I1(n1[28]), 
            .CO(n28099));
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n16544), .D(\neo_pixel_transmitter.done_N_576 ), 
            .R(n36917));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_11_lut (.I0(n11), .I1(bit_ctr[9]), .I2(GND_net), .I3(n27886), 
            .O(n40172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_513[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n28097), .O(n21_adj_4194)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n28097), .I0(timer[27]), .I1(n1[27]), 
            .CO(n28098));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n29362), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n28096), .O(one_wire_N_513[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_8 (.CI(n29362), .I0(n2904), .I1(n2918), .CO(n29363));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n29361), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_3 (.CI(n29148), .I0(n1809), .I1(n43088), .CO(n29149));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n43088), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_28 (.CI(n28096), .I0(timer[26]), .I1(n1[26]), 
            .CO(n28097));
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n43088), 
            .CO(n29148));
    SB_CARRY mod_5_add_2009_7 (.CI(n29361), .I0(n2905), .I1(n2918), .CO(n29362));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n29147), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n29146), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n29360), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n29146), .I0(n1698), .I1(n1730), .CO(n29147));
    SB_CARRY mod_5_add_2009_6 (.CI(n29360), .I0(n2906), .I1(n2918), .CO(n29361));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n29145), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n29145), .I0(n1699), .I1(n1730), .CO(n29146));
    SB_LUT4 add_21_33_lut (.I0(n19), .I1(bit_ctr[31]), .I2(GND_net), .I3(n27908), 
            .O(n40192)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n29359), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n29144), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n29359), .I0(n2907), .I1(n2918), .CO(n29360));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n28095), .O(one_wire_N_513[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n29358), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n29144), .I0(n1700), .I1(n1730), .CO(n29145));
    SB_CARRY sub_14_add_2_27 (.CI(n28095), .I0(timer[25]), .I1(n1[25]), 
            .CO(n28096));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n29143), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n28094), .O(one_wire_N_513[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n29358), .I0(n2908), .I1(n2918), .CO(n29359));
    SB_CARRY mod_5_add_1205_11 (.CI(n29143), .I0(n1701), .I1(n1730), .CO(n29144));
    SB_LUT4 add_21_32_lut (.I0(n19), .I1(bit_ctr[30]), .I2(GND_net), .I3(n27907), 
            .O(n40191)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n43087), 
            .I3(n29357), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n29142), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_3 (.CI(n29357), .I0(n2909), .I1(n43087), .CO(n29358));
    SB_CARRY mod_5_add_1205_10 (.CI(n29142), .I0(n1702), .I1(n1730), .CO(n29143));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n43087), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n43087), 
            .CO(n29357));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n29141), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n29356), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n29141), .I0(n1703), .I1(n1730), .CO(n29142));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n29140), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_26 (.CI(n28094), .I0(timer[24]), .I1(n1[24]), 
            .CO(n28095));
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_513[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n28093), .O(n30_adj_4202)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n29355), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n29355), .I0(n2787), .I1(n2819), .CO(n29356));
    SB_CARRY mod_5_add_1205_8 (.CI(n29140), .I0(n1704), .I1(n1730), .CO(n29141));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n29139), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_32 (.CI(n27907), .I0(bit_ctr[30]), .I1(GND_net), .CO(n27908));
    SB_LUT4 add_21_31_lut (.I0(n19), .I1(bit_ctr[29]), .I2(GND_net), .I3(n27906), 
            .O(n40190)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1205_7 (.CI(n29139), .I0(n1705), .I1(n1730), .CO(n29140));
    SB_CARRY sub_14_add_2_25 (.CI(n28093), .I0(timer[23]), .I1(n1[23]), 
            .CO(n28094));
    SB_CARRY add_21_31 (.CI(n27906), .I0(bit_ctr[29]), .I1(GND_net), .CO(n27907));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n29354), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n29354), .I0(n2788), .I1(n2819), .CO(n29355));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n29138), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_30_lut (.I0(n19), .I1(bit_ctr[28]), .I2(GND_net), .I3(n27905), 
            .O(n40189)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n29353), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n29353), .I0(n2789), .I1(n2819), .CO(n29354));
    SB_CARRY mod_5_add_1205_6 (.CI(n29138), .I0(n1706), .I1(n1730), .CO(n29139));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n29352), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n29137), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_11 (.CI(n27886), .I0(bit_ctr[9]), .I1(GND_net), .CO(n27887));
    SB_CARRY mod_5_add_1205_5 (.CI(n29137), .I0(n1707), .I1(n1730), .CO(n29138));
    SB_CARRY add_21_30 (.CI(n27905), .I0(bit_ctr[28]), .I1(GND_net), .CO(n27906));
    SB_LUT4 add_21_29_lut (.I0(n19), .I1(bit_ctr[27]), .I2(GND_net), .I3(n27904), 
            .O(n40188)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n29136), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n29352), .I0(n2790), .I1(n2819), .CO(n29353));
    SB_CARRY add_21_29 (.CI(n27904), .I0(bit_ctr[27]), .I1(GND_net), .CO(n27905));
    SB_LUT4 add_21_28_lut (.I0(n19), .I1(bit_ctr[26]), .I2(GND_net), .I3(n27903), 
            .O(n40187)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_28 (.CI(n27903), .I0(bit_ctr[26]), .I1(GND_net), .CO(n27904));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n29351), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n29351), .I0(n2791), .I1(n2819), .CO(n29352));
    SB_CARRY mod_5_add_1205_4 (.CI(n29136), .I0(n1708), .I1(n1730), .CO(n29137));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n43090), 
            .I3(n29135), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_27_lut (.I0(n19), .I1(bit_ctr[25]), .I2(GND_net), .I3(n27902), 
            .O(n40186)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1205_3 (.CI(n29135), .I0(n1709), .I1(n43090), .CO(n29136));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n43090), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n29350), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n43090), 
            .CO(n29135));
    SB_LUT4 add_21_3_lut (.I0(n19), .I1(bit_ctr[1]), .I2(GND_net), .I3(n27878), 
            .O(n40193)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_27 (.CI(n27902), .I0(bit_ctr[25]), .I1(GND_net), .CO(n27903));
    SB_LUT4 add_21_26_lut (.I0(n19), .I1(bit_ctr[24]), .I2(GND_net), .I3(n27901), 
            .O(n40185)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_24_lut (.I0(one_wire_N_513[13]), .I1(timer[22]), 
            .I2(n1[22]), .I3(n28092), .O(n24_adj_4197)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1942_20 (.CI(n29350), .I0(n2792), .I1(n2819), .CO(n29351));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n29349), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n29134), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n29133), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_10_lut (.I0(n11), .I1(bit_ctr[8]), .I2(GND_net), .I3(n27885), 
            .O(n40171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_24 (.CI(n28092), .I0(timer[22]), .I1(n1[22]), 
            .CO(n28093));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_513[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n28091), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_10 (.CI(n27885), .I0(bit_ctr[8]), .I1(GND_net), .CO(n27886));
    SB_CARRY sub_14_add_2_23 (.CI(n28091), .I0(timer[21]), .I1(n1[21]), 
            .CO(n28092));
    SB_CARRY mod_5_add_1942_19 (.CI(n29349), .I0(n2793), .I1(n2819), .CO(n29350));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n29348), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n29348), .I0(n2794), .I1(n2819), .CO(n29349));
    SB_CARRY mod_5_add_1138_13 (.CI(n29133), .I0(n1599), .I1(n1631), .CO(n29134));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n29347), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n29132), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n29132), .I0(n1600), .I1(n1631), .CO(n29133));
    SB_CARRY mod_5_add_1942_17 (.CI(n29347), .I0(n2795), .I1(n2819), .CO(n29348));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n29346), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n29131), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n29131), .I0(n1601), .I1(n1631), .CO(n29132));
    SB_CARRY mod_5_add_1942_16 (.CI(n29346), .I0(n2796), .I1(n2819), .CO(n29347));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n29130), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n29130), .I0(n1602), .I1(n1631), .CO(n29131));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n29345), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n29129), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n29345), .I0(n2797), .I1(n2819), .CO(n29346));
    SB_CARRY mod_5_add_1138_9 (.CI(n29129), .I0(n1603), .I1(n1631), .CO(n29130));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n29344), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n29128), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n29344), .I0(n2798), .I1(n2819), .CO(n29345));
    SB_CARRY mod_5_add_1138_8 (.CI(n29128), .I0(n1604), .I1(n1631), .CO(n29129));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n29343), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n29127), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n29343), .I0(n2799), .I1(n2819), .CO(n29344));
    SB_CARRY mod_5_add_1138_7 (.CI(n29127), .I0(n1605), .I1(n1631), .CO(n29128));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n29342), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n29126), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n29126), .I0(n1606), .I1(n1631), .CO(n29127));
    SB_CARRY add_21_26 (.CI(n27901), .I0(bit_ctr[24]), .I1(GND_net), .CO(n27902));
    SB_CARRY mod_5_add_1942_12 (.CI(n29342), .I0(n2800), .I1(n2819), .CO(n29343));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n29125), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_513[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n28090), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n29341), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_22 (.CI(n28090), .I0(timer[20]), .I1(n1[20]), 
            .CO(n28091));
    SB_CARRY mod_5_add_1138_5 (.CI(n29125), .I0(n1607), .I1(n1631), .CO(n29126));
    SB_CARRY mod_5_add_1942_11 (.CI(n29341), .I0(n2801), .I1(n2819), .CO(n29342));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n29340), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n29124), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n29124), .I0(n1608), .I1(n1631), .CO(n29125));
    SB_CARRY mod_5_add_1942_10 (.CI(n29340), .I0(n2802), .I1(n2819), .CO(n29341));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n43092), 
            .I3(n29123), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n29123), .I0(n1609), .I1(n43092), .CO(n29124));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n28089), .O(one_wire_N_513[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF timer_1177__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n43092), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n29339), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n43092), 
            .CO(n29123));
    SB_CARRY mod_5_add_1942_9 (.CI(n29339), .I0(n2803), .I1(n2819), .CO(n29340));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n29122), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n29338), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n29121), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n29338), .I0(n2804), .I1(n2819), .CO(n29339));
    SB_CARRY mod_5_add_1071_12 (.CI(n29121), .I0(n1500), .I1(n1532), .CO(n29122));
    SB_LUT4 add_21_25_lut (.I0(n19), .I1(bit_ctr[23]), .I2(GND_net), .I3(n27900), 
            .O(n40184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n29337), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_25 (.CI(n27900), .I0(bit_ctr[23]), .I1(GND_net), .CO(n27901));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n29120), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n29337), .I0(n2805), .I1(n2819), .CO(n29338));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n29336), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n29120), .I0(n1501), .I1(n1532), .CO(n29121));
    SB_CARRY sub_14_add_2_21 (.CI(n28089), .I0(timer[19]), .I1(n1[19]), 
            .CO(n28090));
    SB_LUT4 add_21_9_lut (.I0(n19), .I1(bit_ctr[7]), .I2(GND_net), .I3(n27884), 
            .O(n40199)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_6 (.CI(n29336), .I0(n2806), .I1(n2819), .CO(n29337));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n29119), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n29335), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n29335), .I0(n2807), .I1(n2819), .CO(n29336));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n29334), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n29119), .I0(n1502), .I1(n1532), .CO(n29120));
    SB_DFF timer_1177__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1177__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF start_103 (.Q(start), .C(clk32MHz), .D(n33387));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n16831));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n17017));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n29118), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n29334), .I0(n2808), .I1(n2819), .CO(n29335));
    SB_CARRY mod_5_add_1071_9 (.CI(n29118), .I0(n1503), .I1(n1532), .CO(n29119));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n28088), .O(one_wire_N_513[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n28088), .I0(timer[18]), .I1(n1[18]), 
            .CO(n28089));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_513[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n28087), .O(n27_adj_4198)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n28087), .I0(timer[17]), .I1(n1[17]), 
            .CO(n28088));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n43091), 
            .I3(n29333), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n29117), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n29117), .I0(n1504), .I1(n1532), .CO(n29118));
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n28086), .O(one_wire_N_513[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_3 (.CI(n29333), .I0(n2809), .I1(n43091), .CO(n29334));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n29116), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n43091), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_7 (.CI(n29116), .I0(n1505), .I1(n1532), .CO(n29117));
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n43091), 
            .CO(n29333));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n29115), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n29332), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n29115), .I0(n1506), .I1(n1532), .CO(n29116));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n29114), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n29114), .I0(n1507), .I1(n1532), .CO(n29115));
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n29331), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n29113), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n29113), .I0(n1508), .I1(n1532), .CO(n29114));
    SB_CARRY mod_5_add_1875_24 (.CI(n29331), .I0(n2688), .I1(n2720), .CO(n29332));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n43093), 
            .I3(n29112), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_3 (.CI(n29112), .I0(n1509), .I1(n43093), .CO(n29113));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n29330), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n29330), .I0(n2689), .I1(n2720), .CO(n29331));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n43093), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n29329), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n43093), 
            .CO(n29112));
    SB_CARRY mod_5_add_1875_22 (.CI(n29329), .I0(n2690), .I1(n2720), .CO(n29330));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n29328), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n29328), .I0(n2691), .I1(n2720), .CO(n29329));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n29327), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_18 (.CI(n28086), .I0(timer[16]), .I1(n1[16]), 
            .CO(n28087));
    SB_CARRY mod_5_add_1875_20 (.CI(n29327), .I0(n2692), .I1(n2720), .CO(n29328));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n29326), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n29326), .I0(n2693), .I1(n2720), .CO(n29327));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n29325), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n29325), .I0(n2694), .I1(n2720), .CO(n29326));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n29324), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n29324), .I0(n2695), .I1(n2720), .CO(n29325));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n29323), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_3 (.CI(n27878), .I0(bit_ctr[1]), .I1(GND_net), .CO(n27879));
    SB_CARRY mod_5_add_1875_16 (.CI(n29323), .I0(n2696), .I1(n2720), .CO(n29324));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n29322), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n28085), .O(one_wire_N_513[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_15 (.CI(n29322), .I0(n2697), .I1(n2720), .CO(n29323));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n29321), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_17 (.CI(n28085), .I0(timer[15]), .I1(n1[15]), 
            .CO(n28086));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n28084), .O(one_wire_N_513[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_16 (.CI(n28084), .I0(timer[14]), .I1(n1[14]), 
            .CO(n28085));
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n28083), .O(one_wire_N_513[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_14 (.CI(n29321), .I0(n2698), .I1(n2720), .CO(n29322));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n29320), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n29320), .I0(n2699), .I1(n2720), .CO(n29321));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n29319), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n29319), .I0(n2700), .I1(n2720), .CO(n29320));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n29318), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n29318), .I0(n2701), .I1(n2720), .CO(n29319));
    SB_CARRY sub_14_add_2_15 (.CI(n28083), .I0(timer[13]), .I1(n1[13]), 
            .CO(n28084));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n29317), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n29317), .I0(n2702), .I1(n2720), .CO(n29318));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n29316), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n29316), .I0(n2703), .I1(n2720), .CO(n29317));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n29315), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n29315), .I0(n2704), .I1(n2720), .CO(n29316));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n29314), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n29314), .I0(n2705), .I1(n2720), .CO(n29315));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n29313), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n29313), .I0(n2706), .I1(n2720), .CO(n29314));
    SB_CARRY add_21_9 (.CI(n27884), .I0(bit_ctr[7]), .I1(GND_net), .CO(n27885));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n29312), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_5 (.CI(n29312), .I0(n2707), .I1(n2720), .CO(n29313));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n29311), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_24_lut (.I0(n19), .I1(bit_ctr[22]), .I2(GND_net), .I3(n27899), 
            .O(n40183)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1875_4 (.CI(n29311), .I0(n2708), .I1(n2720), .CO(n29312));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n43094), 
            .I3(n29310), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n29310), .I0(n2709), .I1(n43094), .CO(n29311));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n43094), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n43094), 
            .CO(n29310));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n29309), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n29308), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n29308), .I0(n2589), .I1(n2621), .CO(n29309));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n29307), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n29307), .I0(n2590), .I1(n2621), .CO(n29308));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n29306), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n29306), .I0(n2591), .I1(n2621), .CO(n29307));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n29305), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n29305), .I0(n2592), .I1(n2621), .CO(n29306));
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n28082), .O(one_wire_N_513[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n29304), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n29304), .I0(n2593), .I1(n2621), .CO(n29305));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n29303), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n29303), .I0(n2594), .I1(n2621), .CO(n29304));
    SB_LUT4 add_21_2_lut (.I0(n19), .I1(bit_ctr[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n40177)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_8_lut (.I0(n19), .I1(bit_ctr[6]), .I2(GND_net), .I3(n27883), 
            .O(n40198)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n29302), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_14 (.CI(n28082), .I0(timer[12]), .I1(n1[12]), 
            .CO(n28083));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n28081), .O(\one_wire_N_513[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n28312), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n28311), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n28311), .I0(n906), .I1(VCC_net), .CO(n28312));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n35441), .I2(VCC_net), 
            .I3(n28310), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n28081), .I0(timer[11]), .I1(n1[11]), 
            .CO(n28082));
    SB_CARRY mod_5_add_669_5 (.CI(n28310), .I0(n35441), .I1(VCC_net), 
            .CO(n28311));
    SB_CARRY add_21_24 (.CI(n27899), .I0(bit_ctr[22]), .I1(GND_net), .CO(n27900));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n16683), .I2(VCC_net), 
            .I3(n28309), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n28309), .I0(n16683), .I1(VCC_net), 
            .CO(n28310));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n14144), .I2(GND_net), 
            .I3(n28308), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n28308), .I0(n14144), .I1(GND_net), 
            .CO(n28309));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n28308));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4228), .I1(n4_adj_4228), .I2(n1037), 
            .I3(n28307), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n28306), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n28306), .I0(n1005), .I1(n1037), .CO(n28307));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n28305), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n29302), .I0(n2595), .I1(n2621), .CO(n29303));
    SB_CARRY mod_5_add_736_6 (.CI(n28305), .I0(n1006), .I1(n1037), .CO(n28306));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n29301), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n28304), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n28304), .I0(n1007), .I1(n1037), .CO(n28305));
    SB_CARRY add_21_8 (.CI(n27883), .I0(bit_ctr[6]), .I1(GND_net), .CO(n27884));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n28303), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n28303), .I0(n1008), .I1(n1037), .CO(n28304));
    SB_CARRY mod_5_add_1808_16 (.CI(n29301), .I0(n2596), .I1(n2621), .CO(n29302));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n43096), 
            .I3(n28302), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n28302), .I0(n1009), .I1(n43096), .CO(n28303));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n29300), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n43096), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_15 (.CI(n29300), .I0(n2597), .I1(n2621), .CO(n29301));
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n43096), 
            .CO(n28302));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n28080), .O(\one_wire_N_513[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n29299), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n29299), .I0(n2598), .I1(n2621), .CO(n29300));
    SB_CARRY sub_14_add_2_12 (.CI(n28080), .I0(timer[10]), .I1(n1[10]), 
            .CO(n28081));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n29298), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_23_lut (.I0(n19), .I1(bit_ctr[21]), .I2(GND_net), .I3(n27898), 
            .O(n40182)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1808_13 (.CI(n29298), .I0(n2599), .I1(n2621), .CO(n29299));
    SB_CARRY add_21_23 (.CI(n27898), .I0(bit_ctr[21]), .I1(GND_net), .CO(n27899));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n29297), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n29297), .I0(n2600), .I1(n2621), .CO(n29298));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n29296), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n29296), .I0(n2601), .I1(n2621), .CO(n29297));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n29295), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n29295), .I0(n2602), .I1(n2621), .CO(n29296));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n28079), .O(\one_wire_N_513[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n29294), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n29294), .I0(n2603), .I1(n2621), .CO(n29295));
    SB_LUT4 i3_4_lut_4_lut (.I0(n35321), .I1(n14146), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n14146), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n35321), .O(n35441));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n29293), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n29293), .I0(n2604), .I1(n2621), .CO(n29294));
    SB_CARRY sub_14_add_2_11 (.CI(n28079), .I0(timer[9]), .I1(n1[9]), 
            .CO(n28080));
    SB_LUT4 add_21_22_lut (.I0(n19), .I1(bit_ctr[20]), .I2(GND_net), .I3(n27897), 
            .O(n40178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n29292), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n28078), .O(\one_wire_N_513[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_7 (.CI(n29292), .I0(n2605), .I1(n2621), .CO(n29293));
    SB_CARRY sub_14_add_2_10 (.CI(n28078), .I0(timer[8]), .I1(n1[8]), 
            .CO(n28079));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n27878));
    SB_CARRY add_21_22 (.CI(n27897), .I0(bit_ctr[20]), .I1(GND_net), .CO(n27898));
    SB_LUT4 add_21_21_lut (.I0(n19), .I1(bit_ctr[19]), .I2(GND_net), .I3(n27896), 
            .O(n40174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n29291), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n28077), .O(\one_wire_N_513[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_6 (.CI(n29291), .I0(n2606), .I1(n2621), .CO(n29292));
    SB_CARRY sub_14_add_2_9 (.CI(n28077), .I0(timer[7]), .I1(n1[7]), .CO(n28078));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n29290), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n28076), .O(\one_wire_N_513[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n28076), .I0(timer[6]), .I1(n1[6]), .CO(n28077));
    SB_CARRY add_21_21 (.CI(n27896), .I0(bit_ctr[19]), .I1(GND_net), .CO(n27897));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n28075), .O(\one_wire_N_513[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n28075), .I0(timer[5]), .I1(n1[5]), .CO(n28076));
    SB_CARRY mod_5_add_1808_5 (.CI(n29290), .I0(n2607), .I1(n2621), .CO(n29291));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n29289), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n28074), .O(one_wire_N_513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_20_lut (.I0(n19), .I1(bit_ctr[18]), .I2(GND_net), .I3(n27895), 
            .O(n40173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_6 (.CI(n28074), .I0(timer[4]), .I1(n1[4]), .CO(n28075));
    SB_CARRY mod_5_add_1808_4 (.CI(n29289), .I0(n2608), .I1(n2621), .CO(n29290));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n28073), .O(one_wire_N_513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n43095), 
            .I3(n29288), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i34080_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n24913), .I2(n35437), 
            .I3(bit_ctr[28]), .O(n35321));
    defparam i34080_3_lut_4_lut.LUT_INIT = 16'h9666;
    SB_CARRY add_21_20 (.CI(n27895), .I0(bit_ctr[18]), .I1(GND_net), .CO(n27896));
    SB_CARRY sub_14_add_2_5 (.CI(n28073), .I0(timer[3]), .I1(n1[3]), .CO(n28074));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n28072), .O(one_wire_N_513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_3 (.CI(n29288), .I0(n2609), .I1(n43095), .CO(n29289));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n43095), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_4 (.CI(n28072), .I0(timer[2]), .I1(n1[2]), .CO(n28073));
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4239), .I1(timer[1]), .I2(n1[1]), 
            .I3(n28071), .O(n30241)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_3 (.CI(n28071), .I0(timer[1]), .I1(n1[1]), .CO(n28072));
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n43095), 
            .CO(n29288));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n29287), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n29286), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n29286), .I0(n2490), .I1(n2522), .CO(n29287));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28250), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28249), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n28249), .I0(n1104), .I1(n1136), .CO(n28250));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28248), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n28248), .I0(n1105), .I1(n1136), .CO(n28249));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n29285), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28247), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n28247), .I0(n1106), .I1(n1136), .CO(n28248));
    SB_CARRY mod_5_add_1741_21 (.CI(n29285), .I0(n2491), .I1(n2522), .CO(n29286));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_513[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_adj_4239)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28246), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n29284), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i20037_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n24695));   // verilog/neopixel.v(22[26:36])
    defparam i20037_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i20049_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n24707));
    defparam i20049_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1500 (.I0(n1405), .I1(n24707), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4240));
    defparam i6_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1501 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4241));
    defparam i7_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1502 (.I0(n17_adj_4241), .I1(n1408), .I2(n16_adj_4240), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1502.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1503 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4242));
    defparam i14_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1504 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4243));
    defparam i18_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1505 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42));
    defparam i16_4_lut_adj_1505.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1506 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4244));
    defparam i17_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1507 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4245));
    defparam i15_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_4246));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4242), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4247));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut_adj_1508 (.I0(n41_adj_4245), .I1(n43_adj_4244), .I2(n42), 
            .I3(n44_adj_4243), .O(n50));
    defparam i24_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4248));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37_adj_4248), .I1(n50), .I2(n46_adj_4247), 
            .I3(n38_adj_4246), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36315_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43077));
    defparam i36315_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1509 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4249));
    defparam i1_2_lut_adj_1509.LUT_INIT = 16'heeee;
    SB_LUT4 i20031_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n24689));
    defparam i20031_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1510 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_4249), 
            .O(n30_adj_4250));
    defparam i13_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1511 (.I0(n2098), .I1(n24689), .I2(n2094), .I3(n2099), 
            .O(n28_adj_4251));
    defparam i11_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1512 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4252));
    defparam i12_4_lut_adj_1512.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1513 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4253));
    defparam i10_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1514 (.I0(n27_adj_4253), .I1(n29_adj_4252), .I2(n28_adj_4251), 
            .I3(n30_adj_4250), .O(n2126));
    defparam i16_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_LUT4 i36316_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43078));
    defparam i36316_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1515 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4254));
    defparam i10_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1516 (.I0(n2203), .I1(n28_adj_4254), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4255));
    defparam i14_4_lut_adj_1516.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1517 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4256));
    defparam i12_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i36333_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43095));
    defparam i36333_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13_4_lut_adj_1518 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4257));
    defparam i13_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1519 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4258));
    defparam i11_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1520 (.I0(n29_adj_4258), .I1(n31_adj_4257), .I2(n30_adj_4256), 
            .I3(n32_adj_4255), .O(n2225));
    defparam i17_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut_adj_1521 (.I0(n3084), .I1(n3085), .I2(n3097), .I3(n3096), 
            .O(n42_adj_4259));
    defparam i15_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1522 (.I0(n3108), .I1(n3101), .I2(n3104), .I3(n3094), 
            .O(n46_adj_4260));
    defparam i19_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1523 (.I0(n3100), .I1(n3089), .I2(n3093), .I3(n3103), 
            .O(n44_adj_4261));
    defparam i17_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1524 (.I0(n3099), .I1(n3092), .I2(n3098), .I3(n3083), 
            .O(n45_adj_4262));
    defparam i18_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1525 (.I0(n3090), .I1(n3087), .I2(n3095), .I3(n3091), 
            .O(n43_adj_4263));
    defparam i16_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(n3106), .I1(n3086), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_4264));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i21_4_lut_adj_1526 (.I0(n3102), .I1(n42_adj_4259), .I2(n3088), 
            .I3(n3107), .O(n48_adj_4265));
    defparam i21_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1527 (.I0(n43_adj_4263), .I1(n45_adj_4262), .I2(n44_adj_4261), 
            .I3(n46_adj_4260), .O(n52));
    defparam i25_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_3_lut (.I0(n3105), .I1(bit_ctr[4]), .I2(n3109), .I3(GND_net), 
            .O(n39_adj_4266));
    defparam i12_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i26_4_lut_adj_1528 (.I0(n39_adj_4266), .I1(n52), .I2(n48_adj_4265), 
            .I3(n40_adj_4264), .O(n3116));
    defparam i26_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i36314_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43076));
    defparam i36314_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut_adj_1529 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4267));
    defparam i3_2_lut_adj_1529.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1530 (.I0(bit_ctr[12]), .I1(n22_adj_4267), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4268));
    defparam i11_4_lut_adj_1530.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1531 (.I0(n2294), .I1(n30_adj_4268), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4269));
    defparam i15_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1532 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4270));
    defparam i13_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1533 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4271));
    defparam i14_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1534 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4272));
    defparam i12_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1535 (.I0(n31_adj_4272), .I1(n33_adj_4271), .I2(n32_adj_4270), 
            .I3(n34_adj_4269), .O(n2324));
    defparam i18_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36334_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43096));
    defparam i36334_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36299_2_lut (.I0(n31213), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i36299_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i36313_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43075));
    defparam i36313_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36301_2_lut (.I0(n31213), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i36301_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n31213), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31377_3_lut (.I0(n905), .I1(n906), .I2(n35441), .I3(GND_net), 
            .O(n38080));
    defparam i31377_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n38080), .I2(n16683), .I3(n14144), 
            .O(n31213));
    defparam i4_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n31213), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n14144), .I1(n971[27]), .I2(n31213), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31379_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n38082));
    defparam i31379_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1536 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_4273));
    defparam i2_3_lut_adj_1536.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut_adj_1537 (.I0(n31213), .I1(n6_adj_4273), .I2(n1005), 
            .I3(n38082), .O(n1037));
    defparam i3_4_lut_adj_1537.LUT_INIT = 16'hfdfc;
    SB_LUT4 i36297_2_lut (.I0(n31213), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4228));   // verilog/neopixel.v(22[26:36])
    defparam i36297_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1538 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n14144));
    defparam i1_2_lut_adj_1538.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i19996_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i19996_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut_adj_1539 (.I0(n708), .I1(n24695), .I2(n35339), .I3(n608), 
            .O(n35437));
    defparam i2_4_lut_adj_1539.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_adj_1540 (.I0(bit_ctr[28]), .I1(n35437), .I2(GND_net), 
            .I3(GND_net), .O(n14146));
    defparam i1_2_lut_adj_1540.LUT_INIT = 16'h9999;
    SB_LUT4 i31286_3_lut (.I0(n35437), .I1(n708), .I2(n35339), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam i31286_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1541 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4274));
    defparam i14_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1542 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4275));
    defparam i3_3_lut_adj_1542.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1543 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4276));
    defparam i12_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1544 (.I0(n25_adj_4275), .I1(n36_adj_4274), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4277));
    defparam i18_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1545 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4278));
    defparam i16_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4276), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4279));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1546 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4280));
    defparam i15_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1547 (.I0(n37_adj_4280), .I1(n39_adj_4279), .I2(n38_adj_4278), 
            .I3(n40_adj_4277), .O(n2621));
    defparam i21_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i36332_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43094));
    defparam i36332_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36331_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43093));
    defparam i36331_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4281));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1548 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4282));
    defparam i15_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i20165_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n24823));
    defparam i20165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1549 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n24823), 
            .O(n36_adj_4283));
    defparam i13_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1550 (.I0(n2700), .I1(n38_adj_4282), .I2(n28_adj_4281), 
            .I3(n2705), .O(n42_adj_4284));
    defparam i19_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1551 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4285));
    defparam i17_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1552 (.I0(n2687), .I1(n36_adj_4283), .I2(n2703), 
            .I3(n2695), .O(n41_adj_4286));
    defparam i18_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1553 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4287));
    defparam i16_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1554 (.I0(n39_adj_4287), .I1(n41_adj_4286), .I2(n40_adj_4285), 
            .I3(n42_adj_4284), .O(n2720));
    defparam i22_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36329_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43091));
    defparam i36329_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1555 (.I0(n1505), .I1(bit_ctr[20]), .I2(n1509), 
            .I3(GND_net), .O(n12_adj_4288));
    defparam i1_3_lut_adj_1555.LUT_INIT = 16'heaea;
    SB_LUT4 i7_4_lut_adj_1556 (.I0(n1506), .I1(n1508), .I2(n1503), .I3(n1501), 
            .O(n18_adj_4289));
    defparam i7_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1557 (.I0(n1504), .I1(n1500), .I2(n1502), .I3(n1507), 
            .O(n19_adj_4290));
    defparam i8_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1558 (.I0(n19_adj_4290), .I1(n1499), .I2(n18_adj_4289), 
            .I3(n12_adj_4288), .O(n1532));
    defparam i10_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36330_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43092));
    defparam i36330_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1559 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4291));
    defparam i8_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1560 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4292));
    defparam i1_3_lut_adj_1560.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4293));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1561 (.I0(n13_adj_4292), .I1(n20_adj_4291), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4294));
    defparam i10_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1562 (.I0(n1601), .I1(n22_adj_4294), .I2(n18_adj_4293), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36328_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43090));
    defparam i36328_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1563 (.I0(n2791), .I1(n2805), .I2(n2801), .I3(n2806), 
            .O(n40_adj_4295));
    defparam i16_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1564 (.I0(n2796), .I1(n2787), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4296));
    defparam i14_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1565 (.I0(n2799), .I1(n2798), .I2(n2803), .I3(n2794), 
            .O(n39_adj_4297));
    defparam i15_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1566 (.I0(n2804), .I1(n2786), .I2(n2795), .I3(n2797), 
            .O(n37_adj_4298));
    defparam i13_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2793), .I1(n2802), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4299));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1567 (.I0(n2800), .I1(n2789), .I2(n2807), .I3(n2792), 
            .O(n42_adj_4300));
    defparam i18_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1568 (.I0(n37_adj_4298), .I1(n39_adj_4297), .I2(n38_adj_4296), 
            .I3(n40_adj_4295), .O(n46_adj_4301));
    defparam i22_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2790), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4302));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut (.I0(n33_adj_4302), .I1(n46_adj_4301), .I2(n42_adj_4300), 
            .I3(n34_adj_4299), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36325_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43087));
    defparam i36325_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1569 (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_4303));
    defparam i4_3_lut_adj_1569.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1570 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4304));
    defparam i8_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1571 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4305));
    defparam i7_3_lut_adj_1571.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1572 (.I0(n21_adj_4304), .I1(n17_adj_4303), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4306));
    defparam i11_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1573 (.I0(n1700), .I1(n24_adj_4306), .I2(n20_adj_4305), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28756_2_lut (.I0(one_wire_N_513[4]), .I1(n35378), .I2(GND_net), 
            .I3(GND_net), .O(n35457));
    defparam i28756_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i130_4_lut (.I0(n24733), .I1(n35483), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n103));
    defparam i130_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1574 (.I0(n35481), .I1(n35457), .I2(n4), .I3(n34616), 
            .O(n34539));
    defparam i1_4_lut_adj_1574.LUT_INIT = 16'h1505;
    SB_LUT4 i1_4_lut_adj_1575 (.I0(n15538), .I1(\state[0] ), .I2(n34539), 
            .I3(n103), .O(n16544));
    defparam i1_4_lut_adj_1575.LUT_INIT = 16'h5150;
    SB_LUT4 i96_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_576 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i96_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20155_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n24813));
    defparam i20155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut_adj_1576 (.I0(n3202), .I1(n3195), .I2(n3205), .I3(n3204), 
            .O(n20_adj_4307));
    defparam i8_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1577 (.I0(n3198), .I1(n3186), .I2(n24813), .I3(n3194), 
            .O(n19_adj_4308));
    defparam i7_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1578 (.I0(n3191), .I1(n3207), .I2(n3187), .I3(n3203), 
            .O(n21_adj_4309));
    defparam i9_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(n21_adj_4309), .I1(n3189), .I2(n19_adj_4308), 
            .I3(n20_adj_4307), .O(n18_adj_4310));
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1580 (.I0(n3190), .I1(n3185), .I2(n3192), .I3(n18_adj_4310), 
            .O(n30_adj_4311));
    defparam i13_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1581 (.I0(n3183), .I1(n3188), .I2(n3208), .I3(n3200), 
            .O(n28_adj_4312));
    defparam i11_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1582 (.I0(n3182), .I1(n3196), .I2(n3197), .I3(n3199), 
            .O(n29_adj_4313));
    defparam i12_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1583 (.I0(n3193), .I1(n3184), .I2(n3206), .I3(n3201), 
            .O(n27_adj_4314));
    defparam i10_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1584 (.I0(n27_adj_4314), .I1(n29_adj_4313), .I2(n28_adj_4312), 
            .I3(n30_adj_4311), .O(n24877));
    defparam i16_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i20075_3_lut (.I0(\one_wire_N_513[9] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[10] ), .I3(GND_net), .O(n24733));
    defparam i20075_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i234_2_lut (.I0(n24853), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1166));   // verilog/neopixel.v(103[9] 111[12])
    defparam i234_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1585 (.I0(n4_adj_4315), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(n1166), .O(n16754));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1585.LUT_INIT = 16'h0a3a;
    SB_LUT4 i1_4_lut_adj_1586 (.I0(\state[0] ), .I1(n4_adj_4315), .I2(n1166), 
            .I3(\state[1] ), .O(n16530));
    defparam i1_4_lut_adj_1586.LUT_INIT = 16'hafcc;
    SB_LUT4 color_bit_I_0_i2_3_lut (.I0(\color[2] ), .I1(\color[3] ), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n2_adj_4316));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1587 (.I0(\color[4] ), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4317));
    defparam i1_2_lut_adj_1587.LUT_INIT = 16'h2222;
    SB_LUT4 i34329_4_lut (.I0(\color[1] ), .I1(n2_adj_4316), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n41093));   // verilog/neopixel.v(22[26:36])
    defparam i34329_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 color_bit_I_0_i7_4_lut (.I0(n41093), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(n4_adj_4317), .O(n7_adj_4318));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i7_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i31333_4_lut (.I0(\state_3__N_362[1] ), .I1(n3209), .I2(bit_ctr[3]), 
            .I3(n24877), .O(n38035));
    defparam i31333_4_lut.LUT_INIT = 16'hbeee;
    SB_LUT4 i3_4_lut_adj_1588 (.I0(n38035), .I1(n7_adj_4318), .I2(bit_ctr[3]), 
            .I3(n24877), .O(state_3__N_362[0]));
    defparam i3_4_lut_adj_1588.LUT_INIT = 16'h4004;
    SB_LUT4 i1_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n24907), .I3(GND_net), .O(n4_adj_4315));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i20195_2_lut_4_lut (.I0(\one_wire_N_513[9] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[10] ), .I3(n15538), .O(n24853));
    defparam i20195_2_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 i28782_2_lut_3_lut (.I0(n35481), .I1(one_wire_N_513[4]), .I2(n35378), 
            .I3(GND_net), .O(n35483));
    defparam i28782_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i20253_2_lut_3_lut (.I0(n24695), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n24913));   // verilog/neopixel.v(22[26:36])
    defparam i20253_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i34084_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n35437), .I2(bit_ctr[27]), 
            .I3(n838), .O(n16683));
    defparam i34084_3_lut_4_lut.LUT_INIT = 16'h6696;
    SB_LUT4 i28644_2_lut_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n24695), .I2(n608), 
            .I3(bit_ctr[28]), .O(n35339));
    defparam i28644_2_lut_3_lut_4_lut.LUT_INIT = 16'h5600;
    SB_LUT4 i2765_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n35437), .I2(bit_ctr[27]), 
            .I3(n35321), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i2765_2_lut_3_lut_4_lut.LUT_INIT = 16'hff60;
    SB_LUT4 i2_3_lut_4_lut (.I0(n24907), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(\state[1] ), .O(n35798));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i23_3_lut_4_lut (.I0(n24891), .I1(one_wire_N_513[4]), .I2(n30086), 
            .I3(\state[0] ), .O(n35367));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf0ee;
    SB_LUT4 mux_662_Mux_0_i3_3_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_662_Mux_0_i3_3_lut_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i1_3_lut_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n34664));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(n15335), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(n4), .O(n15466));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf3f7;
    SB_LUT4 i1_2_lut_4_lut (.I0(n30086), .I1(n15335), .I2(\neo_pixel_transmitter.done ), 
            .I3(start), .O(n1163));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff1f;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(n24695), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hd622;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36326_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43088));
    defparam i36326_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_in_frame[1] , \data_in_frame[17] , clk32MHz, \data_in_frame[2] , 
            GND_net, \data_in_frame[5] , \data_in_frame[3] , rx_data, 
            \data_out_frame[13] , \data_out_frame[15] , \data_in_frame[6] , 
            \data_out_frame[19] , \data_out_frame[18] , \data_out_frame[16] , 
            \data_out_frame[20] , n17581, setpoint, n17582, n17583, 
            n17584, n17585, n17586, n17587, n17574, n17575, n17576, 
            n17577, n17578, \data_out_frame[17] , n17595, n17596, 
            n17593, n17594, n17591, n17592, \data_out_frame[12] , 
            n17588, n17589, n17590, n17579, n17580, n17495, PWMLimit, 
            \data_out_frame[14] , n17496, n17497, n17498, n17499, 
            n17500, n17501, n17487, n17488, n17489, n17490, n17491, 
            n17492, \data_in_frame[10] , n43272, \data_in_frame[19] , 
            \data_in_frame[18] , n17493, n17494, n17479, n17480, n17481, 
            n17482, n17483, n17484, n17485, n17486, \data_out_frame[8] , 
            \data_in_frame[9] , \data_out_frame[7] , \data_in_frame[7] , 
            \data_out_frame[11] , \data_out_frame[6] , \data_out_frame[5] , 
            \data_out_frame[9] , \data_out_frame[10] , n17303, control_mode, 
            n17302, n17301, n17300, n17299, n17298, n17297, n17295, 
            n17294, n17293, n17292, n17291, n17290, n17289, n17288, 
            n17287, n17286, n17285, n17284, n17283, n17282, n17281, 
            n17280, n17279, n17278, rx_data_ready, n17277, n17276, 
            n17275, n17274, \FRAME_MATCHER.state[0] , n36839, n4300, 
            n17273, n17272, n17271, n17270, \data_in_frame[8] , n17269, 
            n17268, \FRAME_MATCHER.state[3] , n17267, n17266, n17265, 
            n17264, n17263, n17262, n17261, n17260, n17259, n17258, 
            n17257, n17256, n17255, n34657, n18962, n63, n17254, 
            n17253, n17252, n17251, n17250, n17249, n17248, n17247, 
            n17246, n17245, n17244, n17243, n17242, n17241, n17240, 
            n17239, n17238, n17237, n17236, n17235, n17234, n17233, 
            n17232, n17231, n17230, n17229, n17228, n17227, n17226, 
            n17225, n17224, n17223, n17222, n17221, n17220, n17219, 
            n17218, n17217, n17216, n17215, n17214, n17213, n17212, 
            n17211, n17210, n17209, n17208, n17207, n17206, n17205, 
            n17204, n17203, n17202, n17201, n17200, n17199, n17198, 
            n17197, n17196, n17195, n17194, n17193, n17192, n17191, 
            n17190, n17189, n17188, n17187, n17186, n17185, n17184, 
            n17183, n17182, n17181, n17180, n17179, n17178, n17177, 
            n17176, n17175, n17174, n17173, n17172, n17171, n17170, 
            n17169, n17165, n17164, \data_in[3] , n17163, n17162, 
            n17161, n17160, n17159, n17158, n17157, n17155, \data_in[2][6] , 
            n17154, \data_in[2][5] , n17153, \data_in[2][4] , \data_in[2][3] , 
            n17151, \data_in[2][2] , \data_in[2][1] , n17149, \data_in[2][0] , 
            n17147, \data_in[1][6] , n13195, \data_in[0] , n17146, 
            \data_in[1][5] , n737, \data_in[1][3] , \data_in[0][5] , 
            \data_in[1][2] , \data_in[0][1] , n17145, \data_in[1][4] , 
            n17144, n17143, \data_in[0][0] , \data_in[1][1] , \data_in[0][4] , 
            \data_in[0][3] , \data_in[0][6] , \data_in[1][0] , n17142, 
            n17141, n17139, n17138, \FRAME_MATCHER.i_31__N_2390 , n2855, 
            n10283, n17137, n17136, n17135, \FRAME_MATCHER.i_31__N_2386 , 
            n122, n17134, n17133, \Ki[7] , n17132, \Ki[6] , n17131, 
            \Ki[5] , n17130, \Ki[4] , n17129, \Ki[3] , n8849, n17128, 
            \Ki[2] , n17127, \Ki[1] , n17126, \Kp[7] , n17125, \Kp[6] , 
            n17124, \Kp[5] , n17123, \Kp[4] , n17122, \Kp[3] , n17121, 
            \Kp[2] , n17120, \Kp[1] , n17119, gearBoxRatio, n17118, 
            n17117, n17116, n4, \FRAME_MATCHER.state_31__N_2426[2] , 
            n7, n17115, n17114, n17113, n17112, n17111, n17110, 
            n17109, n17108, n17107, n17106, n17105, n17104, n17103, 
            n17102, n17101, n17100, n17099, n17098, n17097, n17096, 
            IntegralLimit, n17095, n17094, n17093, n17092, n17091, 
            n17090, n17089, n17088, n17087, n17086, n17085, n17084, 
            n17083, n17082, n17081, n17080, n17079, n17078, n17077, 
            n17076, n17075, n17074, n36885, n4299, n4298, n4309, 
            n4308, n4307, n4311, LED_c, n4310, n4313, n4312, n4315, 
            n4314, n16832, n16986, n33975, n16967, n16965, n16964, 
            n16963, \Ki[0] , n16962, \Kp[0] , n16961, n4292, n4297, 
            n4296, n4295, n4294, n4293, n4306, n4305, n4304, n4303, 
            n4302, n4301, n5, n318, \r_Clock_Count[3] , n16918, 
            r_Bit_Index, n16915, n16911, \r_Clock_Count[1] , n16890, 
            \r_Clock_Count[8] , n16893, \r_Clock_Count[7] , n16905, 
            n16899, \r_Clock_Count[5] , n17029, n17566, r_SM_Main, 
            n26602, n320, VCC_net, n4613, n26612, n16641, n16772, 
            tx_o, tx_enable, n313, n314, n16981, n16979, n316, 
            n3, n29, n16872, \r_Clock_Count[6] , n16869, \r_Clock_Count[7]_adj_3 , 
            n16881, \r_Clock_Count[3]_adj_4 , n16887, \r_Clock_Count[1]_adj_5 , 
            n17005, r_Bit_Index_adj_13, n17002, n17550, r_Rx_Data, 
            PIN_13_N_105, n219, n220, n30, n223, n3_adj_9, n225, 
            n15459, n4_adj_10, n16746, n16635, n17012, n17011, n17010, 
            n17009, n17008, n17007, n17006, n4591, n24014, n4_adj_11, 
            n4_adj_12, n15454) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[17] ;
    input clk32MHz;
    output [7:0]\data_in_frame[2] ;
    input GND_net;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]rx_data;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[20] ;
    input n17581;
    output [23:0]setpoint;
    input n17582;
    input n17583;
    input n17584;
    input n17585;
    input n17586;
    input n17587;
    input n17574;
    input n17575;
    input n17576;
    input n17577;
    input n17578;
    output [7:0]\data_out_frame[17] ;
    input n17595;
    input n17596;
    input n17593;
    input n17594;
    input n17591;
    input n17592;
    output [7:0]\data_out_frame[12] ;
    input n17588;
    input n17589;
    input n17590;
    input n17579;
    input n17580;
    input n17495;
    output [23:0]PWMLimit;
    output [7:0]\data_out_frame[14] ;
    input n17496;
    input n17497;
    input n17498;
    input n17499;
    input n17500;
    input n17501;
    input n17487;
    input n17488;
    input n17489;
    input n17490;
    input n17491;
    input n17492;
    output [7:0]\data_in_frame[10] ;
    input n43272;
    output [7:0]\data_in_frame[19] ;
    output [7:0]\data_in_frame[18] ;
    input n17493;
    input n17494;
    input n17479;
    input n17480;
    input n17481;
    input n17482;
    input n17483;
    input n17484;
    input n17485;
    input n17486;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_in_frame[7] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[10] ;
    input n17303;
    output [7:0]control_mode;
    input n17302;
    input n17301;
    input n17300;
    input n17299;
    input n17298;
    input n17297;
    input n17295;
    input n17294;
    input n17293;
    input n17292;
    input n17291;
    input n17290;
    input n17289;
    input n17288;
    input n17287;
    input n17286;
    input n17285;
    input n17284;
    input n17283;
    input n17282;
    input n17281;
    input n17280;
    input n17279;
    input n17278;
    output rx_data_ready;
    input n17277;
    input n17276;
    input n17275;
    input n17274;
    output \FRAME_MATCHER.state[0] ;
    output n36839;
    output n4300;
    input n17273;
    input n17272;
    input n17271;
    input n17270;
    output [7:0]\data_in_frame[8] ;
    input n17269;
    input n17268;
    output \FRAME_MATCHER.state[3] ;
    input n17267;
    input n17266;
    input n17265;
    input n17264;
    input n17263;
    input n17262;
    input n17261;
    input n17260;
    input n17259;
    input n17258;
    input n17257;
    input n17256;
    input n17255;
    output n34657;
    output n18962;
    output n63;
    input n17254;
    input n17253;
    input n17252;
    input n17251;
    input n17250;
    input n17249;
    input n17248;
    input n17247;
    input n17246;
    input n17245;
    input n17244;
    input n17243;
    input n17242;
    input n17241;
    input n17240;
    input n17239;
    input n17238;
    input n17237;
    input n17236;
    input n17235;
    input n17234;
    input n17233;
    input n17232;
    input n17231;
    input n17230;
    input n17229;
    input n17228;
    input n17227;
    input n17226;
    input n17225;
    input n17224;
    input n17223;
    input n17222;
    input n17221;
    input n17220;
    input n17219;
    input n17218;
    input n17217;
    input n17216;
    input n17215;
    input n17214;
    input n17213;
    input n17212;
    input n17211;
    input n17210;
    input n17209;
    input n17208;
    input n17207;
    input n17206;
    input n17205;
    input n17204;
    input n17203;
    input n17202;
    input n17201;
    input n17200;
    input n17199;
    input n17198;
    input n17197;
    input n17196;
    input n17195;
    input n17194;
    input n17193;
    input n17192;
    input n17191;
    input n17190;
    input n17189;
    input n17188;
    input n17187;
    input n17186;
    input n17185;
    input n17184;
    input n17183;
    input n17182;
    input n17181;
    input n17180;
    input n17179;
    input n17178;
    input n17177;
    input n17176;
    input n17175;
    input n17174;
    input n17173;
    input n17172;
    input n17171;
    input n17170;
    input n17169;
    input n17165;
    input n17164;
    output [7:0]\data_in[3] ;
    input n17163;
    input n17162;
    input n17161;
    input n17160;
    input n17159;
    input n17158;
    input n17157;
    input n17155;
    output \data_in[2][6] ;
    input n17154;
    output \data_in[2][5] ;
    input n17153;
    output \data_in[2][4] ;
    output \data_in[2][3] ;
    input n17151;
    output \data_in[2][2] ;
    output \data_in[2][1] ;
    input n17149;
    output \data_in[2][0] ;
    input n17147;
    output \data_in[1][6] ;
    output n13195;
    output [7:0]\data_in[0] ;
    input n17146;
    output \data_in[1][5] ;
    output n737;
    output \data_in[1][3] ;
    output \data_in[0][5] ;
    output \data_in[1][2] ;
    output \data_in[0][1] ;
    input n17145;
    output \data_in[1][4] ;
    input n17144;
    input n17143;
    output \data_in[0][0] ;
    output \data_in[1][1] ;
    output \data_in[0][4] ;
    output \data_in[0][3] ;
    output \data_in[0][6] ;
    output \data_in[1][0] ;
    input n17142;
    input n17141;
    input n17139;
    input n17138;
    output \FRAME_MATCHER.i_31__N_2390 ;
    output n2855;
    output n10283;
    input n17137;
    input n17136;
    input n17135;
    output \FRAME_MATCHER.i_31__N_2386 ;
    output n122;
    input n17134;
    input n17133;
    output \Ki[7] ;
    input n17132;
    output \Ki[6] ;
    input n17131;
    output \Ki[5] ;
    input n17130;
    output \Ki[4] ;
    input n17129;
    output \Ki[3] ;
    output n8849;
    input n17128;
    output \Ki[2] ;
    input n17127;
    output \Ki[1] ;
    input n17126;
    output \Kp[7] ;
    input n17125;
    output \Kp[6] ;
    input n17124;
    output \Kp[5] ;
    input n17123;
    output \Kp[4] ;
    input n17122;
    output \Kp[3] ;
    input n17121;
    output \Kp[2] ;
    input n17120;
    output \Kp[1] ;
    input n17119;
    output [23:0]gearBoxRatio;
    input n17118;
    input n17117;
    input n17116;
    output n4;
    output \FRAME_MATCHER.state_31__N_2426[2] ;
    output n7;
    input n17115;
    input n17114;
    input n17113;
    input n17112;
    input n17111;
    input n17110;
    input n17109;
    input n17108;
    input n17107;
    input n17106;
    input n17105;
    input n17104;
    input n17103;
    input n17102;
    input n17101;
    input n17100;
    input n17099;
    input n17098;
    input n17097;
    input n17096;
    output [23:0]IntegralLimit;
    input n17095;
    input n17094;
    input n17093;
    input n17092;
    input n17091;
    input n17090;
    input n17089;
    input n17088;
    input n17087;
    input n17086;
    input n17085;
    input n17084;
    input n17083;
    input n17082;
    input n17081;
    input n17080;
    input n17079;
    input n17078;
    input n17077;
    input n17076;
    input n17075;
    input n17074;
    output n36885;
    output n4299;
    output n4298;
    output n4309;
    output n4308;
    output n4307;
    output n4311;
    output LED_c;
    output n4310;
    output n4313;
    output n4312;
    output n4315;
    output n4314;
    input n16832;
    input n16986;
    input n33975;
    input n16967;
    input n16965;
    input n16964;
    input n16963;
    output \Ki[0] ;
    input n16962;
    output \Kp[0] ;
    input n16961;
    output n4292;
    output n4297;
    output n4296;
    output n4295;
    output n4294;
    output n4293;
    output n4306;
    output n4305;
    output n4304;
    output n4303;
    output n4302;
    output n4301;
    output n5;
    output n318;
    output \r_Clock_Count[3] ;
    input n16918;
    output [2:0]r_Bit_Index;
    input n16915;
    input n16911;
    output \r_Clock_Count[1] ;
    input n16890;
    output \r_Clock_Count[8] ;
    input n16893;
    output \r_Clock_Count[7] ;
    input n16905;
    input n16899;
    output \r_Clock_Count[5] ;
    input n17029;
    input n17566;
    output [2:0]r_SM_Main;
    output n26602;
    output n320;
    input VCC_net;
    output n4613;
    output n26612;
    output n16641;
    output n16772;
    output tx_o;
    output tx_enable;
    output n313;
    output n314;
    input n16981;
    input n16979;
    output n316;
    output n3;
    output n29;
    input n16872;
    output \r_Clock_Count[6] ;
    input n16869;
    output \r_Clock_Count[7]_adj_3 ;
    input n16881;
    output \r_Clock_Count[3]_adj_4 ;
    input n16887;
    output \r_Clock_Count[1]_adj_5 ;
    input n17005;
    output [2:0]r_Bit_Index_adj_13;
    input n17002;
    input n17550;
    output r_Rx_Data;
    input PIN_13_N_105;
    output n219;
    output n220;
    output n30;
    output n223;
    output n3_adj_9;
    output n225;
    output n15459;
    output n4_adj_10;
    output n16746;
    output n16635;
    input n17012;
    input n17011;
    input n17010;
    input n17009;
    input n17008;
    input n17007;
    input n17006;
    output n4591;
    output n24014;
    output n4_adj_11;
    output n4_adj_12;
    output n15454;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n13231;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire Kp_23__N_839, n22, n17442, n16104, n20, n17441, n17440, 
        n17439, n6, n15871, n4_c, Kp_23__N_844, n28, n17438;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n10, n34675, n26, Kp_23__N_926, n35069, n34792, n34757, 
        n10_adj_3896, n34639, n17322, n17437, n17436, n17435, n17434, 
        n17433, n17432, n17431, n17430;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    
    wire n17333, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n3_c, n17429, n17428, n17427, n17426, n16353, n29_c, 
        n27939, n27940, n3_adj_3897, n31, n37983;
    wire [31:0]\FRAME_MATCHER.state_31__N_2490 ;
    
    wire n17425, n2_adj_3898, n27938, n2030, n2_adj_3899, n27937, 
        n2_adj_3900, n27936, n1507, n35060, n17351, n17323, n15617, 
        n17350, n34785, n34985, n17349, n17348, n17347, n17346, 
        n17332, n34905, n16423, n15986, n10_adj_3901, n17345, n17344, 
        n17343, n17331, n16026, n35063, n30619, n34870, n16927;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire n17324, n30573, n14, n17629, n17630, n16942, n30534, 
        n34726, n35028, n15, n16457, n35143, n17325, n34976, n16930, 
        n34909, n16999, n16996, n30591, n34912, n17032, n31249, 
        n6_adj_3902, n31226, n35134, n35234, n17476;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    
    wire n17477, n17390, n17389;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n17456, n17457, n17458, n17459, n17460, n17461, n17462, 
        n17388, n17448, n17449, n17450, n17451, n17452, n17453, 
        n17330, n17387, n17478, n17329, n17474, n17475, n17472, 
        n17473, n17470;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    
    wire n17471, n17468, n17469, n17466, n17467, n17328, n17463, 
        n17464, n17465, n17454, n17455, n17444, n17445, n17446, 
        n17447, n17342;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    
    wire n17327, n17326, n17443, n17321, n17320, n17319, n17318, 
        n34813, n6_adj_3903, n1593, n17317, n17316, n17315, n35182, 
        n35004, n34688, n1504, n17314, n17313, n17386, n17385, 
        n17384, n17383, n17382, n17381, n17380, n17379, n17312, 
        n17311, n17310, n14_adj_3904, n17309, n34795, n16476, n35103, 
        n35118, n15_adj_3905, n17404;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    
    wire n17308, n17307, n35072, n16359, n30571, n17306, n17341, 
        n17340, n2_adj_3906, n27935, n34991, n1513, n35214, n15171, 
        n17339, n34997, n1667, n17338, n34740, n12, n34851, n35078, 
        n16, n16166, n35041, n35081, n17, n15831, n30523, n17337, 
        n17336, n17335, n24008, n34654, n17359, n21, n23, n22_adj_3907, 
        n38053, n30_c, n17360, n35031, n28_adj_3908, n17378, n32, 
        n17361, n35258, n35115, n30_adj_3909, n35057, n35141, n15788, 
        n31_adj_3910, n35100, n29_adj_3911, n35201, n17362, n17363, 
        n15923, n34861, n34839, n16259, n35106, n15713, n34874, 
        n30559, n10_adj_3912, n35192, n34835, n16110, n14_adj_3913, 
        n6_adj_3914, n34884, n6_adj_3915, n15591, n34931, n34877, 
        n17364, n1829, n34881, n34832, n6_adj_3916, n15693, n30611, 
        n30613, n6_adj_3917, n17365, n34748, n35208, n34709, n34778, 
        n34718, n35211, n6_adj_3918, n34715, n35038, n34953, n17366, 
        n35151, n8, n34651;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    
    wire n17415, n17416, n34691, n35261, n13862, n17305, n16085, 
        n17304, n16116, n35097, n6_adj_3919, n17296;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    
    wire n17417, n5_c, n6_adj_3920, n34800, n17_adj_3921, n17377, 
        n6_adj_3922, n2_adj_3923, n27934, n34751, n35044, n26_adj_3924, 
        n18, n31_adj_3925;
    wire [0:0]n3241;
    wire [2:0]r_SM_Main_2__N_3323;
    
    wire n3243, n16074, n35051, n16366, n17418, n17419, n34950, 
        n34754, n18_adj_3926, n17420, n17_adj_3927, n15775, n19, 
        n32_adj_3928, n16119, n37, n34769, n34, n17421, n17422, 
        n34816, n36, n35, n39, n41, n37063, n2_adj_3929, n27933, 
        \FRAME_MATCHER.rx_data_ready_prev , n17424, n14_adj_3930, n34643, 
        n9, n34744, n30528, n30543, n17423, n17403, n10_adj_3931, 
        n2_adj_3932, n27932, n34858, n34806, n10_adj_3933, n35019, 
        n34_adj_3934, n22_adj_3935, n23_adj_3936, n38, n34789, n31279, 
        n36_adj_3937, n37_adj_3938, n35195, n35_adj_3939, n34921, 
        n17402, n2_adj_3940, n27931, n35140, n14_adj_3941, n30555, 
        n37194, n16137, n15944, n16_adj_3942, n16286, n15_adj_3943, 
        n16232, n16289, n22_adj_3944, n15939, n15794, n15756, n20_adj_3945, 
        n15803, n24, n15798, n16142, n31_adj_3946, n4291, n17391;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    
    wire n17376, n17375, n17401, n35198, n31275, n12_adj_3947, n35279, 
        n34970, n15165, n15586, n2_adj_3948, n27930, n17400, n6_adj_3949, 
        n34855, n15154, n35066, n10_adj_3950, n29_adj_3951, n47, 
        n34530, n1285, n6_adj_3952, n34957, n2_adj_3953, n27929, 
        n6_adj_3954, n34988, n18_adj_3955, n35166, n19_adj_3956, n17_adj_3957, 
        n18_adj_3958, n2_adj_3959, n27928, n35232, n21_adj_3960, n35146, 
        n20_adj_3961, n35131, n24_adj_3962, n30998, n4_adj_3963, n35380;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n19_adj_3964, n2_adj_3965, n27927, n40561, n5_adj_3966, n38192, 
        n43149, n38193, n101, n38146, n17399, n38148, n43161, 
        n43155, n38147, n17398, n17397, n2_adj_3967, n27926, n19_adj_3968, 
        n40556, n2_adj_3969, n27925, n5_adj_3970, n38189, n43143, 
        n38190, n38143, n38145, n43173, n43167, n38144, n2_adj_3971, 
        n27924, n19_adj_3972, n40551, n5_adj_3973, n2_adj_3974, n27923, 
        n38186, n43137, n38187, n38170, n38172, n43185, n43179, 
        n38171, n19_adj_3975, n6_adj_3976, n5_adj_3977, n38183, n43131, 
        n38184, n38167, n38169, n43197, n43191, n38168, n19_adj_3978, 
        n40513, n19_adj_3979, n6_adj_3980, n5_adj_3981, n5_adj_3982, 
        n38180, n38150, n43125, n38181, n38164, n38166, n43209, 
        n43203, n38165, n43107, n38151, n17396, n38155, n17395, 
        n17374, n38157, n19_adj_3983, n43245, n43239, n38156, n6_adj_3984, 
        n5_adj_3985, n38177, n43119, n38178, n38161, n38163, n43221, 
        n43215, n38162, n34647, n34101, n17394, n19_adj_3986, n40536, 
        n5_adj_3987, n38153, n43113, n38154, n38158, n38160, n43233, 
        n43227, n38159, n40164, n27958, n4_adj_3988, n4368, n30171, 
        n37236, n34673, n34521, n34671, n6_adj_3989, n34772, n35054, 
        n34973, n36175, n7_c, n2_adj_3990, n27922, n2_adj_3991, 
        n27921, n24911, n139, n8_adj_3992, n4_adj_3993, n43479, 
        n15448, n40215, n40163, n27957, \FRAME_MATCHER.i_31__N_2389 , 
        n161, n24117, n13978, n35109, n34803, n10_adj_3994, n15780, 
        n13, n40162, n27956, n4_adj_3995, n34845, n12_adj_3996, 
        n16160, Kp_23__N_896, n34731, n34829, Kp_23__N_893;
    wire [7:0]n7813;
    
    wire n27955, Kp_23__N_858, n17156;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    
    wire n34631, n17405, n22677, n17150, n17406, n17148;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    
    wire n12859, n10_adj_3997;
    wire [7:0]\data_in[0]_c ;   // verilog/coms.v(93[12:19])
    
    wire n14_adj_3998, n15514, n15329, n4_adj_3999, n15342, n20_adj_4000, 
        n19_adj_4001, n38076, n63_adj_4002, n10_adj_4003, n15552, 
        n14_adj_4004, n15_adj_4005, n17140, n27954, n16_adj_4006, 
        n17_adj_4007, n15445, n16_adj_4008, n17_adj_4009, n31_adj_4010, 
        n63_adj_4011, n18_adj_4012, n20_adj_4013, n15_adj_4014, n22667, 
        n41_adj_4015, \FRAME_MATCHER.i_31__N_2392 , n3741, n42, n2720, 
        n43, n34668, n1205, n17_adj_4016, n26928, n34051, n42_adj_4017, 
        n40, n41_adj_4018, n39_adj_4019, n38_adj_4020, n37_adj_4021, 
        n48, n43_adj_4022, n15540, n10_adj_4023, n84, tx_transmit_N_3220, 
        n15437, n42349;
    wire [31:0]n92;
    
    wire n5_adj_4026, n30072, n1, n43474, n35144, n30653, n36946, 
        n30603, n6_adj_4027, n36900, n16_adj_4028, n35034, n17_adj_4029, 
        n6_adj_4030, n36211, n35255, n14_adj_4031, n9_adj_4032, n35276, 
        n35804, n12_adj_4033, n36587, n36281, n7_adj_4034, n18939;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    wire n10_adj_4035, n14_adj_4036, n15_adj_4037, n34523, n8_adj_4038, 
        n7_adj_4039, n6_adj_4040, n27953, n3_adj_4041, n17353, n27952, 
        n17373, n17372, n2_adj_4042, n27951, n17371, n17370, n17369, 
        n3_adj_4043, n3_adj_4044, n3_adj_4045, n3_adj_4046, n3_adj_4047, 
        n3_adj_4048, n3_adj_4049, n3_adj_4050, n3_adj_4051, n3_adj_4052, 
        n3_adj_4053, n3_adj_4054, n3_adj_4055, n3_adj_4056, n3_adj_4057, 
        n3_adj_4058, n3_adj_4059, n2_adj_4060, n3_adj_4061, n2_adj_4062, 
        n3_adj_4063, n2_adj_4064, n3_adj_4065, n2_adj_4066, n3_adj_4067, 
        n2_adj_4068, n3_adj_4069, n2_adj_4070, n3_adj_4071, n2_adj_4072, 
        n3_adj_4073, n2_adj_4074, n3_adj_4075, n2_adj_4076, n3_adj_4077, 
        n2_adj_4078, n3_adj_4079, n2_adj_4080, n3_adj_4081, n2_adj_4082, 
        n3_adj_4083, n3_adj_4084, n16593, n36199, n36969, n34990, 
        n35126, n34910, n33967, n33969, n34111, n33977, n34113, 
        n34043, n7_adj_4085, n8_adj_4086, n34115, n34041, n34117, 
        n34039, n7_adj_4087, n8_adj_4088, n34119, n34037, n34121, 
        n8_adj_4089, n34123, n34035, n34125, n34033, n34127, n34031, 
        n34129, n34029, n7_adj_4090, n8_adj_4091, n34131, n8_adj_4092, 
        n7_adj_4093, n8_adj_4094, n23956, n24611, n7_adj_4095, n8_adj_4096, 
        n34133, n34027, n34135, n34025, n34137, n34023, n34139, 
        n8_adj_4097, n34141, n34021, n34143, n34019, n34145, n34017, 
        n7_adj_4098, n8_adj_4099, n34147, n34015, n34149, n34013, 
        n7_adj_4100, n8_adj_4101, n27950, n34848, n35226, n10_adj_4102, 
        n35240, n17368, n27949, n27942, n27943, n16737, n34864, 
        n12905, n17367, n27948, n27947, n43242, n43236, n43230, 
        n43224, n43218, n43212, n27946, n24524, n15657, n35285, 
        n17414;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    
    wire n17413, n17412, n17411, n17410, n27945, n17393, n27944, 
        n6_adj_4103, n34763, n27941, n43206, n17352, n121, n10_adj_4104, 
        n10_adj_4105, n30585, n37977, n35282, n35243, n17358, n17357, 
        n17356, n43200, n17334, n34693, n34635, n17392, n34627, 
        n17407, n17408, n17409, n34810, n17355, n17354, n34887, 
        n43194, n10_adj_4106, n24172, n43188, n43182, n43176, n22591, 
        n43170, n43164, n43158, n43152, n43146, n43140, n34960, 
        n31273, n12_adj_4107, n8_adj_4108, n31330, n34678, n31269, 
        n34737, n16283, n31234, n35229, n35128, n34901, n31284, 
        n36194, n35137, n35270, n10_adj_4109, n34967, n15990, n6_adj_4110, 
        n34712, n30623, n35022, n35001, Kp_23__N_1353, n36871, n35246, 
        n15671, n35169, n14_adj_4111, n10_adj_4112, n34979, n35774, 
        n16057, n36362, n31332, n6_adj_4113, n35188, n26_adj_4114, 
        n24_adj_4115, n35088, n25, n35025, n34916, n23_adj_4116, 
        n35252, n35012, n16218, n34867, n35172, n35176, n20_adj_4117, 
        n34766, n19_adj_4118, n34702, n16479, n21_adj_4119, n34819, 
        n35112, n35220, n35273, Kp_23__N_969, n35016, n12_adj_4120, 
        n15917, n16391, n35179, n35009, n10_adj_4121, Kp_23__N_1083, 
        n34699, n14_adj_4122, n35084, n15862, n12_adj_4123, n34684, 
        n6_adj_4124, n35047, Kp_23__N_1430, n31345, n30605, n16394, 
        n6_adj_4125, n6_adj_4126, n35160, n35237, n35075, n35157, 
        n12_adj_4127, n14_adj_4128, n10_adj_4129, n31251, n35121, 
        n22_adj_4130, n35163, n32_adj_4131, n36_adj_4132, n34_adj_4133, 
        n35_adj_4134, n16277, n35249, n33, n15828, n28_adj_4135, 
        n35223, n26_adj_4136, n35205, n27, n25_adj_4137, n36545, 
        n34944, n46, n34890, n44, n35091, n45, n35094, n43_adj_4138, 
        n42_adj_4139, n41_adj_4140, n52, n31271, n47_adj_4141, n34994, 
        n20_adj_4142, n34898, n19_adj_4143, n21_adj_4144, n30609, 
        n34940, n8_adj_4145, n16183, n43134, n35148, n34925, n43128, 
        n34825, n34964, n30553, n35264, n6_adj_4147, n10_adj_4148, 
        n31261, n10_adj_4149, n37099, n6_adj_4150, n16400, n6_adj_4151, 
        n35185, n14_adj_4152, n6_adj_4153, n6_adj_4154, n34928, n35267, 
        n34721, n16_adj_4155, n17_adj_4156, n31258, n20_adj_4157, 
        n19_adj_4158, n21_adj_4159, n36828, n8_adj_4160, n12_adj_4161, 
        n36991, n12_adj_4162, n4_adj_4163, n36693, n43740, n14_adj_4164, 
        n13_adj_4165, n12_adj_4166, n36974, n20_adj_4167, n11, n15_adj_4168, 
        n8_adj_4169, n36119, n34935, n36799, n43122, n43116, n43110, 
        n11_adj_4170, n43104, n8_adj_4171;
    
    SB_LUT4 i5_4_lut (.I0(\data_in_frame[1] [7]), .I1(n13231), .I2(\data_in_frame[0] [0]), 
            .I3(Kp_23__N_839), .O(n22));
    defparam i5_4_lut.LUT_INIT = 16'h2112;
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n17442));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_3_lut (.I0(n16104), .I1(\data_in_frame[2] [1]), .I2(Kp_23__N_839), 
            .I3(GND_net), .O(n20));
    defparam i3_3_lut.LUT_INIT = 16'h1414;
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n17441));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n17440));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n17439));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[3] [3]), .I3(n6), .O(n15871));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(n4_c), .I1(n22), .I2(Kp_23__N_844), .I3(\data_in_frame[1] [0]), 
            .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h0440;
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n17438));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut (.I0(Kp_23__N_839), .I1(n10), .I2(n34675), .I3(\data_in_frame[1] [5]), 
            .O(n26));
    defparam i9_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[5] [1]), .I1(Kp_23__N_926), .I2(n35069), 
            .I3(n34792), .O(n34757));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12640_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n17322));
    defparam i12640_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n17437));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n17436));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n17435));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n17434));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n17433));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n17432));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n17431));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n17430));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n17333));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3_c));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n17429));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n17428));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n17427));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n17426));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [6]), .I3(n16353), .O(n29_c));
    defparam i12_4_lut.LUT_INIT = 16'h0080;
    SB_CARRY add_41_21 (.CI(n27939), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n27940));
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[1] [2]), .I1(n28), .I2(n20), 
            .I3(n3_adj_3897), .O(n31));
    defparam i14_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i16_4_lut (.I0(n31), .I1(n29_c), .I2(n37983), .I3(n26), 
            .O(\FRAME_MATCHER.state_31__N_2490 [3]));
    defparam i16_4_lut.LUT_INIT = 16'h0800;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n17425));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_20_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n27938), .O(n2_adj_3898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_20 (.CI(n27938), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n27939));
    SB_LUT4 add_41_19_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n27937), .O(n2_adj_3899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_19 (.CI(n27937), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n27938));
    SB_LUT4 add_41_18_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n27936), .O(n2_adj_3900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[15] [4]), 
            .I2(n1507), .I3(GND_net), .O(n35060));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n17351));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12641_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n17323));
    defparam i12641_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15617));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n17350));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_876 (.I0(\data_out_frame[19] [6]), .I1(n35060), 
            .I2(n34785), .I3(\data_out_frame[19] [5]), .O(n34985));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_876.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n17349));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n17348));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n17347));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n17346));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n17332));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_877 (.I0(\data_out_frame[19] [0]), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n34905));
    defparam i2_3_lut_adj_877.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_878 (.I0(n16423), .I1(n15986), .I2(\data_out_frame[18] [5]), 
            .I3(n34905), .O(n10_adj_3901));
    defparam i4_4_lut_adj_878.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n17345));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n17344));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n17343));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n17331));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_879 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16026));
    defparam i1_2_lut_adj_879.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_880 (.I0(n35063), .I1(\data_out_frame[20] [1]), 
            .I2(n30619), .I3(GND_net), .O(n34870));
    defparam i2_3_lut_adj_880.LUT_INIT = 16'h9696;
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
           .D(n16927));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12642_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n17324));
    defparam i12642_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut (.I0(n30573), .I1(\data_out_frame[20] [5]), .I2(\data_out_frame[18] [4]), 
            .I3(GND_net), .O(n14));   // verilog/coms.v(72[16:43])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
           .D(n17629));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
           .D(n17630));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
           .D(n16942));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut (.I0(n30534), .I1(\data_out_frame[15] [7]), .I2(n34726), 
            .I3(n35028), .O(n15));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n16457), .I2(n14), .I3(\data_out_frame[18] [3]), 
            .O(n35143));   // verilog/coms.v(72[16:43])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12643_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n17325));
    defparam i12643_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_881 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [4]), .I3(\data_out_frame[20] [6]), 
            .O(n34976));
    defparam i3_4_lut_adj_881.LUT_INIT = 16'h6996;
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n17581));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n17582));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n17583));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n17584));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n17585));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n17586));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n17587));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n17574));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n17575));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n17576));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n17577));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n17578));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
           .D(n16930));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_882 (.I0(n34976), .I1(n35143), .I2(\data_out_frame[18] [5]), 
            .I3(GND_net), .O(n34909));
    defparam i2_3_lut_adj_882.LUT_INIT = 16'h9696;
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
           .D(n16999));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
           .D(n16996));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_883 (.I0(n30591), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34912));
    defparam i1_2_lut_adj_883.LUT_INIT = 16'h6666;
    SB_DFF byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
           .D(n17032));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n17595));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n17596));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n17593));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n17594));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n17591));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n17592));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_2_lut (.I0(n31249), .I1(\data_out_frame[12] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3902));
    defparam i2_2_lut.LUT_INIT = 16'h9999;
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n17588));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n17589));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n17590));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n17579));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n17580));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n17495));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut (.I0(n34912), .I1(\data_out_frame[14] [6]), .I2(n6_adj_3902), 
            .I3(n31226), .O(n35134));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n17496));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n17497));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n17498));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n17499));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n17500));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n17501));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n17487));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n17488));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n17489));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n17490));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n17491));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n17492));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_884 (.I0(n30591), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35234));
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n17476));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n17477));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n17390));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n17389));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n43272));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n17456));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n17457));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n17458));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n17459));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n17460));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n17461));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n17462));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n17388));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n17448));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n17449));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n17450));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n17451));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n17452));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n17453));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n17330));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n17493));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n17494));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n17387));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n17478));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n17479));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n17480));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n17481));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n17482));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n17483));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n17484));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n17485));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n17486));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n17329));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n17474));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n17475));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n17472));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n17473));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n17470));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n17471));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n17468));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n17469));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n17466));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n17467));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n17328));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n17463));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n17464));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n17465));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n17454));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n17455));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n17444));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n17445));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n17446));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n17447));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n17342));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n17327));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n17326));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n17325));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n17324));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n17443));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n17323));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n17322));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n17321));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n17320));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n17319));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n17318));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_885 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(n34813), .I3(n6_adj_3903), .O(n1593));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_885.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n17317));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n17316));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n17315));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_886 (.I0(\data_out_frame[8] [4]), .I1(n35182), 
            .I2(n35004), .I3(n34688), .O(n1504));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n17314));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n17313));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n17386));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n17385));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n17384));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n17383));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n17382));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n17381));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n17380));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n17379));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n17312));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_18 (.CI(n27936), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n27937));
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n17311));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n17310));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_adj_887 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[18] [0]), 
            .I2(\data_out_frame[13] [5]), .I3(GND_net), .O(n14_adj_3904));   // verilog/coms.v(72[16:43])
    defparam i5_3_lut_adj_887.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n17309));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_888 (.I0(n34795), .I1(n16476), .I2(n35103), .I3(n35118), 
            .O(n15_adj_3905));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n17404));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n17308));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n17307));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i8_4_lut_adj_889 (.I0(n15_adj_3905), .I1(n35072), .I2(n14_adj_3904), 
            .I3(n16359), .O(n30571));   // verilog/coms.v(72[16:43])
    defparam i8_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n17306));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n17341));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n17340));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_17_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n27935), .O(n2_adj_3906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_890 (.I0(n34991), .I1(\data_out_frame[15] [1]), 
            .I2(n1513), .I3(GND_net), .O(n35214));
    defparam i2_3_lut_adj_890.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_891 (.I0(n15171), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30534));
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n17339));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_892 (.I0(\data_out_frame[13] [2]), .I1(n34997), 
            .I2(\data_out_frame[13] [1]), .I3(GND_net), .O(n1667));   // verilog/coms.v(83[17:63])
    defparam i2_3_lut_adj_892.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n17338));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_adj_893 (.I0(n34740), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n12));
    defparam i5_3_lut_adj_893.LUT_INIT = 16'h9696;
    SB_LUT4 i12644_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n17326));
    defparam i12644_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_894 (.I0(n34851), .I1(\data_out_frame[15] [1]), 
            .I2(n35078), .I3(n34997), .O(n16));
    defparam i6_4_lut_adj_894.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n16166), .I1(n35041), .I2(n35081), .I3(n34991), 
            .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_895 (.I0(n17), .I1(n34740), .I2(n16), .I3(n15831), 
            .O(n30523));
    defparam i9_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n17337));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n17336));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n17335));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12677_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n17359));
    defparam i12677_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14_4_lut_adj_896 (.I0(n21), .I1(n23), .I2(n22_adj_3907), 
            .I3(n38053), .O(n30_c));
    defparam i14_4_lut_adj_896.LUT_INIT = 16'hfeff;
    SB_LUT4 i12678_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n17360));
    defparam i12678_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut (.I0(n31249), .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[11] [0]), 
            .I3(n35031), .O(n28_adj_3908));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n17378));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14_3_lut (.I0(\data_out_frame[14] [5]), .I1(n28_adj_3908), 
            .I2(n30523), .I3(GND_net), .O(n32));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12679_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n17361));
    defparam i12679_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12_4_lut_adj_897 (.I0(\data_out_frame[17] [0]), .I1(n35258), 
            .I2(n30534), .I3(n35115), .O(n30_adj_3909));
    defparam i12_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n35057), .I1(n35141), .I2(n34997), .I3(n15788), 
            .O(n31_adj_3910));
    defparam i13_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_898 (.I0(n35214), .I1(n35100), .I2(\data_out_frame[14] [4]), 
            .I3(\data_out_frame[14] [3]), .O(n29_adj_3911));
    defparam i11_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n29_adj_3911), .I1(n31_adj_3910), .I2(n30_adj_3909), 
            .I3(n32), .O(n35201));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12680_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n17362));
    defparam i12680_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_899 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n15986));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i12681_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n17363));
    defparam i12681_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_900 (.I0(\data_out_frame[18] [3]), .I1(n15923), 
            .I2(GND_net), .I3(GND_net), .O(n34861));
    defparam i1_2_lut_adj_900.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34726));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_902 (.I0(\data_out_frame[6] [5]), .I1(n35103), 
            .I2(n34839), .I3(n16259), .O(n1513));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_903 (.I0(\data_out_frame[11] [5]), .I1(n35106), 
            .I2(n34839), .I3(n15713), .O(n15171));
    defparam i3_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\data_out_frame[13] [6]), .I1(n1513), 
            .I2(GND_net), .I3(GND_net), .O(n35028));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_905 (.I0(n34874), .I1(n35028), .I2(n15171), .I3(GND_net), 
            .O(n30559));
    defparam i2_3_lut_adj_905.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_906 (.I0(n35072), .I1(\data_out_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3912));   // verilog/coms.v(73[16:27])
    defparam i2_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_907 (.I0(n35192), .I1(\data_out_frame[16] [0]), 
            .I2(n34835), .I3(n16110), .O(n14_adj_3913));   // verilog/coms.v(73[16:27])
    defparam i6_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_908 (.I0(\data_out_frame[18] [2]), .I1(n14_adj_3913), 
            .I2(n10_adj_3912), .I3(n34726), .O(n15923));   // verilog/coms.v(73[16:27])
    defparam i7_4_lut_adj_908.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[17] [7]), 
            .I2(n6_adj_3914), .I3(\data_out_frame[16] [0]), .O(n34884));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_909 (.I0(\data_out_frame[20] [4]), .I1(n16423), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3915));
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_910 (.I0(n30559), .I1(n15591), .I2(n34861), .I3(n6_adj_3915), 
            .O(n34931));
    defparam i4_4_lut_adj_910.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_911 (.I0(n34884), .I1(\data_out_frame[20] [3]), 
            .I2(n15923), .I3(GND_net), .O(n34877));
    defparam i2_3_lut_adj_911.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_912 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n15591));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_adj_912.LUT_INIT = 16'h6666;
    SB_LUT4 i12682_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n17364));
    defparam i12682_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1073_2_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1829));   // verilog/coms.v(69[16:27])
    defparam i1073_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34881));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_914 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(n34832), .I3(n6_adj_3916), .O(n15693));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_915 (.I0(n30611), .I1(n15693), .I2(GND_net), 
            .I3(GND_net), .O(n30613));
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_916 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[13] [7]), 
            .I2(n34740), .I3(n6_adj_3917), .O(n16423));
    defparam i4_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i12683_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n17365));
    defparam i12683_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_917 (.I0(\data_out_frame[9] [5]), .I1(n34748), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[7] [4]), .O(n15788));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_918 (.I0(\data_out_frame[12] [0]), .I1(n35208), 
            .I2(n15788), .I3(GND_net), .O(n34709));
    defparam i2_3_lut_adj_918.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_919 (.I0(\data_out_frame[9] [7]), .I1(n34778), 
            .I2(\data_out_frame[10] [0]), .I3(\data_out_frame[12] [1]), 
            .O(n35057));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_920 (.I0(n34718), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n35211));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_920.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_921 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34748));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_921.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_922 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3918));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_922.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_923 (.I0(n34748), .I1(n34715), .I2(n35038), .I3(n6_adj_3918), 
            .O(n34953));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i12684_3_lut_4_lut (.I0(n24008), .I1(n34654), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n17366));
    defparam i12684_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_924 (.I0(\data_out_frame[14] [2]), .I1(n35211), 
            .I2(n35057), .I3(n34709), .O(n16457));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_924.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_925 (.I0(n16457), .I1(n34953), .I2(GND_net), 
            .I3(GND_net), .O(n35151));
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h6666;
    SB_LUT4 i12733_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n17415));
    defparam i12733_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12734_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n17416));
    defparam i12734_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_926 (.I0(n34691), .I1(\data_out_frame[12] [4]), 
            .I2(n30611), .I3(GND_net), .O(n31249));
    defparam i2_3_lut_adj_926.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_927 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16166));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_928 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[10] [5]), .I3(n16166), .O(n34813));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_929 (.I0(n34813), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n35261));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_929.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_930 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n34832));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_930.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_931 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[11] [4]), .I3(n13862), .O(n35106));
    defparam i3_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_932 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[5] [2]), .I3(GND_net), .O(n35208));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_932.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n17305));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16085));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_out_frame[6] [7]), .I1(n34718), 
            .I2(GND_net), .I3(GND_net), .O(n15713));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n17304));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut_adj_935 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[7] [1]), 
            .I2(n15713), .I3(n16085), .O(n34740));
    defparam i2_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_CARRY add_41_17 (.CI(n27935), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n27936));
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n17303));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n17302));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n17301));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n17300));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_936 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35038));
    defparam i1_2_lut_adj_936.LUT_INIT = 16'h6666;
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n17299));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_937 (.I0(\data_out_frame[8] [0]), .I1(n16116), 
            .I2(\data_out_frame[10] [1]), .I3(\data_out_frame[5] [6]), .O(n35097));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_937.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_938 (.I0(\data_out_frame[9] [6]), .I1(n35097), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3919));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_938.LUT_INIT = 16'h6666;
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n17298));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n17297));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
           .D(n17296));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n17295));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n17294));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n17293));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12735_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n17417));
    defparam i12735_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_939 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[9] [5]), .I3(n6_adj_3919), .O(n34715));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n17292));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_4_lut_adj_940 (.I0(n5_c), .I1(\data_in_frame[21] [7]), .I2(n6_adj_3920), 
            .I3(n34800), .O(n17_adj_3921));
    defparam i1_4_lut_adj_940.LUT_INIT = 16'hde7b;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n17377));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_941 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3922));
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n17291));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_16_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n27934), .O(n2_adj_3923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_16_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n17290));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n17289));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_16 (.CI(n27934), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n27935));
    SB_LUT4 i4_4_lut_adj_942 (.I0(n34751), .I1(\data_out_frame[7] [6]), 
            .I2(n35044), .I3(n6_adj_3922), .O(n34691));
    defparam i4_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n17288));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n17287));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n17286));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n17285));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n17284));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n17283));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n17282));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i15_4_lut (.I0(n17_adj_3921), .I1(n30_c), .I2(n26_adj_3924), 
            .I3(n18), .O(n31_adj_3925));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n17281));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n17280));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n17279));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n17278));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSR tx_transmit_3205 (.Q(r_SM_Main_2__N_3323[0]), .C(clk32MHz), 
            .D(n3241[0]), .R(n3243));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_943 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16074));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_out_frame[10] [0]), .I1(n34691), 
            .I2(GND_net), .I3(GND_net), .O(n35051));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_945 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16116));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_945.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_946 (.I0(\data_out_frame[8] [1]), .I1(n16366), 
            .I2(\data_out_frame[5] [6]), .I3(n16116), .O(n34751));   // verilog/coms.v(69[16:62])
    defparam i3_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i12736_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n17418));
    defparam i12736_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_947 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35041));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_947.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_948 (.I0(\data_out_frame[10] [3]), .I1(n35041), 
            .I2(n34751), .I3(\data_out_frame[6] [1]), .O(n30611));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i12737_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n17419));
    defparam i12737_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_949 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35044));
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34950));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34754));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_952 (.I0(n34754), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[6] [5]), .I3(\data_out_frame[6] [3]), .O(n18_adj_3926));   // verilog/coms.v(72[16:27])
    defparam i7_4_lut_adj_952.LUT_INIT = 16'h6996;
    SB_LUT4 i12738_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n17420));
    defparam i12738_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_3_lut (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n17_adj_3927));   // verilog/coms.v(72[16:27])
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_953 (.I0(n34950), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[6] [1]), .I3(n15775), .O(n19));   // verilog/coms.v(72[16:27])
    defparam i8_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_954 (.I0(n35044), .I1(n19), .I2(n17_adj_3927), 
            .I3(n18_adj_3926), .O(n32_adj_3928));   // verilog/coms.v(71[16:34])
    defparam i10_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_955 (.I0(n16119), .I1(\data_out_frame[11] [5]), 
            .I2(n31226), .I3(\data_out_frame[11] [2]), .O(n37));   // verilog/coms.v(71[16:34])
    defparam i15_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_956 (.I0(\data_out_frame[11] [6]), .I1(n34769), 
            .I2(\data_out_frame[9] [3]), .I3(\data_out_frame[9] [4]), .O(n34));   // verilog/coms.v(71[16:34])
    defparam i12_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i12739_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n17421));
    defparam i12739_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12740_3_lut_4_lut (.I0(n8), .I1(n34651), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n17422));
    defparam i12740_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_957 (.I0(\data_out_frame[11] [4]), .I1(n34816), 
            .I2(n35051), .I3(n16074), .O(n36));   // verilog/coms.v(71[16:34])
    defparam i14_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_958 (.I0(n35182), .I1(\data_out_frame[9] [1]), 
            .I2(n34715), .I3(\data_out_frame[11] [3]), .O(n35));   // verilog/coms.v(71[16:34])
    defparam i13_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i17_3_lut (.I0(n35004), .I1(n34), .I2(\data_out_frame[7] [4]), 
            .I3(GND_net), .O(n39));   // verilog/coms.v(71[16:34])
    defparam i17_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(\data_out_frame[8] [1]), .I2(n32_adj_3928), 
            .I3(n34839), .O(n41));   // verilog/coms.v(71[16:34])
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n41), .I1(n39), .I2(n35), .I3(n36), .O(n37063));   // verilog/coms.v(71[16:34])
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_15_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n27933), .O(n2_adj_3929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_15 (.CI(n27933), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n27934));
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3206  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n17424));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n17277));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_959 (.I0(n35038), .I1(\data_out_frame[12] [4]), 
            .I2(n34740), .I3(\data_out_frame[12] [3]), .O(n14_adj_3930));
    defparam i6_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i12629_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n17311));
    defparam i12629_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12630_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n17312));
    defparam i12630_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 i12631_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n17313));
    defparam i12631_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_961 (.I0(n9), .I1(n14_adj_3930), .I2(n34744), 
            .I3(n37063), .O(n30528));
    defparam i7_4_lut_adj_961.LUT_INIT = 16'h9669;
    SB_LUT4 i12632_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n17314));
    defparam i12632_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_962 (.I0(\data_out_frame[14] [7]), .I1(n30528), 
            .I2(GND_net), .I3(GND_net), .O(n30543));
    defparam i1_2_lut_adj_962.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n17276));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n17423));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n17422));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n17403));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_963 (.I0(n35051), .I1(n34778), .I2(\data_out_frame[14] [4]), 
            .I3(n35208), .O(n10_adj_3931));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_14_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n27932), .O(n2_adj_3932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_964 (.I0(n34858), .I1(\data_in_frame[5] [0]), .I2(n34792), 
            .I3(GND_net), .O(n34806));
    defparam i2_3_lut_adj_964.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_965 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3933));
    defparam i2_2_lut_adj_965.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n17275));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_14 (.CI(n27932), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n27933));
    SB_LUT4 i1_2_lut_adj_966 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34874));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_967 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16476));
    defparam i1_2_lut_adj_967.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_968 (.I0(n34874), .I1(n35019), .I2(n30591), 
            .I3(n30543), .O(n34_adj_3934));
    defparam i13_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_3935));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut_adj_970 (.I0(n23_adj_3936), .I1(n34_adj_3934), .I2(\data_out_frame[17] [4]), 
            .I3(n31249), .O(n38));
    defparam i17_4_lut_adj_970.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_971 (.I0(n34789), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[14] [6]), .I3(n31279), .O(n36_adj_3937));
    defparam i15_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_972 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[15] [6]), .I3(n22_adj_3935), .O(n37_adj_3938));
    defparam i16_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_973 (.I0(\data_out_frame[13] [7]), .I1(n35195), 
            .I2(\data_out_frame[13] [0]), .I3(n34881), .O(n35_adj_3939));
    defparam i14_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n35_adj_3939), .I1(n37_adj_3938), .I2(n36_adj_3937), 
            .I3(n38), .O(n34921));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12633_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n17315));
    defparam i12633_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n17402));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_13_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n27931), .O(n2_adj_3940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_13_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n17274));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_974 (.I0(\data_out_frame[17] [1]), .I1(n34921), 
            .I2(GND_net), .I3(GND_net), .O(n35140));
    defparam i1_2_lut_adj_974.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_975 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [3]), .O(n14_adj_3941));
    defparam i6_4_lut_adj_975.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_976 (.I0(\data_in_frame[0] [2]), .I1(n14_adj_3941), 
            .I2(n10_adj_3933), .I3(\data_in_frame[0] [1]), .O(n13231));
    defparam i7_4_lut_adj_976.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_977 (.I0(n34806), .I1(n34757), .I2(n15871), .I3(n30555), 
            .O(n37194));
    defparam i3_4_lut_adj_977.LUT_INIT = 16'hefff;
    SB_LUT4 i3_2_lut (.I0(n16137), .I1(n15944), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_3942));   // verilog/coms.v(228[9:81])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_978 (.I0(n16286), .I1(n15_adj_3943), .I2(n16232), 
            .I3(n16289), .O(n22_adj_3944));   // verilog/coms.v(228[9:81])
    defparam i9_4_lut_adj_978.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n15939), .I1(n15794), .I2(n15756), .I3(GND_net), 
            .O(n20_adj_3945));   // verilog/coms.v(228[9:81])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_979 (.I0(n15803), .I1(n22_adj_3944), .I2(n16_adj_3942), 
            .I3(n37194), .O(n24));   // verilog/coms.v(228[9:81])
    defparam i11_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_980 (.I0(n15798), .I1(n24), .I2(n20_adj_3945), 
            .I3(n16142), .O(n31_adj_3946));   // verilog/coms.v(228[9:81])
    defparam i12_4_lut_adj_980.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_981 (.I0(\FRAME_MATCHER.state [1]), .I1(n31_adj_3946), 
            .I2(n13231), .I3(GND_net), .O(n4291));
    defparam i2_3_lut_adj_981.LUT_INIT = 16'h0202;
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n17391));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n17376));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n17375));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n17401));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut_adj_982 (.I0(n35198), .I1(n35258), .I2(n31275), .I3(n35140), 
            .O(n12_adj_3947));
    defparam i5_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_983 (.I0(\data_out_frame[12] [5]), .I1(n12_adj_3947), 
            .I2(n35279), .I3(n34970), .O(n15165));
    defparam i6_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n15586));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n13862));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_LUT4 i12634_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n17316));
    defparam i12634_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_986 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16119));
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_CARRY add_41_13 (.CI(n27931), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n27932));
    SB_LUT4 add_41_12_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n27930), .O(n2_adj_3948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_12 (.CI(n27930), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n27931));
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n17400));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_987 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34769));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h6666;
    SB_LUT4 i12635_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n17317));
    defparam i12635_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16359));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_989 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16259));
    defparam i1_2_lut_adj_989.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_990 (.I0(\data_out_frame[7] [1]), .I1(n35118), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3949));
    defparam i1_2_lut_adj_990.LUT_INIT = 16'h6666;
    SB_LUT4 i12636_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34643), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n17318));
    defparam i12636_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_991 (.I0(n16259), .I1(\data_out_frame[8] [6]), 
            .I2(n34855), .I3(n6_adj_3949), .O(n15154));
    defparam i4_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_992 (.I0(n15154), .I1(n1507), .I2(GND_net), .I3(GND_net), 
            .O(n35066));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h6666;
    SB_LUT4 i12693_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n17375));
    defparam i12693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34688));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_994 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35195));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16366));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_996 (.I0(n29_adj_3951), .I1(n47), .I2(n34530), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n36839));
    defparam i3_4_lut_adj_996.LUT_INIT = 16'hfffb;
    SB_LUT4 mux_1046_i9_3_lut (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4291), .I3(GND_net), .O(n4300));
    defparam mux_1046_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12694_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n17376));
    defparam i12694_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_997 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15775));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_998 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [0]), 
            .I2(n35195), .I3(\data_out_frame[12] [7]), .O(n34851));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i529_2_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1285));   // verilog/coms.v(69[16:27])
    defparam i529_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_999 (.I0(\data_out_frame[15] [3]), .I1(n1285), 
            .I2(n35115), .I3(n6_adj_3952), .O(n34957));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_11_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n27929), .O(n2_adj_3953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_adj_1000 (.I0(n34957), .I1(n30619), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3954));
    defparam i2_2_lut_adj_1000.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[19] [6]), 
            .I2(n6_adj_3954), .I3(n34795), .O(n34988));
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'h9669;
    SB_CARRY add_41_11 (.CI(n27929), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n27930));
    SB_LUT4 i7_4_lut_adj_1002 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [1]), 
            .I2(n35063), .I3(\data_out_frame[18] [4]), .O(n18_adj_3955));
    defparam i7_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1003 (.I0(n35166), .I1(n16476), .I2(n34953), 
            .I3(\data_out_frame[18] [1]), .O(n19_adj_3956));
    defparam i8_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1004 (.I0(n19_adj_3956), .I1(n35134), .I2(n17_adj_3957), 
            .I3(n18_adj_3955), .O(n18_adj_3958));
    defparam i5_4_lut_adj_1004.LUT_INIT = 16'h9669;
    SB_LUT4 add_41_10_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n27928), .O(n2_adj_3959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut_adj_1005 (.I0(n31279), .I1(n34909), .I2(n35232), 
            .I3(\data_out_frame[20] [7]), .O(n21_adj_3960));
    defparam i8_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_adj_1006 (.I0(n15165), .I1(n35146), .I2(\data_out_frame[19] [7]), 
            .I3(GND_net), .O(n20_adj_3961));
    defparam i7_3_lut_adj_1006.LUT_INIT = 16'h6969;
    SB_LUT4 i11_4_lut_adj_1007 (.I0(n21_adj_3960), .I1(n16026), .I2(n18_adj_3958), 
            .I3(n35131), .O(n24_adj_3962));
    defparam i11_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_CARRY add_41_10 (.CI(n27928), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n27929));
    SB_LUT4 i12_4_lut_adj_1008 (.I0(n34985), .I1(n24_adj_3962), .I2(n20_adj_3961), 
            .I3(n15617), .O(n30998));
    defparam i12_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3963));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'heeee;
    SB_LUT4 i28681_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n34530), .I2(GND_net), 
            .I3(GND_net), .O(n35380));
    defparam i28681_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n17273));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3964));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_41_9_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n27927), .O(n2_adj_3965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_9 (.CI(n27927), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n27928));
    SB_LUT4 i33797_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n40561));   // verilog/coms.v(104[34:55])
    defparam i33797_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3966));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31430_4_lut (.I0(n19_adj_3964), .I1(\data_out_frame[22] [7]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38192));
    defparam i31430_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n17272));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i31431_3_lut (.I0(n43149), .I1(n38192), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38193));
    defparam i31431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31384_4_lut (.I0(n5_adj_3966), .I1(n40561), .I2(n101), .I3(byte_transmit_counter[0]), 
            .O(n38146));
    defparam i31384_4_lut.LUT_INIT = 16'haca0;
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n17399));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i31386_4_lut (.I0(n38146), .I1(n38193), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38148));
    defparam i31386_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31385_3_lut (.I0(n43161), .I1(n43155), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38147));
    defparam i31385_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n17398));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n17397));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n17271));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n17270));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12695_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n17377));
    defparam i12695_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_8_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n27926), .O(n2_adj_3967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3968));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_41_8 (.CI(n27926), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n27927));
    SB_LUT4 i33792_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n40556));   // verilog/coms.v(104[34:55])
    defparam i33792_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i12696_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n17378));
    defparam i12696_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_7_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n27925), .O(n2_adj_3969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_7 (.CI(n27925), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n27926));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3970));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31427_4_lut (.I0(n19_adj_3968), .I1(\data_out_frame[22] [6]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38189));
    defparam i31427_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31428_3_lut (.I0(n43143), .I1(n38189), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38190));
    defparam i31428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12697_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n17379));
    defparam i12697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31381_4_lut (.I0(n5_adj_3970), .I1(n40556), .I2(n101), .I3(byte_transmit_counter[0]), 
            .O(n38143));
    defparam i31381_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31383_4_lut (.I0(n38143), .I1(n38190), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38145));
    defparam i31383_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31382_3_lut (.I0(n43173), .I1(n43167), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38144));
    defparam i31382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_41_6_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n27924), .O(n2_adj_3971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3972));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40551));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3973));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_41_6 (.CI(n27924), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n27925));
    SB_LUT4 add_41_5_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n27923), .O(n2_adj_3974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i31424_4_lut (.I0(n19_adj_3972), .I1(\data_out_frame[22] [5]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38186));
    defparam i31424_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31425_3_lut (.I0(n43137), .I1(n38186), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38187));
    defparam i31425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12698_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n17380));
    defparam i12698_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31408_4_lut (.I0(n5_adj_3973), .I1(byte_transmit_counter[0]), 
            .I2(n101), .I3(n40551), .O(n38170));
    defparam i31408_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31410_4_lut (.I0(n38170), .I1(n38187), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38172));
    defparam i31410_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31409_3_lut (.I0(n43185), .I1(n43179), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38171));
    defparam i31409_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_41_5 (.CI(n27923), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n27924));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3975));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3976));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3977));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31421_4_lut (.I0(n19_adj_3975), .I1(\data_out_frame[22] [4]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38183));
    defparam i31421_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12699_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n17381));
    defparam i12699_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31422_3_lut (.I0(n43131), .I1(n38183), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38184));
    defparam i31422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31405_3_lut (.I0(n5_adj_3977), .I1(n6_adj_3976), .I2(n101), 
            .I3(GND_net), .O(n38167));
    defparam i31405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31407_4_lut (.I0(n38167), .I1(n38184), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38169));
    defparam i31407_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31406_3_lut (.I0(n43197), .I1(n43191), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38168));
    defparam i31406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3978));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_3_lut (.I0(\data_out_frame[5] [0]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40513));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3979));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3980));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3981));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3982));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31418_4_lut (.I0(n19_adj_3979), .I1(\data_out_frame[22] [3]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38180));
    defparam i31418_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31388_4_lut (.I0(n19_adj_3978), .I1(\data_out_frame[22] [0]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38150));
    defparam i31388_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31419_3_lut (.I0(n43125), .I1(n38180), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38181));
    defparam i31419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31402_3_lut (.I0(n5_adj_3981), .I1(n6_adj_3980), .I2(n101), 
            .I3(GND_net), .O(n38164));
    defparam i31402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31404_4_lut (.I0(n38164), .I1(n38181), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38166));
    defparam i31404_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12700_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34643), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n17382));
    defparam i12700_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31403_3_lut (.I0(n43209), .I1(n43203), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38165));
    defparam i31403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31389_3_lut (.I0(n43107), .I1(n38150), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38151));
    defparam i31389_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n17396));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i31393_4_lut (.I0(n5_adj_3982), .I1(byte_transmit_counter[0]), 
            .I2(n101), .I3(n40513), .O(n38155));
    defparam i31393_4_lut.LUT_INIT = 16'haca0;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n17395));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n17374));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i31395_4_lut (.I0(n38155), .I1(n38151), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38157));
    defparam i31395_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3983));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31394_3_lut (.I0(n43245), .I1(n43239), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38156));
    defparam i31394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n6_adj_3984));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha003;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3985));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31415_4_lut (.I0(n19_adj_3983), .I1(\data_out_frame[22] [2]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38177));
    defparam i31415_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31416_3_lut (.I0(n43119), .I1(n38177), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38178));
    defparam i31416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31399_3_lut (.I0(n5_adj_3985), .I1(n6_adj_3984), .I2(n101), 
            .I3(GND_net), .O(n38161));
    defparam i31399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31401_4_lut (.I0(n38161), .I1(n38178), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38163));
    defparam i31401_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31400_3_lut (.I0(n43221), .I1(n43215), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38162));
    defparam i31400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(\data_in_frame[0] [0]), 
            .I3(rx_data[0]), .O(n34101));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n17394));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n17269));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3986));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33773_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n40536));   // verilog/coms.v(104[34:55])
    defparam i33773_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3987));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31391_4_lut (.I0(n19_adj_3986), .I1(\data_out_frame[22] [1]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n38153));
    defparam i31391_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31392_3_lut (.I0(n43113), .I1(n38153), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38154));
    defparam i31392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31396_4_lut (.I0(n5_adj_3987), .I1(n40536), .I2(n101), .I3(byte_transmit_counter[0]), 
            .O(n38158));
    defparam i31396_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31398_4_lut (.I0(n38158), .I1(n38154), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n38160));
    defparam i31398_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31397_3_lut (.I0(n43233), .I1(n43227), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n38159));
    defparam i31397_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n17268));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_3279_9_lut (.I0(n4_adj_3988), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n27958), .O(n40164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n4368));   // verilog/coms.v(110[11:16])
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_4_lut_adj_1011 (.I0(\FRAME_MATCHER.state[3] ), .I1(n30171), 
            .I2(n4_adj_3963), .I3(n35380), .O(n37236));
    defparam i3_4_lut_adj_1011.LUT_INIT = 16'h0004;
    SB_LUT4 i12622_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n17304));
    defparam i12622_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1012 (.I0(n34673), .I1(n34521), .I2(n34671), 
            .I3(n6_adj_3989), .O(n34530));
    defparam i4_4_lut_adj_1012.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(n13231), .I1(n31_adj_3925), .I2(n31_adj_3946), 
            .I3(\FRAME_MATCHER.state [1]), .O(n29_adj_3951));   // verilog/coms.v(110[11:16])
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34675));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1016 (.I0(\data_in_frame[4] [2]), .I1(n34675), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[1] [6]), .O(n15798));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1017 (.I0(\data_in_frame[5] [4]), .I1(n34772), 
            .I2(\data_in_frame[3] [2]), .I3(GND_net), .O(n35054));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1017.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1018 (.I0(\data_in_frame[3] [7]), .I1(n34973), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[4] [1]), .O(n15794));   // verilog/coms.v(228[9:81])
    defparam i3_4_lut_adj_1018.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1019 (.I0(\FRAME_MATCHER.state[0] ), .I1(n36175), 
            .I2(n29_adj_3951), .I3(\FRAME_MATCHER.state [2]), .O(n7_c));
    defparam i1_4_lut_adj_1019.LUT_INIT = 16'h8ccc;
    SB_LUT4 add_41_4_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n27922), .O(n2_adj_3990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_4 (.CI(n27922), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n27923));
    SB_LUT4 i12623_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n17305));
    defparam i12623_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_41_3_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n27921), .O(n2_adj_3991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1020 (.I0(n24911), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n7_c), .I3(n139), .O(n8_adj_3992));
    defparam i3_4_lut_adj_1020.LUT_INIT = 16'h11b1;
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n17267));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_1021 (.I0(n3243), .I1(n8_adj_3992), .I2(n4368), 
            .I3(n4_adj_3993), .O(n43479));
    defparam i4_4_lut_adj_1021.LUT_INIT = 16'h0444;
    SB_LUT4 i33782_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state_31__N_2490 [3]), 
            .I2(n15448), .I3(n4_adj_3963), .O(n40215));   // verilog/coms.v(126[12] 289[6])
    defparam i33782_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_CARRY add_41_3 (.CI(n27921), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n27922));
    SB_LUT4 add_3279_8_lut (.I0(\FRAME_MATCHER.i_31__N_2389 ), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n27957), .O(n40163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1022 (.I0(\data_in_frame[1] [2]), .I1(n35054), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n15939));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1022.LUT_INIT = 16'h9696;
    SB_LUT4 i12624_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n17306));
    defparam i12624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12626_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n17308));
    defparam i12626_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_3279_8 (.CI(n27957), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n27958));
    SB_LUT4 add_41_2_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_2_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n17266));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n17265));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n27921));
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n17264));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n17263));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n17262));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n17261));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n17260));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n17259));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n17258));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n17257));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n17256));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n17255));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12627_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n17309));
    defparam i12627_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i22317_3_lut (.I0(byte_transmit_counter[7]), .I1(n40164), .I2(n24117), 
            .I3(GND_net), .O(n17630));
    defparam i22317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22311_3_lut (.I0(byte_transmit_counter[6]), .I1(n40163), .I2(n24117), 
            .I3(GND_net), .O(n17629));
    defparam i22311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n139));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(\FRAME_MATCHER.state[0] ), .I1(n15448), 
            .I2(GND_net), .I3(GND_net), .O(n34657));   // verilog/coms.v(193[5:24])
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1025 (.I0(n18962), .I1(n34657), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(GND_net), .O(n63));   // verilog/coms.v(193[5:24])
    defparam i2_3_lut_adj_1025.LUT_INIT = 16'hefef;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(n34858), .I3(GND_net), .O(n30555));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1026 (.I0(n13978), .I1(n35109), .I2(n34803), 
            .I3(\data_in_frame[1] [1]), .O(n10_adj_3994));   // verilog/coms.v(68[16:27])
    defparam i4_4_lut_adj_1026.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1027 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[2] [6]), .I3(n15780), .O(n13));   // verilog/coms.v(69[16:69])
    defparam i5_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n17254));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n17253));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n17252));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n17251));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n17250));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n17249));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n17248));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n17247));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n17246));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n17245));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_3279_7_lut (.I0(\FRAME_MATCHER.i_31__N_2389 ), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n27956), .O(n40162)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_7_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n17244));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n17243));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n17242));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n17241));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n17240));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n17239));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n17238));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n17237));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n17236));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n17235));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n17234));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n17233));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n17232));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n17231));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n17230));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n17229));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n17228));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n17227));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n17226));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n17225));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n17224));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n17223));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n17222));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n17221));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12628_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n17310));
    defparam i12628_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n17220));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n17219));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n17218));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n17217));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n17216));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n17215));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n17214));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n17213));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n17212));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n17211));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n17210));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n17209));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n17208));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n17207));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n17206));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n17205));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n17204));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n17203));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n17202));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n17201));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n17200));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n17199));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n17198));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n17197));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n17196));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n17195));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n17194));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n17193));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n17192));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n17191));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i22303_3_lut (.I0(byte_transmit_counter[5]), .I1(n40162), .I2(n24117), 
            .I3(GND_net), .O(n16927));
    defparam i22303_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_4_lut_adj_1028 (.I0(n4_adj_3995), .I1(n34845), .I2(n16104), 
            .I3(\data_in_frame[3] [0]), .O(n12_adj_3996));   // verilog/coms.v(69[16:69])
    defparam i5_4_lut_adj_1028.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1029 (.I0(\data_in_frame[3] [3]), .I1(n12_adj_3996), 
            .I2(n35109), .I3(n16160), .O(Kp_23__N_896));   // verilog/coms.v(69[16:69])
    defparam i6_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n34731));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1031 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[5] [7]), .O(n34829));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\data_in_frame[3] [5]), .I1(n34829), 
            .I2(GND_net), .I3(GND_net), .O(n16289));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1033 (.I0(\data_in_frame[4] [7]), .I1(Kp_23__N_896), 
            .I2(GND_net), .I3(GND_net), .O(n16232));
    defparam i1_2_lut_adj_1033.LUT_INIT = 16'h6666;
    SB_LUT4 equal_1174_i15_2_lut (.I0(Kp_23__N_893), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3943));   // verilog/coms.v(228[9:81])
    defparam equal_1174_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i17953_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34647), .I2(\data_in_frame[0] [4]), 
            .I3(rx_data[4]), .O(n17307));
    defparam i17953_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n17190));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_3279_7 (.CI(n27956), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n27957));
    SB_LUT4 add_3279_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n27955), .O(n7813[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n17189));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n17188));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n17187));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n17186));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n17185));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n17184));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n17183));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n17182));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n17181));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n17180));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n17179));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n17178));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n17177));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n17176));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n17175));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n17174));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_1034 (.I0(n34772), .I1(n4_c), .I2(\data_in_frame[3] [0]), 
            .I3(GND_net), .O(n34858));   // verilog/coms.v(69[16:69])
    defparam i2_3_lut_adj_1034.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n17173));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 Kp_23__N_858_I_0_2_lut (.I0(Kp_23__N_858), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_926));   // verilog/coms.v(69[16:69])
    defparam Kp_23__N_858_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n17172));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n17171));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n17170));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n17169));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n17165));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n17164));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n17163));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n17162));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n17161));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n17160));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n17159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n17158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n17157));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n17156));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2][6] ), .C(clk32MHz), .D(n17155));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12723_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n17405));
    defparam i12723_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i22 (.Q(\data_in[2][5] ), .C(clk32MHz), .D(n17154));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2][4] ), .C(clk32MHz), .D(n17153));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2][3] ), .C(clk32MHz), .D(n22677));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2][2] ), .C(clk32MHz), .D(n17151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2][1] ), .C(clk32MHz), .D(n17150));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12724_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n17406));
    defparam i12724_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i17 (.Q(\data_in[2][0] ), .C(clk32MHz), .D(n17149));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n17148));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1][6] ), .C(clk32MHz), .D(n17147));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state_31__N_2490 [3]), 
            .I2(n12859), .I3(n34530), .O(n13195));   // verilog/coms.v(126[12] 289[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i2_2_lut_adj_1035 (.I0(\data_in[2][3] ), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3997));
    defparam i2_2_lut_adj_1035.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1036 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0]_c [7]), .O(n14_adj_3998));
    defparam i6_4_lut_adj_1036.LUT_INIT = 16'hfeff;
    SB_DFF data_in_0___i14 (.Q(\data_in[1][5] ), .C(clk32MHz), .D(n17146));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut_adj_1037 (.I0(\data_in[3] [6]), .I1(n14_adj_3998), 
            .I2(n10_adj_3997), .I3(\data_in[2][1] ), .O(n15514));
    defparam i7_4_lut_adj_1037.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(n15329), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3999));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'heeee;
    SB_LUT4 i19405_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3999), .I3(\FRAME_MATCHER.i [1]), .O(n737));   // verilog/coms.v(154[9:60])
    defparam i19405_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i12717_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n17399));
    defparam i12717_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1039 (.I0(n15342), .I1(n15514), .I2(\data_in[1][3] ), 
            .I3(\data_in[0][5] ), .O(n20_adj_4000));
    defparam i8_4_lut_adj_1039.LUT_INIT = 16'hefff;
    SB_LUT4 i7_4_lut_adj_1040 (.I0(\data_in[2][5] ), .I1(\data_in[1][6] ), 
            .I2(\data_in[3] [7]), .I3(\data_in[2][6] ), .O(n19_adj_4001));
    defparam i7_4_lut_adj_1040.LUT_INIT = 16'hfffd;
    SB_LUT4 i31373_4_lut (.I0(\data_in[2][0] ), .I1(\data_in[1][2] ), .I2(\data_in[3] [2]), 
            .I3(\data_in[0][1] ), .O(n38076));
    defparam i31373_4_lut.LUT_INIT = 16'h8000;
    SB_DFF data_in_0___i13 (.Q(\data_in[1][4] ), .C(clk32MHz), .D(n17145));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1][3] ), .C(clk32MHz), .D(n17144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1][2] ), .C(clk32MHz), .D(n17143));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i11_3_lut (.I0(n38076), .I1(n19_adj_4001), .I2(n20_adj_4000), 
            .I3(GND_net), .O(n63_adj_4002));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i4_4_lut_adj_1041 (.I0(\data_in[1] [7]), .I1(\data_in[0][0] ), 
            .I2(\data_in[1][1] ), .I3(\data_in[0][4] ), .O(n10_adj_4003));
    defparam i4_4_lut_adj_1041.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1042 (.I0(\data_in[3] [4]), .I1(n10_adj_4003), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n15552));
    defparam i5_3_lut_adj_1042.LUT_INIT = 16'hdfdf;
    SB_CARRY add_3279_6 (.CI(n27955), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n27956));
    SB_LUT4 i5_3_lut_adj_1043 (.I0(\data_in[0][3] ), .I1(\data_in[1][4] ), 
            .I2(\data_in[1][5] ), .I3(GND_net), .O(n14_adj_4004));
    defparam i5_3_lut_adj_1043.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1044 (.I0(\data_in[0][6] ), .I1(n15552), .I2(\data_in[2][4] ), 
            .I3(\data_in[1][0] ), .O(n15_adj_4005));
    defparam i6_4_lut_adj_1044.LUT_INIT = 16'hfeff;
    SB_DFF data_in_0___i10 (.Q(\data_in[1][1] ), .C(clk32MHz), .D(n17142));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1][0] ), .C(clk32MHz), .D(n17141));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0]_c [7]), .C(clk32MHz), .D(n17140));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0][6] ), .C(clk32MHz), .D(n17139));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i8_4_lut_adj_1045 (.I0(n15_adj_4005), .I1(\data_in[3] [0]), 
            .I2(n14_adj_4004), .I3(\data_in[2][2] ), .O(n15342));
    defparam i8_4_lut_adj_1045.LUT_INIT = 16'hfbff;
    SB_DFF data_in_0___i6 (.Q(\data_in[0][5] ), .C(clk32MHz), .D(n17138));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_3279_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n27954), .O(n7813[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1046 (.I0(\data_in[1][2] ), .I1(\data_in[1][6] ), 
            .I2(\data_in[2][0] ), .I3(\data_in[2][5] ), .O(n16_adj_4006));
    defparam i6_4_lut_adj_1046.LUT_INIT = 16'hfffb;
    SB_LUT4 i7_4_lut_adj_1047 (.I0(\data_in[2][6] ), .I1(\data_in[3] [2]), 
            .I2(\data_in[0][1] ), .I3(\data_in[0][5] ), .O(n17_adj_4007));
    defparam i7_4_lut_adj_1047.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1048 (.I0(n17_adj_4007), .I1(\data_in[1][3] ), 
            .I2(n16_adj_4006), .I3(\data_in[3] [7]), .O(n15445));
    defparam i9_4_lut_adj_1048.LUT_INIT = 16'hfeff;
    SB_LUT4 i12718_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n17400));
    defparam i12718_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1049 (.I0(n15445), .I1(\data_in[0]_c [7]), .I2(\data_in[3] [3]), 
            .I3(n15342), .O(n16_adj_4008));
    defparam i6_4_lut_adj_1049.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1050 (.I0(\data_in[3] [6]), .I1(\data_in[0] [2]), 
            .I2(\data_in[2][3] ), .I3(\data_in[2][1] ), .O(n17_adj_4009));
    defparam i7_4_lut_adj_1050.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_3_lut_adj_1051 (.I0(\FRAME_MATCHER.i_31__N_2390 ), .I1(n2855), 
            .I2(n10283), .I3(GND_net), .O(n31_adj_4010));   // verilog/coms.v(113[11:12])
    defparam i1_3_lut_adj_1051.LUT_INIT = 16'h2020;
    SB_DFF data_in_0___i5 (.Q(\data_in[0][4] ), .C(clk32MHz), .D(n17137));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0][3] ), .C(clk32MHz), .D(n17136));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_1052 (.I0(n17_adj_4009), .I1(\data_in[3] [5]), 
            .I2(n16_adj_4008), .I3(\data_in[3] [1]), .O(n63_adj_4011));
    defparam i9_4_lut_adj_1052.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1053 (.I0(\data_in[2][4] ), .I1(\data_in[0][3] ), 
            .I2(\data_in[1][5] ), .I3(n15552), .O(n18_adj_4012));
    defparam i7_4_lut_adj_1053.LUT_INIT = 16'hfffd;
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n17135));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_1054 (.I0(\data_in[0][6] ), .I1(n18_adj_4012), 
            .I2(\data_in[2][2] ), .I3(n15445), .O(n20_adj_4013));
    defparam i9_4_lut_adj_1054.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1][0] ), .I1(\data_in[3] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4014));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1055 (.I0(n15_adj_4014), .I1(n20_adj_4013), .I2(n15514), 
            .I3(\data_in[1][4] ), .O(n22667));
    defparam i10_4_lut_adj_1055.LUT_INIT = 16'hfeff;
    SB_LUT4 i55_3_lut (.I0(\FRAME_MATCHER.i_31__N_2386 ), .I1(n737), .I2(n10283), 
            .I3(GND_net), .O(n41_adj_4015));   // verilog/coms.v(113[11:12])
    defparam i55_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_3_lut_adj_1056 (.I0(\FRAME_MATCHER.state [2]), .I1(n22667), 
            .I2(n63_adj_4011), .I3(GND_net), .O(n122));
    defparam i1_3_lut_adj_1056.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_3_lut_adj_1057 (.I0(\FRAME_MATCHER.i_31__N_2392 ), .I1(n10283), 
            .I2(n3741), .I3(GND_net), .O(n42));   // verilog/coms.v(113[11:12])
    defparam i1_3_lut_adj_1057.LUT_INIT = 16'h0808;
    SB_LUT4 i57_2_lut (.I0(n10283), .I1(n2720), .I2(GND_net), .I3(GND_net), 
            .O(n43));
    defparam i57_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_0___i2 (.Q(\data_in[0][1] ), .C(clk32MHz), .D(n17134));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n17133));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n17132));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n17131));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n17130));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n17129));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4246_2_lut (.I0(n63_adj_4002), .I1(n737), .I2(GND_net), .I3(GND_net), 
            .O(n8849));   // verilog/coms.v(154[6] 156[9])
    defparam i4246_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(n41_adj_4015), .I1(n31_adj_4010), .I2(GND_net), 
            .I3(GND_net), .O(n34668));
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'heeee;
    SB_CARRY add_3279_5 (.CI(n27954), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n27955));
    SB_LUT4 i1_3_lut_adj_1059 (.I0(n1205), .I1(\FRAME_MATCHER.i_31__N_2389 ), 
            .I2(n10283), .I3(GND_net), .O(n17_adj_4016));   // verilog/coms.v(113[11:12])
    defparam i1_3_lut_adj_1059.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_adj_1060 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n26928), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2390 ));   // verilog/coms.v(126[12] 289[6])
    defparam i2_3_lut_adj_1060.LUT_INIT = 16'h4040;
    SB_LUT4 i20_4_lut_adj_1061 (.I0(n40215), .I1(n17_adj_4016), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(n34668), .O(n34051));
    defparam i20_4_lut_adj_1061.LUT_INIT = 16'hfaca;
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n17128));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n17127));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n17126));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n17125));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n17124));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n17123));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i17_4_lut_adj_1062 (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_4017));
    defparam i17_4_lut_adj_1062.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1063 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [15]), .I3(\FRAME_MATCHER.i [16]), .O(n40));
    defparam i15_4_lut_adj_1063.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1064 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [30]), .O(n41_adj_4018));
    defparam i16_4_lut_adj_1064.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1065 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [25]), .O(n39_adj_4019));
    defparam i14_4_lut_adj_1065.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n38_adj_4020));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4021));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23_4_lut (.I0(n39_adj_4019), .I1(n41_adj_4018), .I2(n40), 
            .I3(n42_adj_4017), .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [27]), .O(n43_adj_4022));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n43_adj_4022), .I1(n48), .I2(n37_adj_4021), 
            .I3(n38_adj_4020), .O(n15540));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12719_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n17401));
    defparam i12719_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19408_4_lut (.I0(n10_adj_4023), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n15540), .O(n3741));   // verilog/coms.v(248[9:58])
    defparam i19408_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i12720_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n17402));
    defparam i12720_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n17122));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n17121));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n17120));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n17119));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n17118));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1066 (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/coms.v(100[12:33])
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h8888;
    SB_LUT4 i36287_4_lut (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[5]), 
            .I2(n84), .I3(byte_transmit_counter[6]), .O(tx_transmit_N_3220));
    defparam i36287_4_lut.LUT_INIT = 16'h0001;
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n17117));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n17116));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut_adj_1067 (.I0(n15437), .I1(n42349), .I2(n2030), .I3(n34657), 
            .O(n2720));
    defparam i2_4_lut_adj_1067.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_3_lut_adj_1068 (.I0(n2720), .I1(n1205), .I2(\FRAME_MATCHER.i_31__N_2389 ), 
            .I3(GND_net), .O(n4));
    defparam i1_3_lut_adj_1068.LUT_INIT = 16'heaea;
    SB_LUT4 select_365_Select_2_i7_3_lut (.I0(\FRAME_MATCHER.state_31__N_2426[2] ), 
            .I1(\FRAME_MATCHER.i_31__N_2392 ), .I2(n3741), .I3(GND_net), 
            .O(n7));
    defparam select_365_Select_2_i7_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n17115));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n17114));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n17113));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 select_365_Select_1_i5_4_lut (.I0(n63_adj_4002), .I1(\FRAME_MATCHER.i_31__N_2390 ), 
            .I2(n2855), .I3(n92[1]), .O(n5_adj_4026));
    defparam select_365_Select_1_i5_4_lut.LUT_INIT = 16'hccc4;
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n17112));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n17111));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n17110));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n17109));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12721_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n17403));
    defparam i12721_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n17108));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12722_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34631), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n17404));
    defparam i12722_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1069 (.I0(n63), .I1(n30072), .I2(n1), .I3(n5_adj_4026), 
            .O(n43474));
    defparam i3_4_lut_adj_1069.LUT_INIT = 16'hfffd;
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n17107));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n17106));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n17105));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n17104));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n17103));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n17102));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n17101));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n17100));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n17099));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n17098));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n17097));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n17096));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n17095));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n17094));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n17093));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1070 (.I0(n34931), .I1(n35143), .I2(GND_net), 
            .I3(GND_net), .O(n35144));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n17092));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n17091));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n17090));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n17089));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n17088));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n17087));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n17086));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n17085));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n17084));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_1071 (.I0(\data_out_frame[19] [5]), .I1(n34957), 
            .I2(\data_out_frame[19] [4]), .I3(n30653), .O(n36946));
    defparam i3_4_lut_adj_1071.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(n30523), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n30603));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1073 (.I0(\data_out_frame[17] [1]), .I1(n15617), 
            .I2(n35198), .I3(n6_adj_4027), .O(n36900));
    defparam i4_4_lut_adj_1073.LUT_INIT = 16'h9669;
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n17083));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n17082));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n17081));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n17080));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n17079));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n17078));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n17077));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n17076));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n17075));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n17074));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_1074 (.I0(\data_out_frame[17] [2]), .I1(n35066), 
            .I2(n1593), .I3(n35261), .O(n16_adj_4028));
    defparam i6_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1075 (.I0(n34970), .I1(n35214), .I2(n15171), 
            .I3(n35034), .O(n17_adj_4029));
    defparam i7_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1076 (.I0(n17_adj_4029), .I1(n1504), .I2(n16_adj_4028), 
            .I3(n1667), .O(n30653));
    defparam i9_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(n30653), .I1(n35134), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4030));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [2]), 
            .I2(n1829), .I3(n6_adj_4030), .O(n36211));
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35034));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1080 (.I0(n35279), .I1(n34912), .I2(n35255), 
            .I3(n30611), .O(n14_adj_4031));
    defparam i6_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1081 (.I0(n9_adj_4032), .I1(n14_adj_4031), .I2(n35276), 
            .I3(n31275), .O(n35804));
    defparam i7_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1082 (.I0(n34905), .I1(n35151), .I2(\data_out_frame[19] [1]), 
            .I3(n31275), .O(n12_adj_4033));
    defparam i5_4_lut_adj_1082.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1083 (.I0(\data_out_frame[16] [6]), .I1(n12_adj_4033), 
            .I2(n35234), .I3(n15165), .O(n36587));
    defparam i6_4_lut_adj_1083.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1084 (.I0(\data_out_frame[20] [7]), .I1(n35166), 
            .I2(n34976), .I3(n15986), .O(n36281));
    defparam i3_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1085 (.I0(n31_adj_3925), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4034));   // verilog/coms.v(126[12] 289[6])
    defparam i2_2_lut_adj_1085.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1086 (.I0(n7_adj_4034), .I1(n18939), .I2(n13231), 
            .I3(\FRAME_MATCHER.state [2]), .O(n36885));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1086.LUT_INIT = 16'hfeff;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38148), .I3(n38147), .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38145), .I3(n38144), .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38172), .I3(n38171), .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38169), .I3(n38168), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38166), .I3(n38165), .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38163), .I3(n38162), .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 mux_1046_i8_3_lut (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4291), .I3(GND_net), .O(n4299));
    defparam mux_1046_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1087 (.I0(\FRAME_MATCHER.state [11]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(\FRAME_MATCHER.state [9]), .I3(\FRAME_MATCHER.state [10]), 
            .O(n10_adj_4035));
    defparam i4_4_lut_adj_1087.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1088 (.I0(\FRAME_MATCHER.state [15]), .I1(n10_adj_4035), 
            .I2(\FRAME_MATCHER.state [8]), .I3(GND_net), .O(n34673));
    defparam i5_3_lut_adj_1088.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut_adj_1089 (.I0(\FRAME_MATCHER.state [17]), .I1(\FRAME_MATCHER.state [31]), 
            .I2(\FRAME_MATCHER.state [27]), .I3(GND_net), .O(n14_adj_4036));
    defparam i5_3_lut_adj_1089.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1090 (.I0(\FRAME_MATCHER.state [23]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [25]), .I3(\FRAME_MATCHER.state [22]), 
            .O(n15_adj_4037));
    defparam i6_4_lut_adj_1090.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1091 (.I0(n15_adj_4037), .I1(\FRAME_MATCHER.state [26]), 
            .I2(n14_adj_4036), .I3(\FRAME_MATCHER.state [28]), .O(n34523));
    defparam i8_4_lut_adj_1091.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1092 (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n34671));
    defparam i3_4_lut_adj_1092.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1093 (.I0(\FRAME_MATCHER.state [24]), .I1(\FRAME_MATCHER.state [19]), 
            .I2(\FRAME_MATCHER.state [20]), .I3(GND_net), .O(n8_adj_4038));
    defparam i3_3_lut_adj_1093.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_adj_1094 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [18]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4039));
    defparam i2_2_lut_adj_1094.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1095 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(n7_adj_4039), .I3(n8_adj_4038), .O(n34521));   // verilog/coms.v(126[12] 289[6])
    defparam i2_4_lut_adj_1095.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1096 (.I0(n34521), .I1(n34671), .I2(n34523), 
            .I3(n6_adj_4040), .O(n15448));
    defparam i4_4_lut_adj_1096.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n18962));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38157), .I3(n38156), .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 mux_1046_i7_3_lut (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4291), .I3(GND_net), .O(n4298));
    defparam mux_1046_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n38160), .I3(n38159), .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i12260_4_lut_4_lut (.I0(n24117), .I1(\FRAME_MATCHER.i_31__N_2389 ), 
            .I2(n7813[3]), .I3(byte_transmit_counter[3]), .O(n16942));
    defparam i12260_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 mux_1046_i18_3_lut (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4291), .I3(GND_net), .O(n4309));
    defparam mux_1046_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12248_4_lut_4_lut (.I0(n24117), .I1(\FRAME_MATCHER.i_31__N_2389 ), 
            .I2(n7813[4]), .I3(byte_transmit_counter[4]), .O(n16930));
    defparam i12248_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 i12317_4_lut_4_lut (.I0(n24117), .I1(\FRAME_MATCHER.i_31__N_2389 ), 
            .I2(n7813[1]), .I3(byte_transmit_counter[1]), .O(n16999));
    defparam i12317_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_LUT4 mux_1046_i17_3_lut (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4291), .I3(GND_net), .O(n4308));
    defparam mux_1046_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3279_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n27953), .O(n7813[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3279_4 (.CI(n27953), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n27954));
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3991), .S(n3_adj_4041));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n17353));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_3279_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n27952), .O(n7813[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3279_3 (.CI(n27952), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n27953));
    SB_LUT4 add_3279_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3220), .I3(GND_net), .O(n7813[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3279_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3279_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3220), 
            .CO(n27952));
    SB_LUT4 i12314_4_lut_4_lut (.I0(n24117), .I1(\FRAME_MATCHER.i_31__N_2389 ), 
            .I2(n7813[2]), .I3(byte_transmit_counter[2]), .O(n16996));
    defparam i12314_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n17373));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n17372));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_33_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n27951), .O(n2_adj_4042)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_33_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n17371));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n17370));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n17369));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3990), .S(n3_adj_4043));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3974), .S(n3_adj_4044));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3971), .S(n3_adj_4045));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3969), .S(n3_adj_4046));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3967), .S(n3_adj_4047));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3965), .S(n3_adj_4048));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3959), .S(n3_adj_4049));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3953), .S(n3_adj_4050));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3948), .S(n3_adj_4051));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3940), .S(n3_adj_4052));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3932), .S(n3_adj_4053));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3929), .S(n3_adj_4054));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3923), .S(n3_adj_4055));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3906), .S(n3_adj_4056));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3900), .S(n3_adj_4057));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_3899), .S(n3_adj_4058));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3898), .S(n3_adj_4059));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4060), .S(n3_adj_4061));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4062), .S(n3_adj_4063));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4064), .S(n3_adj_4065));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4066), .S(n3_adj_4067));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4068), .S(n3_adj_4069));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4070), .S(n3_adj_4071));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4072), .S(n3_adj_4073));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4074), .S(n3_adj_4075));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4076), .S(n3_adj_4077));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4078), .S(n3_adj_4079));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4080), .S(n3_adj_4081));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4082), .S(n3_adj_4083));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4042), .S(n3_adj_4084));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n16593), .D(n36281));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_1046_i16_3_lut (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4291), .I3(GND_net), .O(n4307));
    defparam mux_1046_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n16593), .D(n36199));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n16593), .D(n36587));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n16593), .D(n35804));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n16593), .D(n36211));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n16593), .D(n36900));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n16593), .D(n36946));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n16593), .D(n36969));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n16593), .D(n30998));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n16593), .D(n34990));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n16593), .D(n35232));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n16593), .D(n35126));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n16593), .D(n35146));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n16593), .D(n35144));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n16593), .D(n34910));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n33967), .S(n43474));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n33969), .S(n34051));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n34111), .S(n33977));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n34113), .S(n34043));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n7_adj_4085), .S(n8_adj_4086));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n34115), .S(n34041));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n34117), .S(n34039));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n7_adj_4087), .S(n8_adj_4088));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n34119), .S(n34037));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n34121), .S(n8_adj_4089));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n34123), .S(n34035));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n34125), .S(n34033));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n34127), .S(n34031));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n34129), .S(n34029));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n7_adj_4090), .S(n8_adj_4091));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n34131), .S(n8_adj_4092));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n7_adj_4093), .S(n8_adj_4094));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n23956), .S(n24611));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n7_adj_4095), .S(n8_adj_4096));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n34133), .S(n34027));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n34135), .S(n34025));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n34137), .S(n34023));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n34139), .S(n8_adj_4097));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n34141), .S(n34021));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n34143), .S(n34019));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n34145), .S(n34017));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n7_adj_4098), .S(n8_adj_4099));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n34147), .S(n34015));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n34149), .S(n34013));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_4100), .S(n8_adj_4101));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_32_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n27950), .O(n2_adj_4082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_1098 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[12] [6]), .I3(\data_in_frame[12] [7]), .O(n34848));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[6] [3]), .I3(GND_net), .O(n35226));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [0]), 
            .I2(n10_adj_4102), .I3(n15871), .O(n35240));   // verilog/coms.v(83[17:28])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n17368));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12350_4_lut_4_lut (.I0(n24117), .I1(\FRAME_MATCHER.i_31__N_2389 ), 
            .I2(n7813[0]), .I3(byte_transmit_counter[0]), .O(n17032));
    defparam i12350_4_lut_4_lut.LUT_INIT = 16'hea40;
    SB_CARRY add_41_32 (.CI(n27950), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n27951));
    SB_LUT4 mux_1046_i20_3_lut (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4291), .I3(GND_net), .O(n4311));
    defparam mux_1046_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_41_31_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n27949), .O(n2_adj_4080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_24 (.CI(n27942), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n27943));
    SB_DFFESR LED_3208 (.Q(LED_c), .C(clk32MHz), .E(n43479), .D(n16737), 
            .R(n37236));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_1099 (.I0(\data_in_frame[5] [3]), .I1(n34864), 
            .I2(Kp_23__N_926), .I3(n13978), .O(n15944));
    defparam i3_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_CARRY add_41_31 (.CI(n27949), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n27950));
    SB_LUT4 i1_2_lut_adj_1100 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n12905));
    defparam i1_2_lut_adj_1100.LUT_INIT = 16'heeee;
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n17367));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n17366));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_1046_i19_3_lut (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4291), .I3(GND_net), .O(n4310));
    defparam mux_1046_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_41_30_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n27948), .O(n2_adj_4078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_30_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n17365));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n17421));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n17420));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_30 (.CI(n27948), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n27949));
    SB_LUT4 add_41_29_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n27947), .O(n2_adj_4076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_29 (.CI(n27947), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n27948));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n43242));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n43242_bdd_4_lut (.I0(n43242), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n43245));
    defparam n43242_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36457 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n43236));
    defparam byte_transmit_counter_0__bdd_4_lut_36457.LUT_INIT = 16'he4aa;
    SB_LUT4 n43236_bdd_4_lut (.I0(n43236), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n43239));
    defparam n43236_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36452 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n43230));
    defparam byte_transmit_counter_0__bdd_4_lut_36452.LUT_INIT = 16'he4aa;
    SB_LUT4 n43230_bdd_4_lut (.I0(n43230), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n43233));
    defparam n43230_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36447 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n43224));
    defparam byte_transmit_counter_0__bdd_4_lut_36447.LUT_INIT = 16'he4aa;
    SB_LUT4 n43224_bdd_4_lut (.I0(n43224), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n43227));
    defparam n43224_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36442 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n43218));
    defparam byte_transmit_counter_0__bdd_4_lut_36442.LUT_INIT = 16'he4aa;
    SB_LUT4 n43218_bdd_4_lut (.I0(n43218), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n43221));
    defparam n43218_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36437 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n43212));
    defparam byte_transmit_counter_0__bdd_4_lut_36437.LUT_INIT = 16'he4aa;
    SB_LUT4 add_41_28_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n27946), .O(n2_adj_4074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_28_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n17419));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n17418));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n17417));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n17416));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n17415));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_1046_i22_3_lut (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4291), .I3(GND_net), .O(n4313));
    defparam mux_1046_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1046_i21_3_lut (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4291), .I3(GND_net), .O(n4312));
    defparam mux_1046_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1046_i24_3_lut (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4291), .I3(GND_net), .O(n4315));
    defparam mux_1046_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20251_2_lut (.I0(n24524), .I1(n34530), .I2(GND_net), .I3(GND_net), 
            .O(n24911));
    defparam i20251_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[8] [3]), .I1(n15657), .I2(n16289), 
            .I3(\data_in_frame[12] [7]), .O(n35285));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 n43212_bdd_4_lut (.I0(n43212), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n43215));
    defparam n43212_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_41_28 (.CI(n27946), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n27947));
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n17414));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n17413));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n17412));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n17411));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n17410));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n17364));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n17363));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n17362));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_41_27_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n27945), .O(n2_adj_4072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_27_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n17361));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n17393));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_41_27 (.CI(n27945), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n27946));
    SB_LUT4 add_41_26_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n27944), .O(n2_adj_4070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1101 (.I0(\data_in_frame[8] [3]), .I1(n15657), 
            .I2(n16289), .I3(\data_in_frame[19] [6]), .O(n6_adj_4103));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1102 (.I0(\data_in_frame[4] [3]), .I1(n34763), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[2] [1]), .O(n16137));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_CARRY add_41_26 (.CI(n27944), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n27945));
    SB_LUT4 add_41_25_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n27943), .O(n2_adj_4068)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_25 (.CI(n27943), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n27944));
    SB_LUT4 add_41_24_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n27942), .O(n2_adj_4066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_22 (.CI(n27940), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n27941));
    SB_LUT4 add_41_23_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n27941), .O(n2_adj_4064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_23 (.CI(n27941), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n27942));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36432 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n43206));
    defparam byte_transmit_counter_0__bdd_4_lut_36432.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n17352));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n43206_bdd_4_lut (.I0(n43206), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n43209));
    defparam n43206_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i35596_2_lut (.I0(n30171), .I1(n34530), .I2(GND_net), .I3(GND_net), 
            .O(n3243));
    defparam i35596_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i18035_3_lut (.I0(\data_in[0]_c [7]), .I1(\data_in[1] [7]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n17140));   // verilog/coms.v(88[7:20])
    defparam i18035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1103 (.I0(n121), .I1(n84), .I2(byte_transmit_counter[5]), 
            .I3(byte_transmit_counter[6]), .O(n10_adj_4104));
    defparam i4_4_lut_adj_1103.LUT_INIT = 16'h0002;
    SB_LUT4 mux_1046_i23_3_lut (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4291), .I3(GND_net), .O(n4314));
    defparam mux_1046_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1104 (.I0(n30998), .I1(n34988), .I2(n30603), 
            .I3(n34985), .O(n36969));
    defparam i2_3_lut_4_lut_adj_1104.LUT_INIT = 16'h9669;
    SB_LUT4 i18032_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17148));   // verilog/coms.v(88[7:20])
    defparam i18032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18034_3_lut (.I0(\data_in[2][1] ), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17150));   // verilog/coms.v(88[7:20])
    defparam i18034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18014_3_lut (.I0(\data_in[2][3] ), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22677));   // verilog/coms.v(88[7:20])
    defparam i18014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18033_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17156));   // verilog/coms.v(88[7:20])
    defparam i18033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut_adj_1105 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[10] [2]), 
            .I2(n15944), .I3(n10_adj_4105), .O(n30585));   // verilog/coms.v(83[17:28])
    defparam i5_3_lut_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i12614_3_lut_4_lut (.I0(n30998), .I1(n34988), .I2(n16593), 
            .I3(\data_out_frame[22] [0]), .O(n17296));
    defparam i12614_3_lut_4_lut.LUT_INIT = 16'h6f60;
    SB_LUT4 mux_757_i1_4_lut (.I0(n37977), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n24911), .I3(n10_adj_4104), .O(n3241[0]));   // verilog/coms.v(144[4] 288[11])
    defparam mux_757_i1_4_lut.LUT_INIT = 16'h5c0c;
    SB_LUT4 i2_3_lut_4_lut_adj_1106 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[10] [2]), 
            .I2(n15756), .I3(n35282), .O(n35243));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n17360));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n17359));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n16104));   // verilog/coms.v(73[16:43])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[0] [4]), .O(Kp_23__N_893));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_22_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n27940), .O(n2_adj_4062)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_22_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n17358));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n17357));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n17356));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36427 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n43200));
    defparam byte_transmit_counter_0__bdd_4_lut_36427.LUT_INIT = 16'he4aa;
    SB_LUT4 n43200_bdd_4_lut (.I0(n43200), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n43203));
    defparam n43200_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16160));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3995));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n16832));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_858), 
            .I2(GND_net), .I3(GND_net), .O(n34845));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n17334));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1110 (.I0(n34816), .I1(n35081), .I2(\data_out_frame[14] [6]), 
            .I3(n31249), .O(n34970));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1111 (.I0(n34816), .I1(n35081), .I2(n30611), 
            .I3(GND_net), .O(n31226));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1111.LUT_INIT = 16'h9696;
    SB_LUT4 add_41_21_lut (.I0(n2030), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n27939), .O(n2_adj_4060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_1112 (.I0(n34816), .I1(n35081), .I2(n34851), 
            .I3(n16110), .O(n35115));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1113 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n16353));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut_adj_1113.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1114 (.I0(n34789), .I1(n35066), .I2(\data_out_frame[19] [7]), 
            .I3(\data_out_frame[17] [6]), .O(n30619));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i31281_3_lut_4_lut (.I0(\data_in_frame[2] [3]), .I1(n34693), 
            .I2(n4_adj_3995), .I3(\data_in_frame[0] [6]), .O(n37983));   // verilog/coms.v(163[9:87])
    defparam i31281_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i12710_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n17392));
    defparam i12710_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1115 (.I0(\data_in_frame[2] [3]), .I1(n34693), 
            .I2(\data_in_frame[4] [5]), .I3(n16104), .O(n16142));   // verilog/coms.v(163[9:87])
    defparam i2_3_lut_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i12711_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n17393));
    defparam i12711_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12725_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n17407));
    defparam i12725_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12726_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n17408));
    defparam i12726_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n16986));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12727_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n17409));
    defparam i12727_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n17409));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n17408));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n17407));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n17406));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12728_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n17410));
    defparam i12728_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12729_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n17411));
    defparam i12729_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12730_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n17412));
    defparam i12730_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12731_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n17413));
    defparam i12731_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12732_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34627), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n17414));
    defparam i12732_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n33975));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n16967));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n34101));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n16965));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0][0] ), .C(clk32MHz), .D(n16964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n16963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n16962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n16961));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1116 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34810));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i12712_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n17394));
    defparam i12712_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n17392));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12713_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n17395));
    defparam i12713_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(150[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12714_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n17396));
    defparam i12714_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n17355));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n17354));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n17405));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n34887));   // verilog/coms.v(228[9:81])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i12715_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n17397));
    defparam i12715_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12716_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n17398));
    defparam i12716_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12709_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34635), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n17391));
    defparam i12709_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1118 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[17] [4]), .I3(GND_net), .O(n6_adj_3952));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1118.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1119 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[10] [6]), .O(n35182));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36422 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n43194));
    defparam byte_transmit_counter_0__bdd_4_lut_36422.LUT_INIT = 16'he4aa;
    SB_LUT4 i12685_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n17367));
    defparam i12685_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12686_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n17368));
    defparam i12686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12687_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n17369));
    defparam i12687_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12688_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n17370));
    defparam i12688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12689_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n17371));
    defparam i12689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12690_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n17372));
    defparam i12690_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12691_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n17373));
    defparam i12691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12692_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34647), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n17374));
    defparam i12692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12761_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n17443));
    defparam i12761_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12764_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n17446));
    defparam i12764_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12763_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n17445));
    defparam i12763_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12762_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n17444));
    defparam i12762_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12757_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n17439));
    defparam i12757_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_1173_i10_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/coms.v(163[9:87])
    defparam equal_1173_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12758_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n17440));
    defparam i12758_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1046_i1_3_lut (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4291), .I3(GND_net), .O(n4292));
    defparam mux_1046_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12759_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n17441));
    defparam i12759_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12760_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34643), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n17442));
    defparam i12760_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n24172), .O(n34643));   // verilog/coms.v(151[7:23])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1120 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n24172), .O(n34647));   // verilog/coms.v(151[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1120.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1121 (.I0(n24172), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n34635));
    defparam i2_2_lut_3_lut_4_lut_adj_1121.LUT_INIT = 16'hf7ff;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1122 (.I0(n24172), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n34627));
    defparam i2_2_lut_3_lut_4_lut_adj_1122.LUT_INIT = 16'hff7f;
    SB_LUT4 n43194_bdd_4_lut (.I0(n43194), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n43197));
    defparam n43194_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1123 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n26928), .I3(GND_net), .O(n4_adj_3988));
    defparam i1_2_lut_3_lut_adj_1123.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1124 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n121));
    defparam i1_2_lut_3_lut_adj_1124.LUT_INIT = 16'h8080;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36417 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n43188));
    defparam byte_transmit_counter_0__bdd_4_lut_36417.LUT_INIT = 16'he4aa;
    SB_LUT4 n43188_bdd_4_lut (.I0(n43188), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n43191));
    defparam n43188_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1125 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n26928), .I3(GND_net), .O(n2030));
    defparam i1_2_lut_3_lut_adj_1125.LUT_INIT = 16'h7070;
    SB_LUT4 i2_3_lut_4_lut_adj_1126 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n15540), .I3(\FRAME_MATCHER.i [4]), .O(n15329));   // verilog/coms.v(151[7:23])
    defparam i2_3_lut_4_lut_adj_1126.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36412 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n43182));
    defparam byte_transmit_counter_0__bdd_4_lut_36412.LUT_INIT = 16'he4aa;
    SB_LUT4 n43182_bdd_4_lut (.I0(n43182), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n43185));
    defparam n43182_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36407 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n43176));
    defparam byte_transmit_counter_0__bdd_4_lut_36407.LUT_INIT = 16'he4aa;
    SB_LUT4 n43176_bdd_4_lut (.I0(n43176), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n43179));
    defparam n43176_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1127 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(GND_net), .O(n10_adj_4106));   // verilog/coms.v(151[7:23])
    defparam i1_2_lut_3_lut_adj_1127.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1128 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(n22591), .I3(GND_net), .O(Kp_23__N_839));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36402 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n43170));
    defparam byte_transmit_counter_0__bdd_4_lut_36402.LUT_INIT = 16'he4aa;
    SB_LUT4 n43170_bdd_4_lut (.I0(n43170), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n43173));
    defparam n43170_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36397 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n43164));
    defparam byte_transmit_counter_0__bdd_4_lut_36397.LUT_INIT = 16'he4aa;
    SB_LUT4 n43164_bdd_4_lut (.I0(n43164), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n43167));
    defparam n43164_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36392 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n43158));
    defparam byte_transmit_counter_0__bdd_4_lut_36392.LUT_INIT = 16'he4aa;
    SB_LUT4 n43158_bdd_4_lut (.I0(n43158), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n43161));
    defparam n43158_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36387 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n43152));
    defparam byte_transmit_counter_0__bdd_4_lut_36387.LUT_INIT = 16'he4aa;
    SB_LUT4 n43152_bdd_4_lut (.I0(n43152), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n43155));
    defparam n43152_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1129 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_adj_1129.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36382 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n43146));
    defparam byte_transmit_counter_0__bdd_4_lut_36382.LUT_INIT = 16'he4aa;
    SB_LUT4 n43146_bdd_4_lut (.I0(n43146), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n43149));
    defparam n43146_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36377 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n43140));
    defparam byte_transmit_counter_0__bdd_4_lut_36377.LUT_INIT = 16'he4aa;
    SB_LUT4 n43140_bdd_4_lut (.I0(n43140), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n43143));
    defparam n43140_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1130 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(n16085), .I3(n35106), .O(n35019));
    defparam i2_3_lut_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i12749_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n17431));
    defparam i12749_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12750_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n17432));
    defparam i12750_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12751_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n17433));
    defparam i12751_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12752_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n17434));
    defparam i12752_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12753_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n17435));
    defparam i12753_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1131 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n34839));
    defparam i1_2_lut_3_lut_adj_1131.LUT_INIT = 16'h9696;
    SB_LUT4 i12754_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n17436));
    defparam i12754_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12755_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n17437));
    defparam i12755_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12756_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34647), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n17438));
    defparam i12756_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1132 (.I0(n24172), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n34639));   // verilog/coms.v(151[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1132.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1133 (.I0(n24172), .I1(\FRAME_MATCHER.i [0]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [1]), .O(n34631));   // verilog/coms.v(151[7:23])
    defparam i2_2_lut_3_lut_4_lut_adj_1133.LUT_INIT = 16'hffdf;
    SB_LUT4 i12741_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n17423));
    defparam i12741_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12742_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n17424));
    defparam i12742_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12743_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n17425));
    defparam i12743_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12744_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n17426));
    defparam i12744_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12745_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n17427));
    defparam i12745_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12746_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n17428));
    defparam i12746_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12747_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n17429));
    defparam i12747_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i12748_3_lut_4_lut (.I0(n24008), .I1(n34651), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n17430));
    defparam i12748_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i19354_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n24008));
    defparam i19354_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 equal_115_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));
    defparam equal_115_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i2036_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_4023));
    defparam i2036_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i19407_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n15329), .I3(\FRAME_MATCHER.i [31]), .O(n2855));
    defparam i19407_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 equal_122_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_3896));   // verilog/coms.v(151[7:23])
    defparam equal_122_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_116_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_3950));   // verilog/coms.v(151[7:23])
    defparam equal_116_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i12652_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n17334));
    defparam i12652_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12645_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n17327));
    defparam i12645_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12646_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n17328));
    defparam i12646_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12647_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n17329));
    defparam i12647_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1046_i6_3_lut (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4291), .I3(GND_net), .O(n4297));
    defparam mux_1046_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12648_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n17330));
    defparam i12648_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n34973));   // verilog/coms.v(228[9:81])
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i12649_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n17331));
    defparam i12649_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12650_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n17332));
    defparam i12650_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12651_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34635), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n17333));
    defparam i12651_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1046_i5_3_lut (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4291), .I3(GND_net), .O(n4296));
    defparam mux_1046_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1046_i4_3_lut (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4291), .I3(GND_net), .O(n4295));
    defparam mux_1046_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1135 (.I0(n35192), .I1(\data_out_frame[14] [0]), 
            .I2(n35019), .I3(n35234), .O(n35166));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1046_i3_3_lut (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4291), .I3(GND_net), .O(n4294));
    defparam mux_1046_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_337_Select_31_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4084));
    defparam select_337_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_30_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4083));
    defparam select_337_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_4_lut_adj_1136 (.I0(n35192), .I1(\data_out_frame[14] [0]), 
            .I2(n35019), .I3(n16423), .O(n30573));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1046_i2_3_lut (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4291), .I3(GND_net), .O(n4293));
    defparam mux_1046_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_337_Select_29_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4081));
    defparam select_337_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_28_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4079));
    defparam select_337_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 mux_1046_i15_3_lut (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4291), .I3(GND_net), .O(n4306));
    defparam mux_1046_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_337_Select_27_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4077));
    defparam select_337_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 mux_1046_i14_3_lut (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4291), .I3(GND_net), .O(n4305));
    defparam mux_1046_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_337_Select_26_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4075));
    defparam select_337_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_25_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4073));
    defparam select_337_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 mux_1046_i13_3_lut (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4291), .I3(GND_net), .O(n4304));
    defparam mux_1046_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1046_i12_3_lut (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4291), .I3(GND_net), .O(n4303));
    defparam mux_1046_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_337_Select_24_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4071));
    defparam select_337_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 mux_1046_i11_3_lut (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4291), .I3(GND_net), .O(n4302));
    defparam mux_1046_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1046_i10_3_lut (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4291), .I3(GND_net), .O(n4301));
    defparam mux_1046_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1137 (.I0(n15939), .I1(n34960), .I2(GND_net), 
            .I3(GND_net), .O(n31273));
    defparam i1_2_lut_adj_1137.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1138 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[14] [1]), 
            .I2(n12_adj_4107), .I3(n8_adj_4108), .O(n31330));
    defparam i1_4_lut_adj_1138.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1139 (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[15] [5]), 
            .I2(\data_in_frame[15] [6]), .I3(GND_net), .O(n34678));
    defparam i2_3_lut_adj_1139.LUT_INIT = 16'h9696;
    SB_LUT4 select_337_Select_23_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4069));
    defparam select_337_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_in_frame[15] [7]), .I1(n31269), 
            .I2(GND_net), .I3(GND_net), .O(n34737));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16283));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\data_in_frame[13] [6]), .I1(n31234), 
            .I2(GND_net), .I3(GND_net), .O(n35229));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1143 (.I0(\data_in_frame[16] [1]), .I1(n35128), 
            .I2(n34901), .I3(n31284), .O(n36194));
    defparam i3_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1144 (.I0(n35137), .I1(n35270), .I2(n36194), 
            .I3(n31269), .O(n10_adj_4109));
    defparam i4_4_lut_adj_1144.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1145 (.I0(n16283), .I1(n34967), .I2(n34737), 
            .I3(n31284), .O(n15990));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1145.LUT_INIT = 16'h9669;
    SB_LUT4 select_337_Select_22_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4067));
    defparam select_337_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_21_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4065));
    defparam select_337_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_20_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4063));
    defparam select_337_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1146 (.I0(\data_in_frame[19] [7]), .I1(n15990), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4110));
    defparam i1_2_lut_adj_1146.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1147 (.I0(n34712), .I1(n30623), .I2(n35022), 
            .I3(n6_adj_4110), .O(n35001));
    defparam i4_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_18__7__I_0_3230_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1353));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_18__7__I_0_3230_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_337_Select_19_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4061));
    defparam select_337_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i2_3_lut_adj_1148 (.I0(n36871), .I1(\data_in_frame[17] [2]), 
            .I2(\data_in_frame[17] [1]), .I3(GND_net), .O(n35246));
    defparam i2_3_lut_adj_1148.LUT_INIT = 16'h6969;
    SB_LUT4 select_337_Select_18_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4059));
    defparam select_337_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1149 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35270));
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h6666;
    SB_LUT4 select_337_Select_17_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4058));
    defparam select_337_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_16_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4057));
    defparam select_337_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i3_4_lut_adj_1150 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[13] [7]), .I3(\data_in_frame[13] [6]), .O(n15671));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 select_337_Select_15_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4056));
    defparam select_337_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_14_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4055));
    defparam select_337_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i6_4_lut_adj_1151 (.I0(n35270), .I1(\data_in_frame[17] [5]), 
            .I2(n35169), .I3(\data_in_frame[17] [6]), .O(n14_adj_4111));
    defparam i6_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1152 (.I0(\data_in_frame[13] [3]), .I1(n14_adj_4111), 
            .I2(n10_adj_4112), .I3(n34979), .O(n35774));
    defparam i7_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(n15671), .I1(n16057), .I2(GND_net), 
            .I3(GND_net), .O(n34901));
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 select_337_Select_13_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4054));
    defparam select_337_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_12_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4053));
    defparam select_337_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1154 (.I0(n36362), .I1(n31332), .I2(GND_net), 
            .I3(GND_net), .O(n35169));
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1155 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(\data_in_frame[18] [2]), .I3(GND_net), .O(n6_adj_4113));
    defparam i2_3_lut_adj_1155.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1156 (.I0(\data_in_frame[18] [5]), .I1(n6_adj_4113), 
            .I2(Kp_23__N_1353), .I3(\data_in_frame[18] [4]), .O(n34712));
    defparam i3_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 select_337_Select_11_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4052));
    defparam select_337_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i11_4_lut_adj_1157 (.I0(n31234), .I1(n15794), .I2(n35188), 
            .I3(\data_in_frame[13] [1]), .O(n26_adj_4114));   // verilog/coms.v(74[16:43])
    defparam i11_4_lut_adj_1157.LUT_INIT = 16'h9669;
    SB_LUT4 select_337_Select_10_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4051));
    defparam select_337_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_9_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4050));
    defparam select_337_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i9_4_lut_adj_1158 (.I0(\data_in_frame[13] [7]), .I1(n34712), 
            .I2(n35169), .I3(\data_in_frame[15] [3]), .O(n24_adj_4115));   // verilog/coms.v(74[16:43])
    defparam i9_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1159 (.I0(n35088), .I1(\data_in_frame[13] [6]), 
            .I2(n34901), .I3(n35774), .O(n25));   // verilog/coms.v(74[16:43])
    defparam i10_4_lut_adj_1159.LUT_INIT = 16'h9669;
    SB_LUT4 i8_3_lut (.I0(n35025), .I1(n34916), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n23_adj_4116));   // verilog/coms.v(74[16:43])
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut_adj_1160 (.I0(n23_adj_4116), .I1(n25), .I2(n24_adj_4115), 
            .I3(n26_adj_4114), .O(n30623));   // verilog/coms.v(74[16:43])
    defparam i14_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35088));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1162 (.I0(\data_in_frame[8] [7]), .I1(n35252), 
            .I2(n35012), .I3(n16218), .O(n34867));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n34979));
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1164 (.I0(n35172), .I1(\data_in_frame[13] [2]), 
            .I2(n16142), .I3(n35176), .O(n20_adj_4117));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 select_337_Select_8_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4049));
    defparam select_337_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i7_4_lut_adj_1165 (.I0(\data_in_frame[19] [5]), .I1(n35240), 
            .I2(n34766), .I3(\data_in_frame[6] [6]), .O(n19_adj_4118));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1166 (.I0(n34979), .I1(\data_in_frame[6] [4]), 
            .I2(n34702), .I3(n16479), .O(n21_adj_4119));   // verilog/coms.v(74[16:43])
    defparam i9_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1167 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n15788), .I3(n35211), .O(n35192));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 select_337_Select_7_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4048));
    defparam select_337_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i11_3_lut_adj_1168 (.I0(n21_adj_4119), .I1(n19_adj_4118), .I2(n20_adj_4117), 
            .I3(GND_net), .O(n34819));   // verilog/coms.v(74[16:43])
    defparam i11_3_lut_adj_1168.LUT_INIT = 16'h9696;
    SB_LUT4 select_337_Select_6_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4047));
    defparam select_337_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i4_4_lut_adj_1169 (.I0(n34848), .I1(n16286), .I2(n35112), 
            .I3(n6_adj_4103), .O(n35220));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 select_337_Select_5_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4046));
    defparam select_337_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_4_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4045));
    defparam select_337_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 select_337_Select_3_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4044));
    defparam select_337_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i2_3_lut_4_lut_adj_1170 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[13] [5]), .I3(n15586), .O(n34997));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1171 (.I0(\data_in_frame[6] [5]), .I1(n35285), 
            .I2(n35273), .I3(Kp_23__N_969), .O(n35025));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1172 (.I0(n35016), .I1(n35025), .I2(\data_in_frame[15] [2]), 
            .I3(n35012), .O(n12_adj_4120));   // verilog/coms.v(73[16:43])
    defparam i5_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1173 (.I0(n15917), .I1(n12_adj_4120), .I2(n35172), 
            .I3(\data_in_frame[11] [0]), .O(n16391));   // verilog/coms.v(73[16:43])
    defparam i6_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 select_337_Select_2_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4043));
    defparam select_337_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_in_frame[17] [3]), .I1(n16391), 
            .I2(GND_net), .I3(GND_net), .O(n35179));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 select_337_Select_1_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4041));
    defparam select_337_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i2_2_lut_adj_1175 (.I0(\data_in_frame[10] [3]), .I1(n35009), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4121));   // verilog/coms.v(83[17:28])
    defparam i2_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1176 (.I0(Kp_23__N_1083), .I1(n34699), .I2(n35179), 
            .I3(n15939), .O(n14_adj_4122));   // verilog/coms.v(83[17:28])
    defparam i6_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1177 (.I0(\data_in_frame[19] [4]), .I1(n14_adj_4122), 
            .I2(n10_adj_4121), .I3(n35243), .O(n35084));   // verilog/coms.v(83[17:28])
    defparam i7_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 select_337_Select_0_i3_2_lut_4_lut (.I0(n18962), .I1(n2030), 
            .I2(n18939), .I3(\FRAME_MATCHER.i [0]), .O(n3_c));
    defparam select_337_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'h3200;
    SB_LUT4 i1_2_lut_3_lut_adj_1178 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15448), 
            .I2(n121), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2389 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1178.LUT_INIT = 16'h1010;
    SB_LUT4 i5_4_lut_adj_1179 (.I0(n15862), .I1(\data_in_frame[17] [4]), 
            .I2(n35220), .I3(n34819), .O(n12_adj_4123));   // verilog/coms.v(71[16:42])
    defparam i5_4_lut_adj_1179.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1180 (.I0(n34867), .I1(n12_adj_4123), .I2(n35088), 
            .I3(n16391), .O(n34800));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34684));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1182 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15448), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n139), .O(n15437));   // verilog/coms.v(126[12] 289[6])
    defparam i2_3_lut_4_lut_adj_1182.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_adj_1183 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[14] [0]), .I3(GND_net), .O(n35128));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35172));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1185 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[8] [5]), 
            .I2(\data_in_frame[8] [6]), .I3(\data_in_frame[11] [0]), .O(n35188));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1186 (.I0(\data_in_frame[13] [2]), .I1(n35188), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[11] [1]), .O(n35252));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4124));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1188 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[11] [1]), 
            .I2(\data_in_frame[10] [7]), .I3(n6_adj_4124), .O(n34702));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(n15794), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35016));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1190 (.I0(n15798), .I1(n35047), .I2(n35016), 
            .I3(n34702), .O(Kp_23__N_1430));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1191 (.I0(n31269), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n31345));
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(n30605), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34967));
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1193 (.I0(n16394), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[8] [3]), .I3(\data_in_frame[12] [5]), .O(n10_adj_4102));
    defparam i4_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1194 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15448), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n18939));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1194.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1195 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[15] [6]), .I3(\data_out_frame[13] [4]), 
            .O(n35072));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1196 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15448), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n26928));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1196.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1197 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(n34523), .I3(GND_net), .O(n6_adj_3989));
    defparam i1_2_lut_3_lut_adj_1197.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1198 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [13]), 
            .I2(n34673), .I3(GND_net), .O(n6_adj_4040));
    defparam i1_2_lut_3_lut_adj_1198.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n34766));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1200 (.I0(n15_adj_3943), .I1(n16142), .I2(\data_in_frame[11] [2]), 
            .I3(n6_adj_4125), .O(n35047));   // verilog/coms.v(77[16:35])
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(n15803), .I1(n16137), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_969));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1202 (.I0(Kp_23__N_969), .I1(\data_in_frame[8] [6]), 
            .I2(n35047), .I3(n6_adj_4126), .O(n16057));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i12789_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n17471));
    defparam i12789_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35160));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(\data_in_frame[6] [6]), .I1(n15803), 
            .I2(GND_net), .I3(GND_net), .O(n35237));
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35075));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i12791_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n17473));
    defparam i12791_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1206 (.I0(n35075), .I1(n35157), .I2(\data_in_frame[11] [4]), 
            .I3(n34806), .O(n12_adj_4127));
    defparam i5_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1207 (.I0(\data_in_frame[7] [2]), .I1(n12_adj_4127), 
            .I2(n35237), .I3(\data_in_frame[9] [2]), .O(n31234));
    defparam i6_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1208 (.I0(n35160), .I1(n16137), .I2(n34806), 
            .I3(\data_in_frame[9] [1]), .O(n14_adj_4128));
    defparam i6_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1209 (.I0(\data_in_frame[1] [2]), .I1(n34973), 
            .I2(n34887), .I3(n34810), .O(Kp_23__N_858));   // verilog/coms.v(71[16:34])
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1210 (.I0(n16232), .I1(n14_adj_4128), .I2(n10_adj_4129), 
            .I3(\data_in_frame[6] [6]), .O(n31251));
    defparam i7_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i12790_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n17472));
    defparam i12790_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(\data_in_frame[13] [3]), .I1(Kp_23__N_1430), 
            .I2(GND_net), .I3(GND_net), .O(n15862));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1212 (.I0(\data_in_frame[13] [5]), .I1(n31251), 
            .I2(n31234), .I3(\data_in_frame[11] [3]), .O(n30605));
    defparam i3_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i12793_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n17475));
    defparam i12793_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1213 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n35078));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_LUT4 i12792_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n17474));
    defparam i12792_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12796_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n17478));
    defparam i12796_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1214 (.I0(\data_in_frame[13] [4]), .I1(n31251), 
            .I2(\data_in_frame[11] [3]), .I3(n16057), .O(n36362));
    defparam i3_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i12795_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n17477));
    defparam i12795_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1215 (.I0(n36362), .I1(n34916), .I2(\data_in_frame[15] [7]), 
            .I3(GND_net), .O(n35137));
    defparam i2_3_lut_adj_1215.LUT_INIT = 16'h6969;
    SB_LUT4 i12794_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34627), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n17476));
    defparam i12794_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12701_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n17383));
    defparam i12701_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35121));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1217 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4130));
    defparam i2_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1218 (.I0(n35163), .I1(\data_in_frame[15] [2]), 
            .I2(n35121), .I3(\data_in_frame[15] [1]), .O(n32_adj_4131));
    defparam i12_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1219 (.I0(\data_in_frame[17] [0]), .I1(n32_adj_4131), 
            .I2(n22_adj_4130), .I3(n35137), .O(n36_adj_4132));
    defparam i16_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1220 (.I0(\data_in_frame[16] [7]), .I1(n35240), 
            .I2(\data_in_frame[14] [7]), .I3(n34967), .O(n34_adj_4133));
    defparam i14_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1221 (.I0(n15794), .I1(\data_in_frame[14] [1]), 
            .I2(\data_in_frame[16] [5]), .I3(\data_in_frame[14] [0]), .O(n35_adj_4134));
    defparam i15_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1222 (.I0(n16277), .I1(n35249), .I2(\data_in_frame[14] [6]), 
            .I3(\data_in_frame[16] [3]), .O(n33));
    defparam i13_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15828));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n34763));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i19_4_lut_adj_1225 (.I0(n33), .I1(n35_adj_4134), .I2(n34_adj_4133), 
            .I3(n36_adj_4132), .O(n36871));
    defparam i19_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1226 (.I0(n15944), .I1(n30555), .I2(\data_in_frame[4] [6]), 
            .I3(\data_in_frame[6] [7]), .O(n28_adj_4135));
    defparam i12_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1227 (.I0(n35223), .I1(n34806), .I2(n34803), 
            .I3(\data_in_frame[6] [5]), .O(n26_adj_4136));
    defparam i10_4_lut_adj_1227.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1228 (.I0(n35226), .I1(n34829), .I2(n35205), 
            .I3(n34731), .O(n27));
    defparam i11_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1229 (.I0(\data_in_frame[6] [1]), .I1(n35054), 
            .I2(\data_in_frame[3] [4]), .I3(n15657), .O(n25_adj_4137));
    defparam i9_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1230 (.I0(n25_adj_4137), .I1(n27), .I2(n26_adj_4136), 
            .I3(n28_adj_4135), .O(n36545));
    defparam i15_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1231 (.I0(n34944), .I1(\data_in_frame[11] [4]), 
            .I2(n34848), .I3(\data_in_frame[10] [2]), .O(n46));
    defparam i19_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1232 (.I0(n34890), .I1(\data_in_frame[11] [3]), 
            .I2(\data_in_frame[9] [6]), .I3(\data_in_frame[12] [2]), .O(n44));
    defparam i17_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1233 (.I0(n35282), .I1(n35160), .I2(n35252), 
            .I3(n35091), .O(n45));
    defparam i18_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1234 (.I0(n36545), .I1(n35273), .I2(n31345), 
            .I3(n35094), .O(n43_adj_4138));
    defparam i16_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1235 (.I0(n35047), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[13] [3]), .I3(n35172), .O(n42_adj_4139));
    defparam i15_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i12702_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n17384));
    defparam i12702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_3_lut_adj_1236 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[15] [0]), 
            .I2(\data_in_frame[16] [4]), .I3(GND_net), .O(n41_adj_4140));
    defparam i14_3_lut_adj_1236.LUT_INIT = 16'h9696;
    SB_LUT4 i12703_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n17385));
    defparam i12703_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i25_4_lut (.I0(n43_adj_4138), .I1(n45), .I2(n44), .I3(n46), 
            .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12704_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n17386));
    defparam i12704_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20_4_lut_adj_1237 (.I0(n15794), .I1(n15671), .I2(n31271), 
            .I3(\data_in_frame[12] [3]), .O(n47_adj_4141));
    defparam i20_4_lut_adj_1237.LUT_INIT = 16'h9669;
    SB_LUT4 i26_4_lut (.I0(n47_adj_4141), .I1(n52), .I2(n41_adj_4140), 
            .I3(n42_adj_4139), .O(n35249));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12705_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n17387));
    defparam i12705_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1238 (.I0(\data_in_frame[15] [4]), .I1(n35249), 
            .I2(n36871), .I3(n34994), .O(n20_adj_4142));
    defparam i8_4_lut_adj_1238.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1239 (.I0(n34898), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[18] [7]), .I3(n35176), .O(n19_adj_4143));
    defparam i7_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1240 (.I0(\data_in_frame[15] [2]), .I1(n15862), 
            .I2(n36362), .I3(\data_in_frame[16] [1]), .O(n21_adj_4144));
    defparam i9_4_lut_adj_1240.LUT_INIT = 16'h9669;
    SB_LUT4 i11_3_lut_adj_1241 (.I0(n21_adj_4144), .I1(n19_adj_4143), .I2(n20_adj_4142), 
            .I3(GND_net), .O(n30609));
    defparam i11_3_lut_adj_1241.LUT_INIT = 16'h9696;
    SB_LUT4 i12706_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n17388));
    defparam i12706_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12707_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n17389));
    defparam i12707_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1242 (.I0(\data_in_frame[19] [7]), .I1(n34800), 
            .I2(n34940), .I3(n35084), .O(n8_adj_4145));
    defparam i3_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1243 (.I0(n30623), .I1(n8_adj_4145), .I2(\data_in_frame[19] [2]), 
            .I3(\data_in_frame[19] [1]), .O(n16183));
    defparam i4_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16394));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n15780));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_in_frame[3] [3]), .I1(Kp_23__N_893), 
            .I2(GND_net), .I3(GND_net), .O(n34803));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1247 (.I0(\data_in_frame[12] [3]), .I1(n35091), 
            .I2(n16289), .I3(n16394), .O(n10_adj_4105));
    defparam i4_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1248 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[11] [2]), .O(n34835));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i12708_3_lut_4_lut (.I0(n10_adj_3950), .I1(n34639), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n17390));
    defparam i12708_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16277));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1250 (.I0(n92[1]), .I1(n63_adj_4002), .I2(n4), 
            .I3(GND_net), .O(n33967));   // verilog/coms.v(141[4] 143[7])
    defparam i1_2_lut_3_lut_adj_1250.LUT_INIT = 16'hb0b0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36372 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n43134));
    defparam byte_transmit_counter_0__bdd_4_lut_36372.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_in_frame[11] [7]), .I1(n35148), 
            .I2(GND_net), .I3(GND_net), .O(n31271));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1252 (.I0(\FRAME_MATCHER.i_31__N_2392 ), .I1(n3741), 
            .I2(n4), .I3(GND_net), .O(n5));
    defparam i1_2_lut_3_lut_adj_1252.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16479));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1254 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[12] [0]), 
            .I2(n31271), .I3(n16277), .O(n34925));
    defparam i3_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1255 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[8] [2]), .I3(GND_net), .O(n35282));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1255.LUT_INIT = 16'h9696;
    SB_LUT4 n43134_bdd_4_lut (.I0(n43134), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n43137));
    defparam n43134_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36367 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n43128));
    defparam byte_transmit_counter_0__bdd_4_lut_36367.LUT_INIT = 16'he4aa;
    SB_LUT4 n43128_bdd_4_lut (.I0(n43128), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n43131));
    defparam n43128_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35094));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.i_31__N_2392 ), .I1(n3741), 
            .I2(n63_adj_4002), .I3(n92[1]), .O(n30072));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h2202;
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(n63_adj_4011), .I1(n22667), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n92[1]));   // verilog/coms.v(93[12:19])
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1258 (.I0(n2030), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_3896), 
            .O(n34654));
    defparam i1_2_lut_3_lut_4_lut_adj_1258.LUT_INIT = 16'hfff7;
    SB_LUT4 i2_3_lut_adj_1259 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[7] [5]), .I3(GND_net), .O(n34825));
    defparam i2_3_lut_adj_1259.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1260 (.I0(Kp_23__N_896), .I1(n34757), .I2(\data_in_frame[4] [7]), 
            .I3(GND_net), .O(n35223));
    defparam i2_3_lut_adj_1260.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1261 (.I0(n30573), .I1(n16457), .I2(n34953), 
            .I3(n34909), .O(n34910));
    defparam i1_2_lut_3_lut_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(n34757), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35157));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n34964));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1264 (.I0(n30555), .I1(n34806), .I2(\data_in_frame[7] [3]), 
            .I3(GND_net), .O(n30553));
    defparam i2_3_lut_adj_1264.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1265 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[7] [3]), .I3(GND_net), .O(n35264));
    defparam i2_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1266 (.I0(n2030), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_3950), 
            .O(n34651));
    defparam i1_2_lut_3_lut_4_lut_adj_1266.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_adj_1267 (.I0(n63_adj_4011), .I1(n22667), .I2(n63_adj_4002), 
            .I3(GND_net), .O(n10283));   // verilog/coms.v(93[12:19])
    defparam i1_2_lut_3_lut_adj_1267.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4147));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1269 (.I0(n30553), .I1(n15_adj_3943), .I2(n34890), 
            .I3(n6_adj_4147), .O(n35148));
    defparam i4_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1270 (.I0(n35223), .I1(n34825), .I2(n15871), 
            .I3(n35264), .O(n10_adj_4148));
    defparam i4_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n34693));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1272 (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[14] [1]), 
            .I2(\data_in_frame[14] [2]), .I3(n31261), .O(n34994));
    defparam i1_4_lut_adj_1272.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1273 (.I0(\FRAME_MATCHER.state [2]), .I1(n26928), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2386 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1273.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_1274 (.I0(\FRAME_MATCHER.state [2]), .I1(n26928), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2392 ));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1274.LUT_INIT = 16'h4040;
    SB_LUT4 i3_4_lut_adj_1275 (.I0(n16232), .I1(n35148), .I2(n34944), 
            .I3(n15944), .O(n31284));
    defparam i3_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(n34964), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[11] [5]), .I3(n35157), .O(n10_adj_4149));
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1277 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n34013));
    defparam i1_2_lut_3_lut_adj_1277.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_adj_1278 (.I0(n16142), .I1(n10_adj_4149), .I2(n30553), 
            .I3(GND_net), .O(n31269));
    defparam i5_3_lut_adj_1278.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1279 (.I0(n31269), .I1(n31284), .I2(n34994), 
            .I3(\data_in_frame[13] [7]), .O(n37099));
    defparam i3_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1280 (.I0(\data_in_frame[19] [0]), .I1(n34925), 
            .I2(n35163), .I3(n6_adj_4150), .O(n16400));
    defparam i4_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1281 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n34015));
    defparam i1_2_lut_3_lut_adj_1281.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1282 (.I0(n31261), .I1(n30585), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4151));
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1283 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[14] [4]), 
            .I2(\data_in_frame[14] [3]), .I3(n6_adj_4151), .O(n31332));
    defparam i4_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1284 (.I0(\data_in_frame[9] [6]), .I1(n30555), 
            .I2(\data_in_frame[7] [4]), .I3(\data_in_frame[7] [5]), .O(n34960));
    defparam i3_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_858), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[0] [5]), .O(n35069));   // verilog/coms.v(68[16:69])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1285 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n34017));
    defparam i1_2_lut_3_lut_adj_1285.LUT_INIT = 16'he0e0;
    SB_LUT4 data_in_frame_7__7__I_0_2_lut (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1083));   // verilog/coms.v(83[17:28])
    defparam data_in_frame_7__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\data_in_frame[6] [4]), .I1(n16137), 
            .I2(GND_net), .I3(GND_net), .O(n35185));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut_adj_1287 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n16400), .I3(n16183), .O(n6_adj_3920));
    defparam i2_2_lut_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1288 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[20] [4]), .I3(\data_in_frame[18] [2]), .O(n14_adj_4152));
    defparam i5_3_lut_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(n15756), .I1(n15794), .I2(GND_net), 
            .I3(GND_net), .O(n15657));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n34019));
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1291 (.I0(n15756), .I1(n15794), .I2(\data_in_frame[10] [6]), 
            .I3(\data_in_frame[6] [2]), .O(n35012));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1292 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n34021));
    defparam i1_2_lut_3_lut_adj_1292.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(\data_in_frame[14] [6]), .I1(n35285), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4153));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1294 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[17] [2]), 
            .I2(\data_in_frame[10] [5]), .I3(n6_adj_4153), .O(n34699));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1295 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n34023));
    defparam i1_2_lut_3_lut_adj_1295.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1296 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n34025));
    defparam i1_2_lut_3_lut_adj_1296.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1297 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[12] [2]), 
            .I2(\data_in_frame[10] [1]), .I3(n6_adj_4154), .O(n34928));
    defparam i4_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1298 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[14] [4]), .I3(GND_net), .O(n35267));
    defparam i2_3_lut_adj_1298.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35112));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1300 (.I0(\data_in_frame[8] [4]), .I1(n15798), 
            .I2(\data_in_frame[14] [7]), .I3(\data_in_frame[15] [0]), .O(n35009));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n34721));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1302 (.I0(n34721), .I1(\data_in_frame[17] [0]), 
            .I2(n35226), .I3(n35009), .O(n16_adj_4155));
    defparam i6_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1303 (.I0(\data_in_frame[12] [6]), .I1(n35112), 
            .I2(n35267), .I3(n34928), .O(n17_adj_4156));
    defparam i7_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1304 (.I0(n17_adj_4156), .I1(\data_in_frame[14] [6]), 
            .I2(n16_adj_4155), .I3(\data_in_frame[17] [1]), .O(n31258));
    defparam i9_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1305 (.I0(n34699), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[17] [1]), .I3(n35012), .O(n20_adj_4157));   // verilog/coms.v(72[16:43])
    defparam i8_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1306 (.I0(\data_in_frame[19] [3]), .I1(n35185), 
            .I2(\data_in_frame[8] [5]), .I3(\data_in_frame[6] [1]), .O(n19_adj_4158));   // verilog/coms.v(72[16:43])
    defparam i7_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1307 (.I0(n34684), .I1(n30585), .I2(\data_in_frame[14] [5]), 
            .I3(\data_in_frame[13] [0]), .O(n21_adj_4159));   // verilog/coms.v(72[16:43])
    defparam i9_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1308 (.I0(n21_adj_4159), .I1(n19_adj_4158), .I2(n20_adj_4157), 
            .I3(GND_net), .O(n34940));   // verilog/coms.v(72[16:43])
    defparam i11_3_lut_adj_1308.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1309 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n34027));
    defparam i1_2_lut_3_lut_adj_1309.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1310 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n34029));
    defparam i1_2_lut_3_lut_adj_1310.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1311 (.I0(\data_in_frame[21] [4]), .I1(n34940), 
            .I2(n31258), .I3(\data_in_frame[19] [2]), .O(n36828));
    defparam i3_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1312 (.I0(n16183), .I1(\data_in_frame[20] [7]), 
            .I2(n31258), .I3(n30609), .O(n8_adj_4160));
    defparam i1_4_lut_adj_1312.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1313 (.I0(n31332), .I1(\data_in_frame[18] [7]), 
            .I2(n16400), .I3(n37099), .O(n12_adj_4161));
    defparam i5_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1314 (.I0(\data_in_frame[18] [1]), .I1(n35022), 
            .I2(\data_in_frame[18] [2]), .I3(\data_in_frame[20] [3]), .O(n36991));
    defparam i2_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1315 (.I0(n35179), .I1(n35220), .I2(\data_in_frame[20] [0]), 
            .I3(n35001), .O(n12_adj_4162));
    defparam i5_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1316 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[21] [3]), 
            .I2(\data_in_frame[19] [1]), .I3(GND_net), .O(n4_adj_4163));
    defparam i1_3_lut_adj_1316.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1317 (.I0(n34678), .I1(n12_adj_4162), .I2(n35246), 
            .I3(n34916), .O(n36693));
    defparam i6_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i1_rep_142_3_lut (.I0(n16183), .I1(n31258), .I2(n30609), .I3(GND_net), 
            .O(n43740));
    defparam i1_rep_142_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1318 (.I0(n35229), .I1(n34678), .I2(n34867), 
            .I3(\data_in_frame[20] [2]), .O(n14_adj_4164));
    defparam i6_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1319 (.I0(\data_in_frame[18] [1]), .I1(n35121), 
            .I2(n34737), .I3(\data_in_frame[17] [6]), .O(n13_adj_4165));
    defparam i5_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1320 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n34031));
    defparam i1_2_lut_3_lut_adj_1320.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1321 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n34033));
    defparam i1_2_lut_3_lut_adj_1321.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_4_lut_adj_1322 (.I0(n34925), .I1(n31330), .I2(n34928), 
            .I3(n31273), .O(n12_adj_4166));
    defparam i5_4_lut_adj_1322.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n34035));
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_4_lut_adj_1324 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[12] [1]), 
            .I2(n10_adj_4148), .I3(\data_in_frame[11] [7]), .O(n31261));
    defparam i5_3_lut_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1325 (.I0(n34757), .I1(\data_in_frame[7] [4]), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[7] [3]), .O(n34944));
    defparam i1_2_lut_4_lut_adj_1325.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1326 (.I0(n35774), .I1(n35001), .I2(\data_in_frame[20] [1]), 
            .I3(n31332), .O(n36974));
    defparam i3_4_lut_adj_1326.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1327 (.I0(n13_adj_4165), .I1(\data_in_frame[21] [1]), 
            .I2(n14_adj_4164), .I3(n43740), .O(n20_adj_4167));
    defparam i4_4_lut_adj_1327.LUT_INIT = 16'hde7b;
    SB_LUT4 i4_4_lut_adj_1328 (.I0(\data_in_frame[18] [5]), .I1(n16286), 
            .I2(\data_in_frame[18] [4]), .I3(\data_in_frame[20] [6]), .O(n11));
    defparam i4_4_lut_adj_1328.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1329 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n34037));
    defparam i1_2_lut_3_lut_adj_1329.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1330 (.I0(\data_in_frame[4] [7]), .I1(Kp_23__N_896), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n34890));
    defparam i1_2_lut_3_lut_adj_1330.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1331 (.I0(n34901), .I1(\data_in_frame[18] [3]), 
            .I2(n31330), .I3(n34898), .O(n15_adj_4168));
    defparam i6_4_lut_adj_1331.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_1332 (.I0(n37099), .I1(n15990), .I2(\data_in_frame[20] [5]), 
            .I3(GND_net), .O(n8_adj_4169));
    defparam i3_3_lut_adj_1332.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1333 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(n34845), .I3(n4_adj_3995), .O(n34864));
    defparam i1_2_lut_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1334 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(n35267), .I3(GND_net), .O(n35163));
    defparam i1_2_lut_3_lut_adj_1334.LUT_INIT = 16'h9696;
    SB_LUT4 i8_4_lut_adj_1335 (.I0(n15_adj_4168), .I1(n30605), .I2(n14_adj_4152), 
            .I3(n31269), .O(n36119));
    defparam i8_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1336 (.I0(\data_in_frame[19] [1]), .I1(n34935), 
            .I2(n30609), .I3(\data_in_frame[21] [2]), .O(n36799));
    defparam i3_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36362 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n43122));
    defparam byte_transmit_counter_0__bdd_4_lut_36362.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1337 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n34039));
    defparam i1_2_lut_3_lut_adj_1337.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n34041));
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'he0e0;
    SB_LUT4 i31351_4_lut (.I0(n34819), .I1(n36828), .I2(n35084), .I3(\data_in_frame[21] [6]), 
            .O(n38053));
    defparam i31351_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n34043));
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'he0e0;
    SB_LUT4 n43122_bdd_4_lut (.I0(n43122), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n43125));
    defparam n43122_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1340 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[9] [7]), .I3(\data_in_frame[7] [5]), .O(n35091));
    defparam i1_2_lut_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1341 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n3_adj_3897));   // verilog/coms.v(163[9:87])
    defparam i1_2_lut_3_lut_adj_1341.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1342 (.I0(\data_in_frame[18] [5]), .I1(n36991), 
            .I2(n12_adj_4161), .I3(n8_adj_4160), .O(n22_adj_3907));
    defparam i6_4_lut_adj_1342.LUT_INIT = 16'hedde;
    SB_LUT4 i7_4_lut_adj_1343 (.I0(n36119), .I1(\data_in_frame[18] [3]), 
            .I2(n8_adj_4169), .I3(\data_in_frame[18] [4]), .O(n23));
    defparam i7_4_lut_adj_1343.LUT_INIT = 16'hd77d;
    SB_LUT4 i5_4_lut_adj_1344 (.I0(n36799), .I1(\data_in_frame[21] [5]), 
            .I2(n34940), .I3(n35084), .O(n21));
    defparam i5_4_lut_adj_1344.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_3_lut_adj_1345 (.I0(\data_in_frame[21] [0]), .I1(n31258), 
            .I2(n30609), .I3(GND_net), .O(n5_c));
    defparam i1_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1346 (.I0(n43), .I1(n34668), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n33977));
    defparam i1_2_lut_3_lut_adj_1346.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_4_lut_adj_1347 (.I0(n31258), .I1(n36693), .I2(n4_adj_4163), 
            .I3(n30609), .O(n18));
    defparam i2_4_lut_adj_1347.LUT_INIT = 16'hdeed;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n7_adj_4100));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36357 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n43116));
    defparam byte_transmit_counter_0__bdd_4_lut_36357.LUT_INIT = 16'he4aa;
    SB_LUT4 n43116_bdd_4_lut (.I0(n43116), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n43119));
    defparam n43116_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1349 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n34149));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1349.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1350 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n34147));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1350.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n7_adj_4098));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n34145));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n34143));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'he0e0;
    SB_LUT4 i10_4_lut_adj_1354 (.I0(n11), .I1(n20_adj_4167), .I2(n36974), 
            .I3(n12_adj_4166), .O(n26_adj_3924));
    defparam i10_4_lut_adj_1354.LUT_INIT = 16'hfefd;
    SB_LUT4 i1_2_lut_3_lut_adj_1355 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n34141));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1355.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n34139));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n34137));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1358 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n34135));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1358.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1359 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n34133));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1359.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36352 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n43110));
    defparam byte_transmit_counter_0__bdd_4_lut_36352.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n7_adj_4095));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_4_lut_adj_1361 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(n30613), .I3(n10_adj_3901), .O(n35131));
    defparam i5_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i19302_2_lut_3_lut (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n23956));   // verilog/coms.v(113[11:12])
    defparam i19302_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n7_adj_4093));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(n30605), .I1(\data_in_frame[13] [3]), 
            .I2(Kp_23__N_1430), .I3(GND_net), .O(n34916));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n34131));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_3_lut_adj_1365 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(\data_in_frame[6] [5]), .I3(GND_net), .O(n10_adj_4129));
    defparam i2_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n7_adj_4090));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1367 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[9] [0]), 
            .I2(n35205), .I3(GND_net), .O(n6_adj_4126));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1367.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [0]), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n6_adj_4125));   // verilog/coms.v(77[16:35])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n34129));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(n15798), .I1(\data_in_frame[6] [4]), 
            .I2(n16137), .I3(n16218), .O(n35205));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(n15798), .I1(\data_in_frame[6] [4]), 
            .I2(n16137), .I3(GND_net), .O(n15917));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1372 (.I0(n16142), .I1(\data_in_frame[6] [6]), 
            .I2(n15803), .I3(GND_net), .O(n16218));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1372.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n35273));
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1374 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[16] [0]), 
            .I2(\data_in_frame[15] [6]), .I3(\data_in_frame[14] [0]), .O(n34898));
    defparam i1_2_lut_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1375 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[15] [1]), .I3(GND_net), .O(n35176));
    defparam i1_2_lut_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 n43110_bdd_4_lut (.I0(n43110), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n43113));
    defparam n43110_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1376 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n34127));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1376.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_4_lut_adj_1377 (.I0(n36871), .I1(\data_in_frame[17] [2]), 
            .I2(\data_in_frame[17] [1]), .I3(Kp_23__N_1430), .O(n10_adj_4112));
    defparam i2_2_lut_4_lut_adj_1377.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n34125));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n34123));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut_adj_1380 (.I0(n13), .I1(n11_adj_4170), .I2(n15828), 
            .I3(n22591), .O(n35109));   // verilog/coms.v(69[16:69])
    defparam i7_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1381 (.I0(\data_in_frame[13] [6]), .I1(n31234), 
            .I2(n10_adj_4109), .I3(\data_in_frame[16] [0]), .O(n35022));
    defparam i5_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n34121));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36347 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n43104));
    defparam byte_transmit_counter_0__bdd_4_lut_36347.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n34119));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'he0e0;
    SB_LUT4 i22_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_844));   // verilog/coms.v(94[12:25])
    defparam i22_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n7_adj_4087));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1385 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n34117));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1385.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n34115));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n7_adj_4085));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n34113));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1389 (.I0(n17_adj_4016), .I1(n42), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n34111));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1389.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1390 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [31]), .O(n8_adj_4101));
    defparam i1_2_lut_4_lut_adj_1390.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1391 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [28]), .O(n8_adj_4099));
    defparam i1_2_lut_4_lut_adj_1391.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1392 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(n15693), .I3(GND_net), .O(n35198));
    defparam i1_2_lut_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(\data_out_frame[13] [2]), .I1(n1504), 
            .I2(n35060), .I3(GND_net), .O(n34795));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1394 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [24]), .O(n8_adj_4097));
    defparam i1_2_lut_4_lut_adj_1394.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1395 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [20]), .O(n8_adj_4096));
    defparam i1_2_lut_4_lut_adj_1395.LUT_INIT = 16'hfe00;
    SB_LUT4 n43104_bdd_4_lut (.I0(n43104), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n43107));
    defparam n43104_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1396 (.I0(\data_out_frame[13] [2]), .I1(n1504), 
            .I2(n34785), .I3(n30571), .O(n35063));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i19953_2_lut_4_lut (.I0(n31_adj_4010), .I1(n41_adj_4015), .I2(n43), 
            .I3(\FRAME_MATCHER.state [19]), .O(n24611));
    defparam i19953_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i5_3_lut_4_lut_adj_1397 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[13] [6]), 
            .I2(n31234), .I3(n31273), .O(n12_adj_4107));
    defparam i5_3_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1398 (.I0(\data_in_frame[11] [7]), .I1(n35148), 
            .I2(n31269), .I3(\data_in_frame[12] [0]), .O(n8_adj_4108));
    defparam i1_2_lut_4_lut_adj_1398.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n16400), .I3(GND_net), .O(n34935));
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1400 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [18]), .O(n8_adj_4094));
    defparam i1_2_lut_4_lut_adj_1400.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1401 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [17]), .O(n8_adj_4092));
    defparam i1_2_lut_4_lut_adj_1401.LUT_INIT = 16'hfe00;
    SB_LUT4 i19517_2_lut_3_lut (.I0(n2030), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n24172));
    defparam i19517_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(n3_adj_3897), .O(n11_adj_4170));   // verilog/coms.v(163[9:87])
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1402 (.I0(n34789), .I1(n15154), .I2(n1507), 
            .I3(n30559), .O(n6_adj_3914));   // verilog/coms.v(73[16:43])
    defparam i2_2_lut_3_lut_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1403 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(n34960), .I3(\data_in_frame[8] [0]), .O(n6_adj_4154));
    defparam i1_2_lut_3_lut_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1404 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [16]), .O(n8_adj_4091));
    defparam i1_2_lut_4_lut_adj_1404.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1405 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [11]), .O(n8_adj_4089));
    defparam i1_2_lut_4_lut_adj_1405.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1406 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [9]), .O(n8_adj_4088));
    defparam i1_2_lut_4_lut_adj_1406.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1407 (.I0(n31_adj_4010), .I1(n41_adj_4015), 
            .I2(n43), .I3(\FRAME_MATCHER.state [6]), .O(n8_adj_4086));
    defparam i1_2_lut_4_lut_adj_1407.LUT_INIT = 16'hfe00;
    SB_LUT4 i12773_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n17455));
    defparam i12773_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1408 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(n34960), .I3(n35243), .O(n6_adj_4150));
    defparam i1_2_lut_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_4_lut (.I0(n24524), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n12905), .O(n30171));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h7775;
    SB_LUT4 i12780_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n17462));
    defparam i12780_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1409 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[5] [6]), .I3(n15780), .O(n16286));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1410 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n24524));
    defparam i2_2_lut_3_lut_adj_1410.LUT_INIT = 16'hfefe;
    SB_LUT4 i12779_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n17461));
    defparam i12779_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12778_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n17460));
    defparam i12778_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12777_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n17459));
    defparam i12777_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12776_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n17458));
    defparam i12776_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12775_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n17457));
    defparam i12775_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12774_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34635), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n17456));
    defparam i12774_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12672_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n17354));
    defparam i12672_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12673_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n17355));
    defparam i12673_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12674_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n17356));
    defparam i12674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12675_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n17357));
    defparam i12675_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12676_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n17358));
    defparam i12676_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12670_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n17352));
    defparam i12670_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1411 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(n35131), .I3(\data_out_frame[20] [7]), .O(n36199));
    defparam i2_3_lut_4_lut_adj_1411.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1412 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(n34921), .I3(GND_net), .O(n9_adj_4032));
    defparam i1_2_lut_3_lut_adj_1412.LUT_INIT = 16'h9696;
    SB_LUT4 i12671_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n17353));
    defparam i12671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(n34744), .I1(\data_out_frame[15] [0]), 
            .I2(\data_out_frame[14] [7]), .I3(GND_net), .O(n35255));
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1414 (.I0(n30523), .I1(\data_out_frame[17] [3]), 
            .I2(n34744), .I3(n35034), .O(n6_adj_4027));
    defparam i1_2_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1415 (.I0(n35063), .I1(\data_out_frame[20] [1]), 
            .I2(n30619), .I3(n34988), .O(n34990));
    defparam i1_2_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i12669_3_lut_4_lut (.I0(n8), .I1(n34654), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n17351));
    defparam i12669_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_365_Select_1_i1_3_lut_4_lut (.I0(n92[1]), .I1(\FRAME_MATCHER.i_31__N_2386 ), 
            .I2(n63_adj_4002), .I3(n737), .O(n1));
    defparam select_365_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i12661_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n17343));
    defparam i12661_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1416 (.I0(\FRAME_MATCHER.state [2]), .I1(n22667), 
            .I2(n63_adj_4011), .I3(n63_adj_4002), .O(\FRAME_MATCHER.state_31__N_2426[2] ));   // verilog/coms.v(141[7:84])
    defparam i1_2_lut_4_lut_adj_1416.LUT_INIT = 16'hb300;
    SB_LUT4 i12662_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n17344));
    defparam i12662_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12663_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n17345));
    defparam i12663_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35585_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(GND_net), .O(n42349));
    defparam i35585_2_lut_3_lut.LUT_INIT = 16'h1e1e;
    SB_LUT4 i1_3_lut_4_lut_adj_1417 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[1]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[3]), 
            .O(n84));   // verilog/coms.v(100[12:33])
    defparam i1_3_lut_4_lut_adj_1417.LUT_INIT = 16'haa80;
    SB_LUT4 i1_3_lut_4_lut_adj_1418 (.I0(\FRAME_MATCHER.state[3] ), .I1(n10283), 
            .I2(n2720), .I3(n42), .O(n33969));
    defparam i1_3_lut_4_lut_adj_1418.LUT_INIT = 16'haa80;
    SB_LUT4 i12664_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n17346));
    defparam i12664_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12665_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n17347));
    defparam i12665_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12666_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n17348));
    defparam i12666_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12667_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n17349));
    defparam i12667_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12668_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34627), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n17350));
    defparam i12668_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12765_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n17447));
    defparam i12765_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12772_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n17454));
    defparam i12772_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12771_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n17453));
    defparam i12771_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12770_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n17452));
    defparam i12770_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12769_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n17451));
    defparam i12769_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1419 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n6));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1419.LUT_INIT = 16'h9696;
    SB_LUT4 i12768_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n17450));
    defparam i12768_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1420 (.I0(n16160), .I1(n35069), .I2(n10_adj_3994), 
            .I3(\data_in_frame[0] [7]), .O(n34792));   // verilog/coms.v(68[16:27])
    defparam i5_3_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i36293_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n16737));
    defparam i36293_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i12767_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n17449));
    defparam i12767_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(\FRAME_MATCHER.state [2]), .I1(n24524), 
            .I2(n34530), .I3(GND_net), .O(n4_adj_3993));   // verilog/coms.v(110[11:16])
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'h5454;
    SB_LUT4 i12766_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34639), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n17448));
    defparam i12766_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1422 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [6]), .I3(n15828), .O(n15756));   // verilog/coms.v(228[9:81])
    defparam i2_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1423 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[2] [3]), 
            .I2(n34693), .I3(n3_adj_3897), .O(n15803));   // verilog/coms.v(72[16:43])
    defparam i2_2_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1424 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state_31__N_2490 [3]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n36175));
    defparam i2_3_lut_4_lut_adj_1424.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_2_lut_4_lut_adj_1425 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n35380), .O(n16593));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_4_lut_adj_1425.LUT_INIT = 16'h0002;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [3]), 
            .I2(n15923), .I3(n35201), .O(n17_adj_3957));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1426 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[9] [0]), .I3(GND_net), .O(n16110));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1426.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1427 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[8] [2]), .O(n34816));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1428 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[10] [4]), .I3(GND_net), .O(n35081));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_1428.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1429 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[15] [5]), .I3(GND_net), .O(n34789));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1430 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(n35100), .I3(\data_out_frame[11] [1]), .O(n1507));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1431 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[11] [2]), .I3(GND_net), .O(n34855));
    defparam i1_2_lut_3_lut_adj_1431.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1432 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n13978));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1432.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1433 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[10] [7]), .I3(n34835), .O(n35100));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1434 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n34772));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1434.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[10] [7]), .I3(GND_net), .O(n15831));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1436 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[9] [2]), .I3(n13862), .O(n35118));
    defparam i2_3_lut_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1437 (.I0(n34884), .I1(\data_out_frame[20] [3]), 
            .I2(n15923), .I3(n34931), .O(n35146));
    defparam i1_2_lut_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1438 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(n35276), .I3(GND_net), .O(n35258));
    defparam i1_2_lut_3_lut_adj_1438.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1439 (.I0(\data_out_frame[14] [5]), .I1(n30611), 
            .I2(n15693), .I3(GND_net), .O(n31275));
    defparam i1_2_lut_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_LUT4 i12783_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n17465));
    defparam i12783_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12782_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n17464));
    defparam i12782_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12781_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n17463));
    defparam i12781_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1440 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n23_adj_3936));
    defparam i2_2_lut_3_lut_adj_1440.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1441 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[12] [3]), 
            .I2(n10_adj_3931), .I3(\data_out_frame[12] [2]), .O(n30591));   // verilog/coms.v(83[17:28])
    defparam i5_3_lut_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i12785_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n17467));
    defparam i12785_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12784_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n17466));
    defparam i12784_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12787_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n17469));
    defparam i12787_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12786_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n17468));
    defparam i12786_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12788_3_lut_4_lut (.I0(n10_adj_4106), .I1(n34631), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n17470));
    defparam i12788_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1442 (.I0(Kp_23__N_844), .I1(n34693), .I2(\data_in_frame[0] [3]), 
            .I3(GND_net), .O(n22591));   // verilog/coms.v(94[12:25])
    defparam i2_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1443 (.I0(n30573), .I1(n16457), .I2(n34953), 
            .I3(GND_net), .O(n31279));
    defparam i1_2_lut_3_lut_adj_1443.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1444 (.I0(n15154), .I1(\data_out_frame[17] [1]), 
            .I2(n34921), .I3(GND_net), .O(n35141));
    defparam i1_2_lut_3_lut_adj_1444.LUT_INIT = 16'h9696;
    SB_LUT4 i22355_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n12859));   // verilog/coms.v(110[11:16])
    defparam i22355_4_lut_4_lut.LUT_INIT = 16'h0102;
    SB_LUT4 i12653_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n17335));
    defparam i12653_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12654_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n17336));
    defparam i12654_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1445 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n35004));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1445.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1446 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[7] [3]), .O(n34718));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1447 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[5] [5]), .O(n34778));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1448 (.I0(\data_out_frame[20] [2]), .I1(n30571), 
            .I2(n34884), .I3(n34877), .O(n35126));
    defparam i1_2_lut_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i12655_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n17337));
    defparam i12655_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12656_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n17338));
    defparam i12656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1449 (.I0(\data_out_frame[12] [5]), .I1(n34813), 
            .I2(\data_out_frame[12] [6]), .I3(\data_out_frame[6] [3]), .O(n34744));
    defparam i1_2_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i12657_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n17339));
    defparam i12657_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12658_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n17340));
    defparam i12658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(\data_out_frame[12] [0]), .I1(n35208), 
            .I2(n15788), .I3(n35031), .O(n6_adj_3917));
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1451 (.I0(\data_out_frame[20] [2]), .I1(n30571), 
            .I2(n34884), .I3(n34870), .O(n35232));
    defparam i1_2_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i12659_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n17341));
    defparam i12659_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12660_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34631), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n17342));
    defparam i12660_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12637_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n17319));
    defparam i12637_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12638_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n17320));
    defparam i12638_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1452 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[11] [7]), .I3(GND_net), .O(n35031));
    defparam i1_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1453 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(n35097), .I3(GND_net), .O(n6_adj_3916));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1453.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1454 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[16] [2]), .I3(GND_net), .O(n35276));
    defparam i1_2_lut_3_lut_adj_1454.LUT_INIT = 16'h9696;
    SB_LUT4 i12639_3_lut_4_lut (.I0(n10_adj_3896), .I1(n34639), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n17321));
    defparam i12639_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1455 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[9] [3]), .I3(\data_out_frame[9] [1]), .O(n35103));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1456 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [5]), 
            .I2(n35201), .I3(GND_net), .O(n35279));
    defparam i1_2_lut_3_lut_adj_1456.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut (.I0(\data_out_frame[14] [7]), .I1(n12), .I2(n8_adj_4171), 
            .I3(GND_net), .O(n34991));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut_adj_1457 (.I0(\data_out_frame[13] [2]), .I1(n34997), 
            .I2(\data_out_frame[13] [1]), .I3(n31226), .O(n8_adj_4171));
    defparam i1_2_lut_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1458 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[17] [5]), .I3(n1593), .O(n34785));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1459 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[11] [0]), .O(n6_adj_3903));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    uart_tx tx (.n318(n318), .r_Clock_Count({Open_7, Open_8, Open_9, 
            Open_10, Open_11, \r_Clock_Count[3] , Open_12, \r_Clock_Count[1] , 
            Open_13}), .GND_net(GND_net), .n16918(n16918), .r_Bit_Index({r_Bit_Index}), 
            .clk32MHz(clk32MHz), .n16915(n16915), .n16911(n16911), .n16890(n16890), 
            .\r_Clock_Count[8] (\r_Clock_Count[8] ), .n16893(n16893), .\r_Clock_Count[7] (\r_Clock_Count[7] ), 
            .n16905(n16905), .n16899(n16899), .\r_Clock_Count[5] (\r_Clock_Count[5] ), 
            .n17029(n17029), .n17566(n17566), .r_SM_Main({r_SM_Main}), 
            .n26602(n26602), .n320(n320), .VCC_net(VCC_net), .tx_data({tx_data}), 
            .n4613(n4613), .n26612(n26612), .n16641(n16641), .n16772(n16772), 
            .tx_o(tx_o), .tx_enable(tx_enable), .n313(n313), .n314(n314), 
            .n16981(n16981), .n16979(n16979), .n316(n316), .n3(n3), 
            .\r_SM_Main_2__N_3323[0] (r_SM_Main_2__N_3323[0]), .n29(n29), 
            .\byte_transmit_counter[7] (byte_transmit_counter[7]), .n37977(n37977), 
            .n15437(n15437), .n63(n63), .n24117(n24117), .tx_transmit_N_3220(tx_transmit_N_3220), 
            .n1205(n1205)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n16872(n16872), .\r_Clock_Count[6] (\r_Clock_Count[6] ), 
            .n16869(n16869), .\r_Clock_Count[7] (\r_Clock_Count[7]_adj_3 ), 
            .n16881(n16881), .\r_Clock_Count[3] (\r_Clock_Count[3]_adj_4 ), 
            .n16887(n16887), .\r_Clock_Count[1] (\r_Clock_Count[1]_adj_5 ), 
            .n17005(n17005), .r_Bit_Index({r_Bit_Index_adj_13}), .n17002(n17002), 
            .n17550(n17550), .rx_data({rx_data}), .r_Rx_Data(r_Rx_Data), 
            .PIN_13_N_105(PIN_13_N_105), .n219(n219), .GND_net(GND_net), 
            .n220(n220), .n30(n30), .n223(n223), .n3(n3_adj_9), .n225(n225), 
            .VCC_net(VCC_net), .rx_data_ready(rx_data_ready), .n15459(n15459), 
            .n4(n4_adj_10), .n16746(n16746), .n16635(n16635), .n17012(n17012), 
            .n17011(n17011), .n17010(n17010), .n17009(n17009), .n17008(n17008), 
            .n17007(n17007), .n17006(n17006), .n4591(n4591), .n24014(n24014), 
            .n4_adj_1(n4_adj_11), .n4_adj_2(n4_adj_12), .n15454(n15454)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n318, r_Clock_Count, GND_net, n16918, r_Bit_Index, 
            clk32MHz, n16915, n16911, n16890, \r_Clock_Count[8] , 
            n16893, \r_Clock_Count[7] , n16905, n16899, \r_Clock_Count[5] , 
            n17029, n17566, r_SM_Main, n26602, n320, VCC_net, tx_data, 
            n4613, n26612, n16641, n16772, tx_o, tx_enable, n313, 
            n314, n16981, n16979, n316, n3, \r_SM_Main_2__N_3323[0] , 
            n29, \byte_transmit_counter[7] , n37977, n15437, n63, 
            n24117, tx_transmit_N_3220, n1205) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output n318;
    output [8:0]r_Clock_Count;
    input GND_net;
    input n16918;
    output [2:0]r_Bit_Index;
    input clk32MHz;
    input n16915;
    input n16911;
    input n16890;
    output \r_Clock_Count[8] ;
    input n16893;
    output \r_Clock_Count[7] ;
    input n16905;
    input n16899;
    output \r_Clock_Count[5] ;
    input n17029;
    input n17566;
    output [2:0]r_SM_Main;
    output n26602;
    output n320;
    input VCC_net;
    input [7:0]tx_data;
    output n4613;
    output n26612;
    output n16641;
    output n16772;
    output tx_o;
    output tx_enable;
    output n313;
    output n314;
    input n16981;
    input n16979;
    output n316;
    output n3;
    input \r_SM_Main_2__N_3323[0] ;
    output n29;
    input \byte_transmit_counter[7] ;
    output n37977;
    input n15437;
    input n63;
    output n24117;
    input tx_transmit_N_3220;
    output n1205;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n27968, n27969, n16908;
    wire [8:0]r_Clock_Count_c;   // verilog/uart_tx.v(32[16:29])
    
    wire n16896, n26643, n17604, n40066, n27967, n27966, n40063, 
        n13073;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n152, n38074, n24585, n10, n219, n18734, n27973, n27972, 
        n16980, tx_active, n36075, n40065, n27971, n27970, n40064, 
        n38173, n38174, n38243, n38242, o_Tx_Serial_N_3351, n8784, 
        n16577, n43098;
    
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n27968), .O(n318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n27968), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n27969));
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n16918));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n16915));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n16911));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count_c[2]), .C(clk32MHz), .D(n16908));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(\r_Clock_Count[8] ), .C(clk32MHz), .D(n16890));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count_c[6]), .C(clk32MHz), .D(n16896));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(\r_Clock_Count[7] ), .C(clk32MHz), .D(n16893));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n16905));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count_c[4]), .C(clk32MHz), .D(n26643));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(\r_Clock_Count[5] ), .C(clk32MHz), .D(n16899));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17029));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count_c[0]), .C(clk32MHz), .D(n17604));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n17566));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_4_lut (.I0(n26602), .I1(r_Clock_Count_c[2]), .I2(GND_net), 
            .I3(n27967), .O(n40066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_4 (.CI(n27967), .I0(r_Clock_Count_c[2]), .I1(GND_net), 
            .CO(n27968));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n27966), .O(n320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n27966), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n27967));
    SB_LUT4 add_59_2_lut (.I0(n26602), .I1(r_Clock_Count_c[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n40063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count_c[0]), .I1(GND_net), 
            .CO(n27966));
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i22081_3_lut (.I0(r_Clock_Count_c[2]), .I1(n40066), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16908));
    defparam i22081_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n152));   // verilog/uart_tx.v(31[16:25])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i195_4_lut (.I0(n152), .I1(r_SM_Main[2]), .I2(n38074), .I3(\r_Clock_Count[7] ), 
            .O(n26602));   // verilog/uart_tx.v(31[16:25])
    defparam i195_4_lut.LUT_INIT = 16'hccce;
    SB_LUT4 i1290_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4613));   // verilog/uart_tx.v(98[36:51])
    defparam i1290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n24585));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count_c[0]), .I1(\r_Clock_Count[5] ), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[1]), .O(n10));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count_c[2]), .I1(n10), .I2(r_Clock_Count_c[4]), 
            .I3(GND_net), .O(n219));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n26612), .O(n16641));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i12090_3_lut (.I0(n16641), .I1(r_SM_Main[1]), .I2(n24585), 
            .I3(GND_net), .O(n16772));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12090_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_2_lut_adj_872 (.I0(r_SM_Main[0]), .I1(n26612), .I2(GND_net), 
            .I3(GND_net), .O(n18734));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_872.LUT_INIT = 16'h8888;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n13073), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22036_3_lut (.I0(r_Clock_Count_c[0]), .I1(n40063), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n17604));
    defparam i22036_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(\r_Clock_Count[8] ), .I2(GND_net), 
            .I3(n27973), .O(n313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(\r_Clock_Count[7] ), .I2(GND_net), 
            .I3(n27972), .O(n314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n16981));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n16980));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n16979));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n36075));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_9 (.CI(n27972), .I0(\r_Clock_Count[7] ), .I1(GND_net), 
            .CO(n27973));
    SB_LUT4 add_59_8_lut (.I0(n26602), .I1(r_Clock_Count_c[6]), .I2(GND_net), 
            .I3(n27971), .O(n40065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_8 (.CI(n27971), .I0(r_Clock_Count_c[6]), .I1(GND_net), 
            .CO(n27972));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(\r_Clock_Count[5] ), .I2(GND_net), 
            .I3(n27970), .O(n316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n27970), .I0(\r_Clock_Count[5] ), .I1(GND_net), 
            .CO(n27971));
    SB_LUT4 add_59_6_lut (.I0(n26602), .I1(r_Clock_Count_c[4]), .I2(GND_net), 
            .I3(n27969), .O(n40064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_6 (.CI(n27969), .I0(r_Clock_Count_c[4]), .I1(GND_net), 
            .CO(n27970));
    SB_LUT4 i31411_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n38173));
    defparam i31411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31412_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n38174));
    defparam i31412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31481_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n38243));
    defparam i31481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31480_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n38242));
    defparam i31480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22099_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3351), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_tx.v(31[16:25])
    defparam i22099_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i1_2_lut_adj_873 (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n8784));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_873.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut_adj_874 (.I0(n8784), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n18734), .O(n16577));
    defparam i2_4_lut_adj_874.LUT_INIT = 16'h3202;
    SB_LUT4 i14531_3_lut (.I0(n16577), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n16980));   // verilog/uart_tx.v(31[16:25])
    defparam i14531_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i22051_3_lut (.I0(r_Clock_Count_c[4]), .I1(n40064), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n26643));
    defparam i22051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24_4_lut (.I0(\r_SM_Main_2__N_3323[0] ), .I1(n24585), .I2(r_SM_Main[1]), 
            .I3(n26612), .O(n29));   // verilog/uart_tx.v(31[16:25])
    defparam i24_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i22066_3_lut (.I0(r_Clock_Count_c[6]), .I1(n40065), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n16896));
    defparam i22066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(n26612), .O(n36075));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i3_3_lut_4_lut (.I0(\r_SM_Main_2__N_3323[0] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n13073));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i31275_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(\byte_transmit_counter[7] ), .I3(GND_net), .O(n37977));
    defparam i31275_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i19462_3_lut_4_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(n15437), .I3(n63), .O(n24117));
    defparam i19462_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(tx_transmit_N_3220), .I3(GND_net), .O(n1205));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i31371_2_lut_3_lut (.I0(r_Clock_Count_c[6]), .I1(\r_Clock_Count[8] ), 
            .I2(n219), .I3(GND_net), .O(n38074));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i31371_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_3_lut_4_lut_adj_875 (.I0(r_Clock_Count_c[6]), .I1(\r_Clock_Count[8] ), 
            .I2(\r_Clock_Count[7] ), .I3(n219), .O(n26612));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_3_lut_4_lut_adj_875.LUT_INIT = 16'hfffe;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n38242), 
            .I2(n38243), .I3(r_Bit_Index[2]), .O(n43098));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n43098_bdd_4_lut (.I0(n43098), .I1(n38174), .I2(n38173), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3351));
    defparam n43098_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n16872, \r_Clock_Count[6] , n16869, \r_Clock_Count[7] , 
            n16881, \r_Clock_Count[3] , n16887, \r_Clock_Count[1] , 
            n17005, r_Bit_Index, n17002, n17550, rx_data, r_Rx_Data, 
            PIN_13_N_105, n219, GND_net, n220, n30, n223, n3, 
            n225, VCC_net, rx_data_ready, n15459, n4, n16746, n16635, 
            n17012, n17011, n17010, n17009, n17008, n17007, n17006, 
            n4591, n24014, n4_adj_1, n4_adj_2, n15454) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n16872;
    output \r_Clock_Count[6] ;
    input n16869;
    output \r_Clock_Count[7] ;
    input n16881;
    output \r_Clock_Count[3] ;
    input n16887;
    output \r_Clock_Count[1] ;
    input n17005;
    output [2:0]r_Bit_Index;
    input n17002;
    input n17550;
    output [7:0]rx_data;
    output r_Rx_Data;
    input PIN_13_N_105;
    output n219;
    input GND_net;
    output n220;
    output n30;
    output n223;
    output n3;
    output n225;
    input VCC_net;
    output rx_data_ready;
    output n15459;
    output n4;
    output n16746;
    output n16635;
    input n17012;
    input n17011;
    input n17010;
    input n17009;
    input n17008;
    input n17007;
    input n17006;
    output n4591;
    output n24014;
    output n4_adj_1;
    output n4_adj_2;
    output n15454;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n17605;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n16878, n17645, n16884, n17552;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n17549, r_Rx_Data_R, n27965, n27964;
    wire [31:0]n194;
    
    wire n27963, n40088, n27962, n27961, n55, n6, n80, n6_adj_3893, 
        n40084, n40067, n27960;
    wire [2:0]r_SM_Main_2__N_3249;
    
    wire n34611, n27959, n34191, n15320, n36763, n61, n18845, 
        n40160, n34620, n40225, n43248, n43251, n16972, n34534, 
        n16563, n23, n36924, n36923, n40226;
    
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n17605));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(\r_Clock_Count[6] ), .C(clk32MHz), .D(n16872));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(\r_Clock_Count[7] ), .C(clk32MHz), .D(n16869));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n16878));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n17645));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n16884));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(\r_Clock_Count[3] ), .C(clk32MHz), .D(n16881));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(\r_Clock_Count[1] ), .C(clk32MHz), .D(n16887));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17005));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17002));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n17552));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17549));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n17550));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_105));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 add_62_9_lut (.I0(GND_net), .I1(\r_Clock_Count[7] ), .I2(GND_net), 
            .I3(n27965), .O(n219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(\r_Clock_Count[6] ), .I2(GND_net), 
            .I3(n27964), .O(n220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_8 (.CI(n27964), .I0(\r_Clock_Count[6] ), .I1(GND_net), 
            .CO(n27965));
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n27963), .O(n194[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n27963), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n27964));
    SB_LUT4 add_62_6_lut (.I0(n30), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n27962), .O(n40088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n27962), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n27963));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(\r_Clock_Count[3] ), .I2(GND_net), 
            .I3(n27961), .O(n223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n27961), .I0(\r_Clock_Count[3] ), .I1(GND_net), 
            .CO(n27962));
    SB_LUT4 i1_2_lut (.I0(\r_Clock_Count[6] ), .I1(\r_Clock_Count[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n55));   // verilog/uart_rx.v(32[17:30])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_860 (.I0(\r_Clock_Count[3] ), .I1(\r_Clock_Count[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/uart_rx.v(32[17:30])
    defparam i1_2_lut_adj_860.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(n6), .O(n80));   // verilog/uart_rx.v(32[17:30])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(n6_adj_3893), 
            .I3(n55), .O(n3));
    defparam i1_4_lut.LUT_INIT = 16'haaea;
    SB_LUT4 i21702_3_lut (.I0(r_Clock_Count[0]), .I1(n40084), .I2(n3), 
            .I3(GND_net), .O(n17605));
    defparam i21702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_62_4_lut (.I0(n30), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n27960), .O(n40067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3249[2]), 
            .R(n34611));   // verilog/uart_rx.v(49[10] 144[8])
    SB_CARRY add_62_4 (.CI(n27960), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n27961));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(\r_Clock_Count[1] ), .I2(GND_net), 
            .I3(n27959), .O(n225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n27959), .I0(\r_Clock_Count[1] ), .I1(GND_net), 
            .CO(n27960));
    SB_LUT4 add_62_2_lut (.I0(n30), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n40084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n27959));
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n34191));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3249[2]), .O(n15320));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_adj_861 (.I0(r_Bit_Index[0]), .I1(n15320), .I2(GND_net), 
            .I3(GND_net), .O(n15459));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_861.LUT_INIT = 16'heeee;
    SB_LUT4 equal_137_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_137_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n36763));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14359_4_lut (.I0(n16746), .I1(n36763), .I2(n16635), .I3(r_Bit_Index[0]), 
            .O(n17549));
    defparam i14359_4_lut.LUT_INIT = 16'h05c0;
    SB_LUT4 i1_2_lut_adj_862 (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3249[2]), 
            .I2(GND_net), .I3(GND_net), .O(n61));
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h8888;
    SB_LUT4 i33795_3_lut (.I0(n18845), .I1(r_Rx_Data), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n40160));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i33795_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i1_4_lut_adj_863 (.I0(r_SM_Main[2]), .I1(n40160), .I2(n61), 
            .I3(r_SM_Main[1]), .O(n17552));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut_adj_863.LUT_INIT = 16'h0544;
    SB_LUT4 i1_2_lut_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(n18845), 
            .I3(GND_net), .O(n34620));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(n80), 
            .I3(r_Clock_Count[5]), .O(n6_adj_3893));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 n43248_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(n40225), 
            .I3(n43248), .O(n43251));   // verilog/uart_rx.v(41[10] 45[8])
    defparam n43248_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n17012));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n17011));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n17010));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n17009));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n17008));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n17007));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n17006));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n16972));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1268_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4591));   // verilog/uart_rx.v(102[36:51])
    defparam i1268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_864 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(GND_net), .O(n34534));
    defparam i2_3_lut_adj_864.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3249[2]), .O(n16635));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3249[2]), 
            .I3(r_SM_Main[0]), .O(n16563));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n16563), 
            .I3(rx_data_ready), .O(n34191));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i36282_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n34611));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i36282_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i12081_3_lut (.I0(n16635), .I1(r_SM_Main[1]), .I2(n34534), 
            .I3(GND_net), .O(n16746));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12081_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_2_lut_adj_865 (.I0(r_SM_Main[2]), .I1(n43251), .I2(GND_net), 
            .I3(GND_net), .O(n16972));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_865.LUT_INIT = 16'h4444;
    SB_LUT4 i21699_3_lut (.I0(r_Clock_Count[2]), .I1(n40067), .I2(n3), 
            .I3(GND_net), .O(n16884));
    defparam i21699_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_866 (.I0(n30), .I1(r_Clock_Count[5]), .I2(n194[5]), 
            .I3(n3), .O(n17645));
    defparam i1_4_lut_adj_866.LUT_INIT = 16'h88a0;
    SB_LUT4 i21705_3_lut (.I0(r_Clock_Count[4]), .I1(n40088), .I2(n3), 
            .I3(GND_net), .O(n16878));
    defparam i21705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_867 (.I0(r_SM_Main[1]), .I1(\r_Clock_Count[6] ), 
            .I2(r_Clock_Count[5]), .I3(\r_Clock_Count[7] ), .O(n23));
    defparam i1_4_lut_adj_867.LUT_INIT = 16'h5554;
    SB_LUT4 i2_4_lut_adj_868 (.I0(r_Clock_Count[5]), .I1(n55), .I2(n80), 
            .I3(r_SM_Main[1]), .O(n36924));
    defparam i2_4_lut_adj_868.LUT_INIT = 16'h1300;
    SB_LUT4 i2_4_lut_adj_869 (.I0(n80), .I1(n23), .I2(n55), .I3(n34620), 
            .O(n36923));
    defparam i2_4_lut_adj_869.LUT_INIT = 16'hffcd;
    SB_LUT4 i2_4_lut_adj_870 (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(n36923), 
            .I3(n36924), .O(n30));
    defparam i2_4_lut_adj_870.LUT_INIT = 16'hffec;
    SB_LUT4 i19360_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n24014));
    defparam i19360_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_132_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_132_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_134_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_134_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_871 (.I0(n15320), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n15454));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_871.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Clock_Count[5]), .I1(\r_Clock_Count[6] ), 
            .I2(\r_Clock_Count[7] ), .I3(n80), .O(r_SM_Main_2__N_3249[2]));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_Clock_Count[5]), .I1(n80), .I2(\r_Clock_Count[6] ), 
            .I3(\r_Clock_Count[7] ), .O(n18845));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i34075_2_lut_3_lut_4_lut (.I0(r_Clock_Count[5]), .I1(n80), .I2(\r_Clock_Count[6] ), 
            .I3(\r_Clock_Count[7] ), .O(n40225));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i34075_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i34126_2_lut_4_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(r_SM_Main_2__N_3249[2]), .O(n40226));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34126_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(r_SM_Main_2__N_3249[2]), .I1(r_SM_Main[1]), 
            .I2(n40226), .I3(r_SM_Main[0]), .O(n43248));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n17519, encoder0_position, clk32MHz, 
            n17520, n17521, n17522, n17523, n17524, n17515, n17516, 
            n17517, n17518, n17513, n17514, n17511, n17512, n17509, 
            n17510, n17507, n17508, n17505, n17506, n17502, n17503, 
            n17504, data_o, n2940, GND_net, count_enable, n16968, 
            n17551, reg_B, n37155, PIN_2_c_0, PIN_1_c_1, n16971) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n17519;
    output [23:0]encoder0_position;
    input clk32MHz;
    input n17520;
    input n17521;
    input n17522;
    input n17523;
    input n17524;
    input n17515;
    input n17516;
    input n17517;
    input n17518;
    input n17513;
    input n17514;
    input n17511;
    input n17512;
    input n17509;
    input n17510;
    input n17507;
    input n17508;
    input n17505;
    input n17506;
    input n17502;
    input n17503;
    input n17504;
    output [1:0]data_o;
    output [23:0]n2940;
    input GND_net;
    output count_enable;
    input n16968;
    input n17551;
    output [1:0]reg_B;
    output n37155;
    input PIN_2_c_0;
    input PIN_1_c_1;
    input n16971;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, n2936, n28046, n28045, n28044, n28043, 
        n28042, n28041, n28040, count_direction, n28039, n28038, 
        n28037, n28036, n28035, n28034, n28033, n28032, n28031, 
        n28030, n28029, n28028, n28027, n28026, n28025, n28024, 
        n28023;
    
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n17519));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n17520));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n17521));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n17522));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n17523));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n17524));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n17515));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n17516));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n17517));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n17518));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n17513));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n17514));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n17511));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n17512));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n17509));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n17510));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n17507));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n17508));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n17505));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n17506));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n17502));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n17503));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n17504));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_628_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2936), 
            .I3(n28046), .O(n2940[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2936), 
            .I3(n28045), .O(n2940[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_24 (.CI(n28045), .I0(encoder0_position[22]), .I1(n2936), 
            .CO(n28046));
    SB_LUT4 add_628_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2936), 
            .I3(n28044), .O(n2940[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_23 (.CI(n28044), .I0(encoder0_position[21]), .I1(n2936), 
            .CO(n28045));
    SB_LUT4 add_628_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2936), 
            .I3(n28043), .O(n2940[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_22 (.CI(n28043), .I0(encoder0_position[20]), .I1(n2936), 
            .CO(n28044));
    SB_LUT4 add_628_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2936), 
            .I3(n28042), .O(n2940[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_21 (.CI(n28042), .I0(encoder0_position[19]), .I1(n2936), 
            .CO(n28043));
    SB_LUT4 add_628_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2936), 
            .I3(n28041), .O(n2940[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_20 (.CI(n28041), .I0(encoder0_position[18]), .I1(n2936), 
            .CO(n28042));
    SB_LUT4 add_628_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2936), 
            .I3(n28040), .O(n2940[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_19 (.CI(n28040), .I0(encoder0_position[17]), .I1(n2936), 
            .CO(n28041));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_628_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2936), 
            .I3(n28039), .O(n2940[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_628_18 (.CI(n28039), .I0(encoder0_position[16]), .I1(n2936), 
            .CO(n28040));
    SB_LUT4 add_628_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2936), 
            .I3(n28038), .O(n2940[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_17 (.CI(n28038), .I0(encoder0_position[15]), .I1(n2936), 
            .CO(n28039));
    SB_LUT4 add_628_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2936), 
            .I3(n28037), .O(n2940[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_16 (.CI(n28037), .I0(encoder0_position[14]), .I1(n2936), 
            .CO(n28038));
    SB_LUT4 add_628_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2936), 
            .I3(n28036), .O(n2940[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_15 (.CI(n28036), .I0(encoder0_position[13]), .I1(n2936), 
            .CO(n28037));
    SB_LUT4 add_628_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2936), 
            .I3(n28035), .O(n2940[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_14 (.CI(n28035), .I0(encoder0_position[12]), .I1(n2936), 
            .CO(n28036));
    SB_LUT4 add_628_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2936), 
            .I3(n28034), .O(n2940[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_13 (.CI(n28034), .I0(encoder0_position[11]), .I1(n2936), 
            .CO(n28035));
    SB_LUT4 add_628_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2936), 
            .I3(n28033), .O(n2940[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_12 (.CI(n28033), .I0(encoder0_position[10]), .I1(n2936), 
            .CO(n28034));
    SB_LUT4 add_628_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2936), 
            .I3(n28032), .O(n2940[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_11 (.CI(n28032), .I0(encoder0_position[9]), .I1(n2936), 
            .CO(n28033));
    SB_LUT4 add_628_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2936), 
            .I3(n28031), .O(n2940[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_10 (.CI(n28031), .I0(encoder0_position[8]), .I1(n2936), 
            .CO(n28032));
    SB_LUT4 add_628_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2936), 
            .I3(n28030), .O(n2940[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_9 (.CI(n28030), .I0(encoder0_position[7]), .I1(n2936), 
            .CO(n28031));
    SB_LUT4 add_628_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2936), 
            .I3(n28029), .O(n2940[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_8 (.CI(n28029), .I0(encoder0_position[6]), .I1(n2936), 
            .CO(n28030));
    SB_LUT4 add_628_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2936), 
            .I3(n28028), .O(n2940[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_7 (.CI(n28028), .I0(encoder0_position[5]), .I1(n2936), 
            .CO(n28029));
    SB_LUT4 add_628_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2936), 
            .I3(n28027), .O(n2940[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_6 (.CI(n28027), .I0(encoder0_position[4]), .I1(n2936), 
            .CO(n28028));
    SB_LUT4 add_628_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2936), 
            .I3(n28026), .O(n2940[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_5 (.CI(n28026), .I0(encoder0_position[3]), .I1(n2936), 
            .CO(n28027));
    SB_LUT4 add_628_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2936), 
            .I3(n28025), .O(n2940[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_4 (.CI(n28025), .I0(encoder0_position[2]), .I1(n2936), 
            .CO(n28026));
    SB_LUT4 add_628_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2936), 
            .I3(n28024), .O(n2940[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_3 (.CI(n28024), .I0(encoder0_position[1]), .I1(n2936), 
            .CO(n28025));
    SB_LUT4 add_628_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n28023), .O(n2940[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_2 (.CI(n28023), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n28024));
    SB_CARRY add_628_1 (.CI(GND_net), .I0(n2936), .I1(n2936), .CO(n28023));
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n16968));   // quad.v(35[10] 41[6])
    SB_LUT4 i900_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2936));   // quad.v(37[5] 40[8])
    defparam i900_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n17551(n17551), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .n37155(n37155), .GND_net(GND_net), 
            .PIN_2_c_0(PIN_2_c_0), .PIN_1_c_1(PIN_1_c_1), .n16971(n16971)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n17551, data_o, clk32MHz, reg_B, n37155, 
            GND_net, PIN_2_c_0, PIN_1_c_1, n16971) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n17551;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    output n37155;
    input GND_net;
    input PIN_2_c_0;
    input PIN_1_c_1;
    input n16971;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3559, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n17551));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1180__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[2]), 
            .I3(GND_net), .O(n37155));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_2_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n37155), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22929_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22929_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR cnt_reg_1180__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1180__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_1_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n16971));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i22938_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22938_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22931_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22931_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n2890, encoder1_position, GND_net, 
            n17542, clk32MHz, n17543, n17544, n17545, n17546, n17547, 
            n17548, n17534, n17535, n17536, n17537, n17538, n17539, 
            n17540, n17541, n17530, n17531, n17532, n17533, n17526, 
            n17527, n17528, n17529, data_o, count_enable, n16970, 
            n17597, PIN_6_c_0, reg_B, PIN_7_c_1, n36606, n16990) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n2890;
    output [23:0]encoder1_position;
    input GND_net;
    input n17542;
    input clk32MHz;
    input n17543;
    input n17544;
    input n17545;
    input n17546;
    input n17547;
    input n17548;
    input n17534;
    input n17535;
    input n17536;
    input n17537;
    input n17538;
    input n17539;
    input n17540;
    input n17541;
    input n17530;
    input n17531;
    input n17532;
    input n17533;
    input n17526;
    input n17527;
    input n17528;
    input n17529;
    output [1:0]data_o;
    output count_enable;
    input n16970;
    input n17597;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    output n36606;
    input n16990;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n2880, n28070, n28069, n28068, n28067, n28066, n28065, 
        n28064, B_delayed, A_delayed, n28063, n28062, n28061, n28060, 
        n28059, n28058, n28057, n28056, n28055, n28054, n28053, 
        n28052, n28051, n28050, n28049, n28048, count_direction, 
        n28047;
    
    SB_LUT4 add_602_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2880), 
            .I3(n28070), .O(n2890[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_602_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2880), 
            .I3(n28069), .O(n2890[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_24 (.CI(n28069), .I0(encoder1_position[22]), .I1(n2880), 
            .CO(n28070));
    SB_LUT4 add_602_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2880), 
            .I3(n28068), .O(n2890[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_23 (.CI(n28068), .I0(encoder1_position[21]), .I1(n2880), 
            .CO(n28069));
    SB_LUT4 add_602_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2880), 
            .I3(n28067), .O(n2890[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_22 (.CI(n28067), .I0(encoder1_position[20]), .I1(n2880), 
            .CO(n28068));
    SB_LUT4 add_602_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2880), 
            .I3(n28066), .O(n2890[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n17542));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n17543));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n17544));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n17545));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n17546));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n17547));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n17548));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n17534));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n17535));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n17536));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n17537));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n17538));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n17539));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n17540));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n17541));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n17530));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n17531));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n17532));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n17533));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n17526));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n17527));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n17528));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n17529));   // quad.v(35[10] 41[6])
    SB_CARRY add_602_21 (.CI(n28066), .I0(encoder1_position[19]), .I1(n2880), 
            .CO(n28067));
    SB_LUT4 add_602_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2880), 
            .I3(n28065), .O(n2890[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_20 (.CI(n28065), .I0(encoder1_position[18]), .I1(n2880), 
            .CO(n28066));
    SB_LUT4 add_602_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2880), 
            .I3(n28064), .O(n2890[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_602_19 (.CI(n28064), .I0(encoder1_position[17]), .I1(n2880), 
            .CO(n28065));
    SB_LUT4 add_602_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2880), 
            .I3(n28063), .O(n2890[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_18 (.CI(n28063), .I0(encoder1_position[16]), .I1(n2880), 
            .CO(n28064));
    SB_LUT4 add_602_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2880), 
            .I3(n28062), .O(n2890[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_17 (.CI(n28062), .I0(encoder1_position[15]), .I1(n2880), 
            .CO(n28063));
    SB_LUT4 add_602_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2880), 
            .I3(n28061), .O(n2890[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_16 (.CI(n28061), .I0(encoder1_position[14]), .I1(n2880), 
            .CO(n28062));
    SB_LUT4 add_602_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2880), 
            .I3(n28060), .O(n2890[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_15 (.CI(n28060), .I0(encoder1_position[13]), .I1(n2880), 
            .CO(n28061));
    SB_LUT4 add_602_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2880), 
            .I3(n28059), .O(n2890[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_14 (.CI(n28059), .I0(encoder1_position[12]), .I1(n2880), 
            .CO(n28060));
    SB_LUT4 add_602_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2880), 
            .I3(n28058), .O(n2890[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_13 (.CI(n28058), .I0(encoder1_position[11]), .I1(n2880), 
            .CO(n28059));
    SB_LUT4 add_602_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2880), 
            .I3(n28057), .O(n2890[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_12 (.CI(n28057), .I0(encoder1_position[10]), .I1(n2880), 
            .CO(n28058));
    SB_LUT4 add_602_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2880), 
            .I3(n28056), .O(n2890[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_11 (.CI(n28056), .I0(encoder1_position[9]), .I1(n2880), 
            .CO(n28057));
    SB_LUT4 add_602_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2880), 
            .I3(n28055), .O(n2890[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_10 (.CI(n28055), .I0(encoder1_position[8]), .I1(n2880), 
            .CO(n28056));
    SB_LUT4 add_602_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2880), 
            .I3(n28054), .O(n2890[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_9 (.CI(n28054), .I0(encoder1_position[7]), .I1(n2880), 
            .CO(n28055));
    SB_LUT4 add_602_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2880), 
            .I3(n28053), .O(n2890[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_8 (.CI(n28053), .I0(encoder1_position[6]), .I1(n2880), 
            .CO(n28054));
    SB_LUT4 add_602_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2880), 
            .I3(n28052), .O(n2890[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_7 (.CI(n28052), .I0(encoder1_position[5]), .I1(n2880), 
            .CO(n28053));
    SB_LUT4 add_602_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2880), 
            .I3(n28051), .O(n2890[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_6 (.CI(n28051), .I0(encoder1_position[4]), .I1(n2880), 
            .CO(n28052));
    SB_LUT4 add_602_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2880), 
            .I3(n28050), .O(n2890[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_5 (.CI(n28050), .I0(encoder1_position[3]), .I1(n2880), 
            .CO(n28051));
    SB_LUT4 add_602_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2880), 
            .I3(n28049), .O(n2890[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_4 (.CI(n28049), .I0(encoder1_position[2]), .I1(n2880), 
            .CO(n28050));
    SB_LUT4 add_602_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2880), 
            .I3(n28048), .O(n2890[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_3 (.CI(n28048), .I0(encoder1_position[1]), .I1(n2880), 
            .CO(n28049));
    SB_LUT4 add_602_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n28047), .O(n2890[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_602_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_602_2 (.CI(n28047), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n28048));
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_602_1 (.CI(GND_net), .I0(n2880), .I1(n2880), .CO(n28047));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n16970));   // quad.v(35[10] 41[6])
    SB_LUT4 i913_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2880));   // quad.v(37[5] 40[8])
    defparam i913_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n17597(n17597), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B}), .PIN_7_c_1(PIN_7_c_1), 
            .GND_net(GND_net), .n36606(n36606), .n16990(n16990)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n17597, data_o, clk32MHz, PIN_6_c_0, reg_B, 
            PIN_7_c_1, GND_net, n36606, n16990) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n17597;
    output [1:0]data_o;
    input clk32MHz;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    input GND_net;
    output n36606;
    input n16990;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3559, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n17597));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_6_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_7_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1181__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n36606), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22951_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22951_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n36606));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFFSR cnt_reg_1181__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1181__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n16990));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i22960_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22960_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22953_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22953_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (VCC_net, GND_net, \Ki[4] , \Kp[3] , \Kp[6] , 
            \Kp[0] , setpoint, \Kp[4] , \Kp[2] , \Kp[1] , \Kp[5] , 
            \Ki[1] , \Ki[0] , \Ki[5] , \Ki[2] , \Ki[3] , PWMLimit, 
            \Ki[6] , IntegralLimit, \Ki[7] , duty, clk32MHz, \Kp[7] , 
            motor_state, n25, n43079) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input VCC_net;
    input GND_net;
    input \Ki[4] ;
    input \Kp[3] ;
    input \Kp[6] ;
    input \Kp[0] ;
    input [23:0]setpoint;
    input \Kp[4] ;
    input \Kp[2] ;
    input \Kp[1] ;
    input \Kp[5] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[5] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input [23:0]PWMLimit;
    input \Ki[6] ;
    input [23:0]IntegralLimit;
    input \Ki[7] ;
    output [23:0]duty;
    input clk32MHz;
    input \Kp[7] ;
    input [23:0]motor_state;
    input n25;
    output n43079;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [23:0]n1;
    
    wire n28156, n29504;
    wire [18:0]n7785;
    
    wire n29505;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3454 ;
    wire [23:0]n1_adj_3891;
    
    wire n28155, n45, n28154;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(31[23:31])
    wire [19:0]n7763;
    
    wire n521, n29503, n448, n29502, n29719;
    wire [21:0]n8013;
    
    wire n29720, n375, n29501;
    wire [47:0]n155;
    
    wire n29718, n302, n29500, n43, n28153, n29717;
    wire [9:0]n8235;
    wire [8:0]n8247;
    
    wire n186, n29886, n229, n29499, n29716, n29887, n156, n29498, 
        n29715, n14, n83, n28015;
    wire [23:0]n2996;
    wire [23:0]n3021;
    
    wire n28016, n41, n28152, n44, n113;
    wire [20:0]n7740;
    
    wire n29497, n29714, n29496;
    wire [23:0]duty_23__N_3478;
    
    wire n28014, n39, n28151, n29713, n29495, n37, n28150, n35, 
        n28149;
    wire [10:0]n8222;
    
    wire n29885, n29494, n29712, n33, n28148, n29884, n29493, 
        n29711, n305, n28013, n29883, n29710, n29882, n29709, 
        n29492, n548, n29881, n4_adj_3565;
    wire [2:0]n8001;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    wire [3:0]n7995;
    
    wire n490, n12;
    wire [23:0]n1_adj_3892;
    
    wire n6_adj_3566, n8_adj_3567, n11, n6_adj_3568, n27680, n475, 
        n29880, n29708, n18, n29491, n13, n29490, n4_adj_3569, 
        n36676, n31, n28147, n29707, n29489, n29488, n29706, n402, 
        n29879, n29705, n329, n29878, n512, n29704, n256, n29877, 
        n77, n8_adj_3570, n378, n439, n29703, n150, n223, n256_adj_3571, 
        n296, n27621, n369, n442, n183_adj_3572, n29876, n41_adj_3573, 
        n110, n366, n29702, n515;
    wire [11:0]n8208;
    
    wire n29875, n29874, n29873, n293, n29701, n107, n29872, n220, 
        n29700, n29487, n147, n29699, n29486, n28012, n38, n29485, 
        n29, n28146;
    wire [23:0]duty_23__N_3355;
    wire [23:0]\PID_CONTROLLER.err_23__N_3379 ;
    
    wire n5_adj_3575, n74, n29871;
    wire [20:0]n8037;
    
    wire n29698, n545, n29870, n29697, n29484, n27, n28145, n472, 
        n29869, n29696, n29695, n518, n29483, n28011, n180, n25_adj_3577, 
        n28144, n445, n29482, n29694, n399, n29868, n372, n29481, 
        n29693, n24213, n253, n326, n299, n29480, n28010, n80, 
        n29692, n11_adj_3579, n29691, n29690, n29689, n153, n29688, 
        n23, n28143, n226, n29479, n29687, n29478, n29867, n29686, 
        n29866, n29685;
    wire [0:0]n6169;
    wire [21:0]n7716;
    
    wire n29477, n29476, n29684, n29865, n21_adj_3581, n28142, n28009;
    wire [23:0]n28;
    
    wire n28742;
    wire [12:0]n8193;
    
    wire n29864, n28741, n29863, n29683, n29475, n28740, n28008, 
        n28739, n29862, n29474, n29473, n29472, n28738, n29471, 
        n29861, n19, n28141, n28737, n98, n29_adj_3584, n451, 
        n29682, n29470, n171, n524, n29681, n244, n29860, n29680, 
        n29469, n28007, n28736, n29468, n28735, n29679, n29467, 
        n29678, n28734, n29859, n29466;
    wire [5:0]n7980;
    
    wire n29677, n29465, n317;
    wire [4:0]n7988;
    
    wire n417, n29676, n542, n29858, n469, n29857, n29464, n344, 
        n29675, n271, n29674, n396, n29856, n28733, n29463, n28732, 
        n198_adj_3589, n29673, n29462, n323, n29855, n250, n29854, 
        n28731, n56, n125, n512_adj_3592, n29461, n439_adj_3595, 
        n29460, n390, n463, n28730, n28729, n28728, n28727, n28726, 
        n366_adj_3596, n29459;
    wire [6:0]n7971;
    
    wire n560, n29672, n17_adj_3597, n28140, n28725, n28006, n177, 
        n29853, n28724, n487, n29671, n293_adj_3599, n29458, n414, 
        n29670, n220_adj_3600, n29457, n28723, n35_adj_3601, n104_adj_3602, 
        n15_adj_3603, n28139;
    wire [13:0]n8177;
    
    wire n29852, n13_adj_3605, n28138, n29851, n147_adj_3607, n29456, 
        n341, n29669, n5_adj_3608, n74_adj_3609, n268, n29668, n28722, 
        n29455, n28721, n28720, n29454, n29453, n195_adj_3610, n29667, 
        n29452, n29850, n29451, n29450, n29449, n53, n122_adj_3612;
    wire [7:0]n7961;
    
    wire n29666, n29849, n557, n29665, n29448, n29447, n484, n29664, 
        n29446, n29445, n29848, n28005, n29444, n411, n29663, 
        n11_adj_3613, n28137, n29847, n29443, n28004, n29846, n338, 
        n29662, n539, n29845, n29442, n265, n29661, n29441, n515_adj_3615, 
        n29440, n9_adj_3616, n28136, n28003, n442_adj_3618, n29439, 
        n466, n29844, n369_adj_3619, n29438, n296_adj_3620, n29437, 
        n192_adj_3621, n29660, n393, n29843, n50, n119_adj_3622, 
        n223_adj_3623, n29436;
    wire [8:0]n7950;
    
    wire n29659, n150_adj_3624, n29435, n29658, n7_adj_3625, n28135, 
        n554, n29657, n8_adj_3626, n77_adj_3627, n320, n29842, n481, 
        n29656, n5_adj_3628, n28134, n247, n29841, n174, n29840, 
        n408, n29655, n335, n29654, n32, n101, n262, n29653, 
        n189_adj_3630, n29652;
    wire [14:0]n8160;
    
    wire n29839, n29838, n47, n116_adj_3631;
    wire [9:0]n7938;
    
    wire n29651, n29650, n29649, n28002, n29837, n536, n551, n29648, 
        n478, n29647, n29836, n405, n29646, n29835, n332, n29645, 
        n3_adj_3634, n28133, n259, n29644, n186_adj_3635, n29643, 
        duty_23__N_3502, n29834, n44_adj_3637, n113_adj_3638, n29833, 
        n29832, n536_adj_3639, n29831, n463_adj_3640, n29830;
    wire [10:0]n7925;
    
    wire n29642, n29641, n390_adj_3641, n29829, n29640, n29639, 
        n317_adj_3642, n29828, n548_adj_3643, n29638, n244_adj_3644, 
        n29827, n171_adj_3645, n29826, n29_adj_3646, n98_adj_3647;
    wire [15:0]n8142;
    
    wire n29825, n475_adj_3648, n29637, n29824, n41_adj_3649, n28001, 
        n402_adj_3650, n29636, n39_adj_3651, n29823, n329_adj_3652, 
        n29635, n256_adj_3653, n29634, n183_adj_3654, n29633, n29822, 
        n41_adj_3655, n110_adj_3656;
    wire [11:0]n7911;
    
    wire n29632, n29631, n29821, n29630, n45_adj_3657, n29820, n29629, 
        n29628, n29819, n545_adj_3659, n29627, n29818, n472_adj_3660, 
        n29626, n43_adj_3661, n399_adj_3662, n29625, n326_adj_3663, 
        n29624, n28000, n29817, n533, n29816, n253_adj_3664, n29623, 
        n460, n29815, n180_adj_3665, n29622, n38_adj_3666, n107_adj_3667;
    wire [12:0]n7896;
    
    wire n29621, n29_adj_3668, n31_adj_3669, n37_adj_3670, n23_adj_3671, 
        n387, n29814, n314, n29813, n25_adj_3672, n241, n29812, 
        n35_adj_3673, n33_adj_3674, n9_adj_3675, n168, n29811, n17_adj_3676, 
        n19_adj_3677, n29620, n21_adj_3678, n26, n95, n29619;
    wire [16:0]n8123;
    
    wire n29810, n29809, n29808, n11_adj_3679, n13_adj_3681, n29807, 
        n15_adj_3682, n29618, n29806, n29805, n29804, n29803, n29617, 
        n29802, n29801, n29616, n530, n29800, n457, n29799, n384, 
        n29798, n311, n29797, n542_adj_3683, n29615, n238, n29796, 
        n27_adj_3684, n40727, n165, n29795, n23_adj_3685, n92, n40697, 
        \PID_CONTROLLER.integral_23__N_3451 , n12_adj_3686, n30, n469_adj_3687, 
        n29614, n40749, n41362, n396_adj_3688, n29613, n323_adj_3689, 
        n29612;
    wire [17:0]n8103;
    
    wire n29794, n29793, n29792, n41354, n250_adj_3690, n29611, 
        n29791, n29790, n42113, n41670, n42216, n6_adj_3691, n41909, 
        n41910, n16_adj_3692, n24_adj_3693, n40629, n8_adj_3694, n40627, 
        n41820, n41115, n4_adj_3695, n41907, n41908, n40689, n177_adj_3697, 
        n29610, n29789, n10_adj_3698, n40683, n42151, n41117, n35_adj_3699, 
        n104_adj_3700, n42284, n42285, n42271;
    wire [13:0]n7880;
    
    wire n29609, n40634, n29788, n42197, n41123, n42199, n29787, 
        n29786, n29608;
    wire [23:0]n257;
    
    wire n41_adj_3701, n39_adj_3703, n45_adj_3705, n43_adj_3706, n37_adj_3707, 
        n29_adj_3708, n31_adj_3709, n23_adj_3710, n25_adj_3711, n35_adj_3712, 
        n33_adj_3714, n11_adj_3715, n13_adj_3716, n15_adj_3717, n27_adj_3719, 
        n9_adj_3720, n17_adj_3721, n19_adj_3722, n21_adj_3724, n40605, 
        n40583, n12_adj_3725, n10_adj_3726, n30_adj_3727, n40623, 
        n41284, n41280, n42099, n41638, n42214, n16_adj_3728, n6_adj_3729, 
        n41860, n41861, n8_adj_3730, n24_adj_3731, n40460, n40453, 
        n41822, n41125, n40103, n4_adj_3732, n41836, n41837, n40522, 
        n40509, n42167, n41127, n42292, n42293, n42262, n40468, 
        n42050, n41133, n42201, n47_adj_3733, n89, n20_adj_3734, 
        n101_adj_3737, n32_adj_3738, n162, n29785, n29607, n28201, 
        n28200, n29606, n174_adj_3741, n247_adj_3743, n235, n320_adj_3744, 
        n29605, n308, n381, n393_adj_3745, n454, n29784, n466_adj_3746, 
        n29604, n29603, n527, n29783, n539_adj_3747, n29602, n29601, 
        n29782, n29600, n29781, n29780, n29599, n29779, n29598, 
        n28199, n29597, n29778;
    wire [14:0]n7863;
    
    wire n29596, n29595, n28198, n28197, n29594, n29593;
    wire [18:0]n8082;
    
    wire n29777, n29776, n28196, n29592, n28195, n29775, n28194, 
        n29591, n29590, n29774, n29589, n29588, n29773, n28193, 
        n28192, n29587, n29586, n28191, n28190, n29772, n29771, 
        n29770, n28189, n29769, n29585, n28188, n29768, n28187, 
        n28186, n28185, n29584, n29767, n29766, n29765, n29583, 
        n29764, n28184;
    wire [15:0]n7845;
    
    wire n29582, n29581, n29763, n28183, n28182, n29580, n29762, 
        n29579, n29578, n28181, n28180, n28179, n232, n29761, 
        n29577, n29576, n159, n29760, n29575, n28178, n28177, 
        n17_adj_3754, n86, n29574, n533_adj_3755, n29573, n28176;
    wire [19:0]n8060;
    
    wire n29759, n460_adj_3757, n29572, n29758, n387_adj_3758, n29571, 
        n314_adj_3759, n29570, n29757, n241_adj_3760, n29569, n168_adj_3761, 
        n29568, n29756, n26_adj_3762, n95_adj_3763, n29755, n17_adj_3764, 
        n9_adj_3765, n11_adj_3766, n40517, n40350, n44041, n41560, 
        n40987, n44023, n40943;
    wire [16:0]n7826;
    
    wire n29567, n41514, n44017, n40812, n40833, n16_adj_3767, n40753, 
        n8_adj_3768, n24_adj_3769, n40873, n41468, n41452, n42133, 
        n41722, n42220, n41037, n44010, n41502, n44005, n12_adj_3770, 
        n40899, n44028, n10_adj_3771, n30_adj_3772, n41766, n40922, 
        n44008, n41760, n44034, n42143, n43999, n42305, n43996, 
        n16_adj_3773, n40875, n24_adj_3774, n6_adj_3775, n41923, n41924, 
        n40877, n8_adj_3776, n43994, n41816, n41095, n4_adj_3777, 
        n41915, n41916, n12_adj_3778, n28175, n40797, n10_adj_3780, 
        n29754, n29566, n29565, n29564, n30_adj_3781, n29563, n29753, 
        n29562, n40803, n42149, n41107, n28174, n29561, n42282, 
        n29752, n29560, n42283, n42273, n29559, n29751, n29558, 
        n530_adj_3783, n29557, n6_adj_3784, n41917, n29750, n457_adj_3785, 
        n29556, n384_adj_3786, n29555, n41918, n311_adj_3787, n29554, 
        n28173, n40757, n41818, n29749, n238_adj_3789, n29553, n41105, 
        n165_adj_3790, n29552, n40759, n42193, n41113, n28172, n42195, 
        n29748, n23_adj_3792, n92_adj_3793, n4_adj_3794;
    wire [17:0]n7806;
    
    wire n29551, n28171, n29747, n29550, n41921, n521_adj_3796, 
        n29746, n29549, n29548, n41922, n28170, n40901, n28169, 
        n28168, n448_adj_3800, n29745, n29547, n42147, n375_adj_3801, 
        n29744, n29546, n41097, n28167, n42280, n29545, n42281, 
        n29544, n302_adj_3803, n29743, n42277, n40884, n42189, n41103, 
        \PID_CONTROLLER.integral_23__N_3453 , n229_adj_3804, n29742, n29543, 
        n42191, n29542, n156_adj_3805, n29741, n29541, n14_adj_3806, 
        n83_adj_3807, n527_adj_3808, n29540, n29740, n454_adj_3809, 
        n29539, n29739, n381_adj_3810, n29538, n28166, n29738, n308_adj_3812, 
        n29537, n29737, n235_adj_3813, n29536, n29736, n162_adj_3814, 
        n29535, n20_adj_3815, n89_adj_3816, n29735, n29534, n29533, 
        n28022, n28165, n29532, n28164, n29734, n29531, n29530, 
        n29733, n29529, n29732, n29528, n29527, n29526, n29731, 
        n29525, n29524, n28021, n29730, n29523, n524_adj_3819, n29522, 
        n29729, n451_adj_3820, n29521, n28020, n28163, n378_adj_3822, 
        n29520, n29728, n28162, n305_adj_3824, n29519, n232_adj_3825, 
        n29518, n29727, n159_adj_3826, n29517, n28019, n17_adj_3827, 
        n86_adj_3828, n518_adj_3829, n29726, n29516, n28161, n29515, 
        n445_adj_3831, n29725, n29514, n40149, n29513, n372_adj_3832, 
        n29724, n28160, n29512, n28159, n28018, n299_adj_3835, n29723, 
        n29511, n28158, n28017, n29510, n28157, n226_adj_3838, n29722, 
        n29509;
    wire [5:0]n8277;
    
    wire n36243, n490_adj_3839, n29920;
    wire [4:0]n8285;
    
    wire n417_adj_3840, n29919, n344_adj_3841, n29918, n271_adj_3842, 
        n29917, n198_adj_3843, n29916, n56_adj_3844, n125_adj_3845;
    wire [6:0]n8268;
    
    wire n560_adj_3846, n29915, n487_adj_3847, n29914, n414_adj_3848, 
        n29913, n341_adj_3849, n29912, n29508, n268_adj_3851, n29911, 
        n195_adj_3852, n29910, n53_adj_3853, n122_adj_3854;
    wire [7:0]n8258;
    
    wire n29909, n557_adj_3855, n29908, n153_adj_3856, n29721, n484_adj_3857, 
        n29907, n411_adj_3858, n29906, n338_adj_3859, n29905, n265_adj_3860, 
        n29904, n29507, n192_adj_3861, n29903, n50_adj_3862, n119_adj_3863, 
        n29902, n29901, n554_adj_3864, n29900, n481_adj_3865, n29899, 
        n408_adj_3866, n29898, n335_adj_3867, n29897, n262_adj_3868, 
        n29896, n189_adj_3869, n29895, n47_adj_3870, n116_adj_3871, 
        n29894, n29506, n29893, n29892, n551_adj_3872, n29891, n478_adj_3873, 
        n29890, n405_adj_3874, n29889, n332_adj_3876, n29888, n11_adj_3877, 
        n80_adj_3878, n259_adj_3879, n27655;
    wire [1:0]n8006;
    
    wire n4_adj_3880;
    wire [3:0]n8292;
    
    wire n6_adj_3881;
    wire [2:0]n8298;
    
    wire n27791, n4_adj_3882, n27825;
    wire [1:0]n8303;
    
    wire n4_adj_3883, n12_adj_3884, n8_adj_3885, n27748, n11_adj_3886, 
        n6_adj_3887, n27850, n18_adj_3888, n13_adj_3889, n4_adj_3890, 
        n27578;
    
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n28156));
    SB_CARRY add_3692_9 (.CI(n29504), .I0(n7785[6]), .I1(GND_net), .CO(n29505));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3891[23]), 
            .I3(n28155), .O(\PID_CONTROLLER.integral_23__N_3454 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_3891[22]), .I3(n28154), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3692_8_lut (.I0(GND_net), .I1(n7785[5]), .I2(n521), .I3(n29503), 
            .O(n7763[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_8 (.CI(n29503), .I0(n7785[5]), .I1(n521), .CO(n29504));
    SB_LUT4 add_3692_7_lut (.I0(GND_net), .I1(n7785[4]), .I2(n448), .I3(n29502), 
            .O(n7763[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_7 (.CI(n29502), .I0(n7785[4]), .I1(n448), .CO(n29503));
    SB_CARRY mult_11_add_1225_23 (.CI(n29719), .I0(n8013[20]), .I1(GND_net), 
            .CO(n29720));
    SB_LUT4 add_3692_6_lut (.I0(GND_net), .I1(n7785[3]), .I2(n375), .I3(n29501), 
            .O(n7763[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_6 (.CI(n29501), .I0(n7785[3]), .I1(n375), .CO(n29502));
    SB_CARRY unary_minus_5_add_3_24 (.CI(n28154), .I0(GND_net), .I1(n1_adj_3891[22]), 
            .CO(n28155));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n8013[19]), .I2(GND_net), 
            .I3(n29718), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n29718), .I0(n8013[19]), .I1(GND_net), 
            .CO(n29719));
    SB_LUT4 add_3692_5_lut (.I0(GND_net), .I1(n7785[2]), .I2(n302), .I3(n29500), 
            .O(n7763[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_3891[21]), .I3(n28153), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n28153), .I0(GND_net), .I1(n1_adj_3891[21]), 
            .CO(n28154));
    SB_CARRY add_3692_5 (.CI(n29500), .I0(n7785[2]), .I1(n302), .CO(n29501));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n8013[18]), .I2(GND_net), 
            .I3(n29717), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_3_lut (.I0(GND_net), .I1(n8247[0]), .I2(n186), .I3(n29886), 
            .O(n8235[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n29717), .I0(n8013[18]), .I1(GND_net), 
            .CO(n29718));
    SB_LUT4 add_3692_4_lut (.I0(GND_net), .I1(n7785[1]), .I2(n229), .I3(n29499), 
            .O(n7763[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n8013[17]), .I2(GND_net), 
            .I3(n29716), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_4 (.CI(n29499), .I0(n7785[1]), .I1(n229), .CO(n29500));
    SB_CARRY add_3724_3 (.CI(n29886), .I0(n8247[0]), .I1(n186), .CO(n29887));
    SB_CARRY mult_11_add_1225_20 (.CI(n29716), .I0(n8013[17]), .I1(GND_net), 
            .CO(n29717));
    SB_LUT4 add_3692_3_lut (.I0(GND_net), .I1(n7785[0]), .I2(n156), .I3(n29498), 
            .O(n7763[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_3 (.CI(n29498), .I0(n7785[0]), .I1(n156), .CO(n29499));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n8013[16]), .I2(GND_net), 
            .I3(n29715), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n7763[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n29498));
    SB_CARRY add_636_18 (.CI(n28015), .I0(n2996[16]), .I1(n3021[16]), 
            .CO(n28016));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_3891[20]), .I3(n28152), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n28152), .I0(GND_net), .I1(n1_adj_3891[20]), 
            .CO(n28153));
    SB_LUT4 add_3724_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n8235[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n29715), .I0(n8013[16]), .I1(GND_net), 
            .CO(n29716));
    SB_LUT4 add_3691_22_lut (.I0(GND_net), .I1(n7763[19]), .I2(GND_net), 
            .I3(n29497), .O(n7740[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n8013[15]), .I2(GND_net), 
            .I3(n29714), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3691_21_lut (.I0(GND_net), .I1(n7763[18]), .I2(GND_net), 
            .I3(n29496), .O(n7740[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_636_17_lut (.I0(GND_net), .I1(n2996[15]), .I2(n3021[15]), 
            .I3(n28014), .O(duty_23__N_3478[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n29886));
    SB_CARRY mult_11_add_1225_18 (.CI(n29714), .I0(n8013[15]), .I1(GND_net), 
            .CO(n29715));
    SB_CARRY add_3691_21 (.CI(n29496), .I0(n7763[18]), .I1(GND_net), .CO(n29497));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_3891[19]), .I3(n28151), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n28151), .I0(GND_net), .I1(n1_adj_3891[19]), 
            .CO(n28152));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n8013[14]), .I2(GND_net), 
            .I3(n29713), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3691_20_lut (.I0(GND_net), .I1(n7763[17]), .I2(GND_net), 
            .I3(n29495), .O(n7740[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_17 (.CI(n28014), .I0(n2996[15]), .I1(n3021[15]), 
            .CO(n28015));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_3891[18]), .I3(n28150), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n28150), .I0(GND_net), .I1(n1_adj_3891[18]), 
            .CO(n28151));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_3891[17]), .I3(n28149), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n28149), .I0(GND_net), .I1(n1_adj_3891[17]), 
            .CO(n28150));
    SB_LUT4 add_3723_12_lut (.I0(GND_net), .I1(n8235[9]), .I2(GND_net), 
            .I3(n29885), .O(n8222[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n29713), .I0(n8013[14]), .I1(GND_net), 
            .CO(n29714));
    SB_CARRY add_3691_20 (.CI(n29495), .I0(n7763[17]), .I1(GND_net), .CO(n29496));
    SB_LUT4 add_3691_19_lut (.I0(GND_net), .I1(n7763[16]), .I2(GND_net), 
            .I3(n29494), .O(n7740[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n8013[13]), .I2(GND_net), 
            .I3(n29712), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_19 (.CI(n29494), .I0(n7763[16]), .I1(GND_net), .CO(n29495));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_3891[16]), .I3(n28148), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3723_11_lut (.I0(GND_net), .I1(n8235[8]), .I2(GND_net), 
            .I3(n29884), .O(n8222[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n29712), .I0(n8013[13]), .I1(GND_net), 
            .CO(n29713));
    SB_LUT4 add_3691_18_lut (.I0(GND_net), .I1(n7763[15]), .I2(GND_net), 
            .I3(n29493), .O(n7740[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n8013[12]), .I2(GND_net), 
            .I3(n29711), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_18 (.CI(n29493), .I0(n7763[15]), .I1(GND_net), .CO(n29494));
    SB_CARRY add_3723_11 (.CI(n29884), .I0(n8235[8]), .I1(GND_net), .CO(n29885));
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_636_16_lut (.I0(GND_net), .I1(n2996[14]), .I2(n3021[14]), 
            .I3(n28013), .O(duty_23__N_3478[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n29711), .I0(n8013[12]), .I1(GND_net), 
            .CO(n29712));
    SB_LUT4 add_3723_10_lut (.I0(GND_net), .I1(n8235[7]), .I2(GND_net), 
            .I3(n29883), .O(n8222[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n8013[11]), .I2(GND_net), 
            .I3(n29710), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_10 (.CI(n29883), .I0(n8235[7]), .I1(GND_net), .CO(n29884));
    SB_LUT4 add_3723_9_lut (.I0(GND_net), .I1(n8235[6]), .I2(GND_net), 
            .I3(n29882), .O(n8222[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n29710), .I0(n8013[11]), .I1(GND_net), 
            .CO(n29711));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n8013[10]), .I2(GND_net), 
            .I3(n29709), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_9 (.CI(n29882), .I0(n8235[6]), .I1(GND_net), .CO(n29883));
    SB_LUT4 add_3691_17_lut (.I0(GND_net), .I1(n7763[14]), .I2(GND_net), 
            .I3(n29492), .O(n7740[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n29709), .I0(n8013[10]), .I1(GND_net), 
            .CO(n29710));
    SB_LUT4 add_3723_8_lut (.I0(GND_net), .I1(n8235[5]), .I2(n548), .I3(n29881), 
            .O(n8222[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_8 (.CI(n29881), .I0(n8235[5]), .I1(n548), .CO(n29882));
    SB_CARRY unary_minus_5_add_3_18 (.CI(n28148), .I0(GND_net), .I1(n1_adj_3891[16]), 
            .CO(n28149));
    SB_LUT4 i2_4_lut (.I0(n4_adj_3565), .I1(\Kp[3] ), .I2(n8001[1]), .I3(\PID_CONTROLLER.err [19]), 
            .O(n7995[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_844 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_844.LUT_INIT = 16'h9c50;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[4]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23011_4_lut (.I0(n7995[2]), .I1(\Kp[4] ), .I2(n6_adj_3566), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_3567));   // verilog/motorControl.v(42[17:23])
    defparam i23011_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11));   // verilog/motorControl.v(42[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23042_4_lut (.I0(n8001[1]), .I1(\Kp[3] ), .I2(n4_adj_3565), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_3568));   // verilog/motorControl.v(42[17:23])
    defparam i23042_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[5]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23077_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n27680));   // verilog/motorControl.v(42[17:23])
    defparam i23077_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3723_7_lut (.I0(GND_net), .I1(n8235[4]), .I2(n475), .I3(n29880), 
            .O(n8222[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n8013[9]), .I2(GND_net), 
            .I3(n29708), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_17 (.CI(n29492), .I0(n7763[14]), .I1(GND_net), .CO(n29493));
    SB_LUT4 i8_4_lut (.I0(n6_adj_3568), .I1(n11), .I2(n8_adj_3567), .I3(n12), 
            .O(n18));   // verilog/motorControl.v(42[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3691_16_lut (.I0(GND_net), .I1(n7763[13]), .I2(GND_net), 
            .I3(n29491), .O(n7740[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13));   // verilog/motorControl.v(42[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY mult_11_add_1225_12 (.CI(n29708), .I0(n8013[9]), .I1(GND_net), 
            .CO(n29709));
    SB_CARRY add_3691_16 (.CI(n29491), .I0(n7763[13]), .I1(GND_net), .CO(n29492));
    SB_LUT4 add_3691_15_lut (.I0(GND_net), .I1(n7763[12]), .I2(GND_net), 
            .I3(n29490), .O(n7740[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut (.I0(n13), .I1(n18), .I2(n27680), .I3(n4_adj_3569), 
            .O(n36676));   // verilog/motorControl.v(42[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_3891[15]), .I3(n28147), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n8013[8]), .I2(GND_net), 
            .I3(n29707), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_15 (.CI(n29490), .I0(n7763[12]), .I1(GND_net), .CO(n29491));
    SB_LUT4 add_3691_14_lut (.I0(GND_net), .I1(n7763[11]), .I2(GND_net), 
            .I3(n29489), .O(n7740[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_7 (.CI(n29880), .I0(n8235[4]), .I1(n475), .CO(n29881));
    SB_CARRY mult_11_add_1225_11 (.CI(n29707), .I0(n8013[8]), .I1(GND_net), 
            .CO(n29708));
    SB_CARRY add_3691_14 (.CI(n29489), .I0(n7763[11]), .I1(GND_net), .CO(n29490));
    SB_LUT4 add_3691_13_lut (.I0(GND_net), .I1(n7763[10]), .I2(GND_net), 
            .I3(n29488), .O(n7740[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n8013[7]), .I2(GND_net), 
            .I3(n29706), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3723_6_lut (.I0(GND_net), .I1(n8235[3]), .I2(n402), .I3(n29879), 
            .O(n8222[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_6 (.CI(n29879), .I0(n8235[3]), .I1(n402), .CO(n29880));
    SB_CARRY mult_11_add_1225_10 (.CI(n29706), .I0(n8013[7]), .I1(GND_net), 
            .CO(n29707));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n8013[6]), .I2(GND_net), 
            .I3(n29705), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n29705), .I0(n8013[6]), .I1(GND_net), 
            .CO(n29706));
    SB_LUT4 add_3723_5_lut (.I0(GND_net), .I1(n8235[2]), .I2(n329), .I3(n29878), 
            .O(n8222[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_5 (.CI(n29878), .I0(n8235[2]), .I1(n329), .CO(n29879));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n8013[5]), .I2(n512), 
            .I3(n29704), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n29704), .I0(n8013[5]), .I1(n512), 
            .CO(n29705));
    SB_LUT4 add_3723_4_lut (.I0(GND_net), .I1(n8235[1]), .I2(n256), .I3(n29877), 
            .O(n8222[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3570));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3723_4 (.CI(n29877), .I0(n8235[1]), .I1(n256), .CO(n29878));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n8013[4]), .I2(n439), 
            .I3(n29703), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i9_3_lut (.I0(n155[8]), .I1(PWMLimit[8]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i9_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23023_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n27621));   // verilog/motorControl.v(42[17:23])
    defparam i23023_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[9]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3723_3_lut (.I0(GND_net), .I1(n8235[0]), .I2(n183_adj_3572), 
            .I3(n29876), .O(n8222[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_13 (.CI(n29488), .I0(n7763[10]), .I1(GND_net), .CO(n29489));
    SB_LUT4 mux_634_i10_3_lut (.I0(n155[9]), .I1(PWMLimit[9]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i10_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3723_3 (.CI(n29876), .I0(n8235[0]), .I1(n183_adj_3572), 
            .CO(n29877));
    SB_LUT4 add_3723_2_lut (.I0(GND_net), .I1(n41_adj_3573), .I2(n110), 
            .I3(GND_net), .O(n8222[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3723_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n29703), .I0(n8013[4]), .I1(n439), 
            .CO(n29704));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n8013[3]), .I2(n366), 
            .I3(n29702), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3723_2 (.CI(GND_net), .I0(n41_adj_3573), .I1(n110), .CO(n29876));
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3722_13_lut (.I0(GND_net), .I1(n8222[10]), .I2(GND_net), 
            .I3(n29875), .O(n8208[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_12_lut (.I0(GND_net), .I1(n8222[9]), .I2(GND_net), 
            .I3(n29874), .O(n8208[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_12 (.CI(n29874), .I0(n8222[9]), .I1(GND_net), .CO(n29875));
    SB_LUT4 add_3722_11_lut (.I0(GND_net), .I1(n8222[8]), .I2(GND_net), 
            .I3(n29873), .O(n8208[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n29702), .I0(n8013[3]), .I1(n366), 
            .CO(n29703));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n8013[2]), .I2(n293), 
            .I3(n29701), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n29701), .I0(n8013[2]), .I1(n293), 
            .CO(n29702));
    SB_CARRY add_3722_11 (.CI(n29873), .I0(n8222[8]), .I1(GND_net), .CO(n29874));
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_636_16 (.CI(n28013), .I0(n2996[14]), .I1(n3021[14]), 
            .CO(n28014));
    SB_LUT4 add_3722_10_lut (.I0(GND_net), .I1(n8222[7]), .I2(GND_net), 
            .I3(n29872), .O(n8208[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n8013[1]), .I2(n220), 
            .I3(n29700), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3691_12_lut (.I0(GND_net), .I1(n7763[9]), .I2(GND_net), 
            .I3(n29487), .O(n7740[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n29700), .I0(n8013[1]), .I1(n220), 
            .CO(n29701));
    SB_CARRY add_3691_12 (.CI(n29487), .I0(n7763[9]), .I1(GND_net), .CO(n29488));
    SB_CARRY add_3722_10 (.CI(n29872), .I0(n8222[7]), .I1(GND_net), .CO(n29873));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n8013[0]), .I2(n147), 
            .I3(n29699), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3691_11_lut (.I0(GND_net), .I1(n7763[8]), .I2(GND_net), 
            .I3(n29486), .O(n7740[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n29699), .I0(n8013[0]), .I1(n147), 
            .CO(n29700));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n28147), .I0(GND_net), .I1(n1_adj_3891[15]), 
            .CO(n28148));
    SB_LUT4 add_636_15_lut (.I0(GND_net), .I1(n2996[13]), .I2(n3021[13]), 
            .I3(n28012), .O(duty_23__N_3478[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_11 (.CI(n29486), .I0(n7763[8]), .I1(GND_net), .CO(n29487));
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3691_10_lut (.I0(GND_net), .I1(n7763[7]), .I2(GND_net), 
            .I3(n29485), .O(n7740[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_634_i11_3_lut (.I0(n155[10]), .I1(PWMLimit[10]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i11_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3691_10 (.CI(n29485), .I0(n7763[7]), .I1(GND_net), .CO(n29486));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_3891[14]), .I3(n28146), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3355[0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_3575), .I2(n74), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_3575), .I1(n74), 
            .CO(n29699));
    SB_LUT4 add_3722_9_lut (.I0(GND_net), .I1(n8222[6]), .I2(GND_net), 
            .I3(n29871), .O(n8208[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_9 (.CI(n29871), .I0(n8222[6]), .I1(GND_net), .CO(n29872));
    SB_LUT4 add_3712_23_lut (.I0(GND_net), .I1(n8037[20]), .I2(GND_net), 
            .I3(n29698), .O(n8013[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_15 (.CI(n28012), .I0(n2996[13]), .I1(n3021[13]), 
            .CO(n28013));
    SB_LUT4 add_3722_8_lut (.I0(GND_net), .I1(n8222[5]), .I2(n545), .I3(n29870), 
            .O(n8208[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3712_22_lut (.I0(GND_net), .I1(n8037[19]), .I2(GND_net), 
            .I3(n29697), .O(n8013[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3691_9_lut (.I0(GND_net), .I1(n7763[6]), .I2(GND_net), 
            .I3(n29484), .O(n7740[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n28146), .I0(GND_net), .I1(n1_adj_3891[14]), 
            .CO(n28147));
    SB_CARRY add_3712_22 (.CI(n29697), .I0(n8037[19]), .I1(GND_net), .CO(n29698));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_3891[13]), .I3(n28145), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n28145), .I0(GND_net), .I1(n1_adj_3891[13]), 
            .CO(n28146));
    SB_CARRY add_3722_8 (.CI(n29870), .I0(n8222[5]), .I1(n545), .CO(n29871));
    SB_LUT4 add_3722_7_lut (.I0(GND_net), .I1(n8222[4]), .I2(n472), .I3(n29869), 
            .O(n8208[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3712_21_lut (.I0(GND_net), .I1(n8037[18]), .I2(GND_net), 
            .I3(n29696), .O(n8013[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_21 (.CI(n29696), .I0(n8037[18]), .I1(GND_net), .CO(n29697));
    SB_CARRY add_3691_9 (.CI(n29484), .I0(n7763[6]), .I1(GND_net), .CO(n29485));
    SB_LUT4 add_3712_20_lut (.I0(GND_net), .I1(n8037[17]), .I2(GND_net), 
            .I3(n29695), .O(n8013[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_7 (.CI(n29869), .I0(n8222[4]), .I1(n472), .CO(n29870));
    SB_LUT4 add_3691_8_lut (.I0(GND_net), .I1(n7763[5]), .I2(n518), .I3(n29483), 
            .O(n7740[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_636_14_lut (.I0(GND_net), .I1(n2996[12]), .I2(n3021[12]), 
            .I3(n28011), .O(duty_23__N_3478[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_20 (.CI(n29695), .I0(n8037[17]), .I1(GND_net), .CO(n29696));
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[10]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_636_14 (.CI(n28011), .I0(n2996[12]), .I1(n3021[12]), 
            .CO(n28012));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_3891[12]), .I3(n28144), .O(n25_adj_3577)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3691_8 (.CI(n29483), .I0(n7763[5]), .I1(n518), .CO(n29484));
    SB_LUT4 add_3691_7_lut (.I0(GND_net), .I1(n7763[4]), .I2(n445), .I3(n29482), 
            .O(n7740[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3712_19_lut (.I0(GND_net), .I1(n8037[16]), .I2(GND_net), 
            .I3(n29694), .O(n8013[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_6_lut (.I0(GND_net), .I1(n8222[3]), .I2(n399), .I3(n29868), 
            .O(n8208[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_7 (.CI(n29482), .I0(n7763[4]), .I1(n445), .CO(n29483));
    SB_CARRY add_3712_19 (.CI(n29694), .I0(n8037[16]), .I1(GND_net), .CO(n29695));
    SB_LUT4 add_3691_6_lut (.I0(GND_net), .I1(n7763[3]), .I2(n372), .I3(n29481), 
            .O(n7740[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_6 (.CI(n29481), .I0(n7763[3]), .I1(n372), .CO(n29482));
    SB_LUT4 add_3712_18_lut (.I0(GND_net), .I1(n8037[15]), .I2(GND_net), 
            .I3(n29693), .O(n8013[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19558_1_lut (.I0(n256_adj_3571), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24213));   // verilog/motorControl.v(46[19:35])
    defparam i19558_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3691_5_lut (.I0(GND_net), .I1(n7763[2]), .I2(n299), .I3(n29480), 
            .O(n7740[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_636_13_lut (.I0(GND_net), .I1(n2996[11]), .I2(n3021[11]), 
            .I3(n28010), .O(duty_23__N_3478[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3712_18 (.CI(n29693), .I0(n8037[15]), .I1(GND_net), .CO(n29694));
    SB_LUT4 add_3712_17_lut (.I0(GND_net), .I1(n8037[14]), .I2(GND_net), 
            .I3(n29692), .O(n8013[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3579));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3712_17 (.CI(n29692), .I0(n8037[14]), .I1(GND_net), .CO(n29693));
    SB_LUT4 add_3712_16_lut (.I0(GND_net), .I1(n8037[13]), .I2(GND_net), 
            .I3(n29691), .O(n8013[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_16 (.CI(n29691), .I0(n8037[13]), .I1(GND_net), .CO(n29692));
    SB_LUT4 add_3712_15_lut (.I0(GND_net), .I1(n8037[12]), .I2(GND_net), 
            .I3(n29690), .O(n8013[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_15 (.CI(n29690), .I0(n8037[12]), .I1(GND_net), .CO(n29691));
    SB_LUT4 add_3712_14_lut (.I0(GND_net), .I1(n8037[11]), .I2(GND_net), 
            .I3(n29689), .O(n8013[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n28144), .I0(GND_net), .I1(n1_adj_3891[12]), 
            .CO(n28145));
    SB_CARRY add_3712_14 (.CI(n29689), .I0(n8037[11]), .I1(GND_net), .CO(n29690));
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3722_6 (.CI(n29868), .I0(n8222[3]), .I1(n399), .CO(n29869));
    SB_LUT4 add_3712_13_lut (.I0(GND_net), .I1(n8037[10]), .I2(GND_net), 
            .I3(n29688), .O(n8013[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_13 (.CI(n29688), .I0(n8037[10]), .I1(GND_net), .CO(n29689));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_3891[11]), .I3(n28143), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3691_5 (.CI(n29480), .I0(n7763[2]), .I1(n299), .CO(n29481));
    SB_CARRY add_636_13 (.CI(n28010), .I0(n2996[11]), .I1(n3021[11]), 
            .CO(n28011));
    SB_LUT4 add_3691_4_lut (.I0(GND_net), .I1(n7763[1]), .I2(n226), .I3(n29479), 
            .O(n7740[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3691_4 (.CI(n29479), .I0(n7763[1]), .I1(n226), .CO(n29480));
    SB_LUT4 add_3712_12_lut (.I0(GND_net), .I1(n8037[9]), .I2(GND_net), 
            .I3(n29687), .O(n8013[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3691_3_lut (.I0(GND_net), .I1(n7763[0]), .I2(n153), .I3(n29478), 
            .O(n7740[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_12 (.CI(n29687), .I0(n8037[9]), .I1(GND_net), .CO(n29688));
    SB_CARRY add_3691_3 (.CI(n29478), .I0(n7763[0]), .I1(n153), .CO(n29479));
    SB_LUT4 add_3691_2_lut (.I0(GND_net), .I1(n11_adj_3579), .I2(n80), 
            .I3(GND_net), .O(n7740[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3691_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_5_lut (.I0(GND_net), .I1(n8222[2]), .I2(n326), .I3(n29867), 
            .O(n8208[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3712_11_lut (.I0(GND_net), .I1(n8037[8]), .I2(GND_net), 
            .I3(n29686), .O(n8013[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_5 (.CI(n29867), .I0(n8222[2]), .I1(n326), .CO(n29868));
    SB_CARRY add_3712_11 (.CI(n29686), .I0(n8037[8]), .I1(GND_net), .CO(n29687));
    SB_LUT4 add_3722_4_lut (.I0(GND_net), .I1(n8222[1]), .I2(n253), .I3(n29866), 
            .O(n8208[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n28143), .I0(GND_net), .I1(n1_adj_3891[11]), 
            .CO(n28144));
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3691_2 (.CI(GND_net), .I0(n11_adj_3579), .I1(n80), .CO(n29478));
    SB_LUT4 add_3712_10_lut (.I0(GND_net), .I1(n8037[7]), .I2(GND_net), 
            .I3(n29685), .O(n8013[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_10 (.CI(n29685), .I0(n8037[7]), .I1(GND_net), .CO(n29686));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n7716[21]), 
            .I2(GND_net), .I3(n29477), .O(n6169[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n24213), .I1(n7716[20]), .I2(GND_net), 
            .I3(n29476), .O(n2996[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3722_4 (.CI(n29866), .I0(n8222[1]), .I1(n253), .CO(n29867));
    SB_LUT4 add_3712_9_lut (.I0(GND_net), .I1(n8037[6]), .I2(GND_net), 
            .I3(n29684), .O(n8013[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3722_3_lut (.I0(GND_net), .I1(n8222[0]), .I2(n180), .I3(n29865), 
            .O(n8208[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3722_3 (.CI(n29865), .I0(n8222[0]), .I1(n180), .CO(n29866));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_3891[10]), .I3(n28142), .O(n21_adj_3581)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_636_12_lut (.I0(GND_net), .I1(n2996[10]), .I2(n3021[10]), 
            .I3(n28009), .O(duty_23__N_3478[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n29476), .I0(n7716[20]), .I1(GND_net), 
            .CO(n29477));
    SB_LUT4 add_3722_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n8208[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3722_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[11]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_634_i12_3_lut (.I0(n155[11]), .I1(PWMLimit[11]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i12_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3722_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n29865));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n28742), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_14_lut (.I0(GND_net), .I1(n8208[11]), .I2(GND_net), 
            .I3(n29864), .O(n8193[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3712_9 (.CI(n29684), .I0(n8037[6]), .I1(GND_net), .CO(n29685));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n28741), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_13_lut (.I0(GND_net), .I1(n8208[10]), .I2(GND_net), 
            .I3(n29863), .O(n8193[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_13 (.CI(n29863), .I0(n8208[10]), .I1(GND_net), .CO(n29864));
    SB_LUT4 add_3712_8_lut (.I0(GND_net), .I1(n8037[5]), .I2(n515), .I3(n29683), 
            .O(n8013[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_24  (.CI(n28741), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n28742));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n24213), .I1(n7716[19]), .I2(GND_net), 
            .I3(n29475), .O(n2996[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n28740), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_636_12 (.CI(n28009), .I0(n2996[10]), .I1(n3021[10]), 
            .CO(n28010));
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_23  (.CI(n28740), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n28741));
    SB_LUT4 add_636_11_lut (.I0(GND_net), .I1(n2996[9]), .I2(n3021[9]), 
            .I3(n28008), .O(duty_23__N_3478[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n28739), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_22  (.CI(n28739), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n28740));
    SB_CARRY add_3712_8 (.CI(n29683), .I0(n8037[5]), .I1(n515), .CO(n29684));
    SB_LUT4 add_3721_12_lut (.I0(GND_net), .I1(n8208[9]), .I2(GND_net), 
            .I3(n29862), .O(n8193[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_12 (.CI(n29862), .I0(n8208[9]), .I1(GND_net), .CO(n29863));
    SB_CARRY mult_10_add_1225_22 (.CI(n29475), .I0(n7716[19]), .I1(GND_net), 
            .CO(n29476));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n24213), .I1(n7716[18]), .I2(GND_net), 
            .I3(n29474), .O(n2996[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_21 (.CI(n29474), .I0(n7716[18]), .I1(GND_net), 
            .CO(n29475));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n24213), .I1(n7716[17]), .I2(GND_net), 
            .I3(n29473), .O(n2996[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_20 (.CI(n29473), .I0(n7716[17]), .I1(GND_net), 
            .CO(n29474));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n28142), .I0(GND_net), .I1(n1_adj_3891[10]), 
            .CO(n28143));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n24213), .I1(n7716[16]), .I2(GND_net), 
            .I3(n29472), .O(n2996[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n28738), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_21  (.CI(n28738), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n28739));
    SB_CARRY add_636_11 (.CI(n28008), .I0(n2996[9]), .I1(n3021[9]), .CO(n28009));
    SB_CARRY mult_10_add_1225_19 (.CI(n29472), .I0(n7716[16]), .I1(GND_net), 
            .CO(n29473));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n24213), .I1(n7716[15]), .I2(GND_net), 
            .I3(n29471), .O(n2996[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_18 (.CI(n29471), .I0(n7716[15]), .I1(GND_net), 
            .CO(n29472));
    SB_LUT4 add_3721_11_lut (.I0(GND_net), .I1(n8208[8]), .I2(GND_net), 
            .I3(n29861), .O(n8193[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_3891[9]), .I3(n28141), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[6]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n28737), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_20  (.CI(n28737), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n28738));
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3584));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3712_7_lut (.I0(GND_net), .I1(n8037[4]), .I2(n442), .I3(n29682), 
            .O(n8013[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n24213), .I1(n7716[14]), .I2(GND_net), 
            .I3(n29470), .O(n2996[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3712_7 (.CI(n29682), .I0(n8037[4]), .I1(n442), .CO(n29683));
    SB_LUT4 add_3712_6_lut (.I0(GND_net), .I1(n8037[3]), .I2(n369), .I3(n29681), 
            .O(n8013[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n29470), .I0(n7716[14]), .I1(GND_net), 
            .CO(n29471));
    SB_CARRY add_3721_11 (.CI(n29861), .I0(n8208[8]), .I1(GND_net), .CO(n29862));
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3712_6 (.CI(n29681), .I0(n8037[3]), .I1(n369), .CO(n29682));
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[7]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3721_10_lut (.I0(GND_net), .I1(n8208[7]), .I2(GND_net), 
            .I3(n29860), .O(n8193[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3712_5_lut (.I0(GND_net), .I1(n8037[2]), .I2(n296), .I3(n29680), 
            .O(n8013[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_5 (.CI(n29680), .I0(n8037[2]), .I1(n296), .CO(n29681));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n24213), .I1(n7716[13]), .I2(GND_net), 
            .I3(n29469), .O(n2996[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_636_10_lut (.I0(GND_net), .I1(n2996[8]), .I2(n3021[8]), 
            .I3(n28007), .O(duty_23__N_3478[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_10 (.CI(n29860), .I0(n8208[7]), .I1(GND_net), .CO(n29861));
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[8]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[9]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n28141), .I0(GND_net), .I1(n1_adj_3891[9]), 
            .CO(n28142));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n28736), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[10]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_19  (.CI(n28736), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n28737));
    SB_CARRY mult_10_add_1225_16 (.CI(n29469), .I0(n7716[13]), .I1(GND_net), 
            .CO(n29470));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n24213), .I1(n7716[12]), .I2(GND_net), 
            .I3(n29468), .O(n2996[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n28735), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n29468), .I0(n7716[12]), .I1(GND_net), 
            .CO(n29469));
    SB_LUT4 add_3712_4_lut (.I0(GND_net), .I1(n8037[1]), .I2(n223), .I3(n29679), 
            .O(n8013[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_4 (.CI(n29679), .I0(n8037[1]), .I1(n223), .CO(n29680));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n24213), .I1(n7716[11]), .I2(GND_net), 
            .I3(n29467), .O(n2996[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3712_3_lut (.I0(GND_net), .I1(n8037[0]), .I2(n150), .I3(n29678), 
            .O(n8013[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_18  (.CI(n28735), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n28736));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n28734), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_9_lut (.I0(GND_net), .I1(n8208[6]), .I2(GND_net), 
            .I3(n29859), .O(n8193[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3712_3 (.CI(n29678), .I0(n8037[0]), .I1(n150), .CO(n29679));
    SB_CARRY mult_10_add_1225_14 (.CI(n29467), .I0(n7716[11]), .I1(GND_net), 
            .CO(n29468));
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_17  (.CI(n28734), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n28735));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n24213), .I1(n7716[10]), .I2(GND_net), 
            .I3(n29466), .O(n2996[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3712_2_lut (.I0(GND_net), .I1(n8_adj_3570), .I2(n77), 
            .I3(GND_net), .O(n8013[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3712_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n29466), .I0(n7716[10]), .I1(GND_net), 
            .CO(n29467));
    SB_CARRY add_3712_2 (.CI(GND_net), .I0(n8_adj_3570), .I1(n77), .CO(n29678));
    SB_LUT4 add_3706_7_lut (.I0(GND_net), .I1(n36676), .I2(n490), .I3(n29677), 
            .O(n7980[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3706_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n24213), .I1(n7716[9]), .I2(GND_net), 
            .I3(n29465), .O(n2996[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3721_9 (.CI(n29859), .I0(n8208[6]), .I1(GND_net), .CO(n29860));
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3706_6_lut (.I0(GND_net), .I1(n7988[3]), .I2(n417), .I3(n29676), 
            .O(n7980[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3706_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_8_lut (.I0(GND_net), .I1(n8208[5]), .I2(n542), .I3(n29858), 
            .O(n8193[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n29465), .I0(n7716[9]), .I1(GND_net), 
            .CO(n29466));
    SB_CARRY add_3721_8 (.CI(n29858), .I0(n8208[5]), .I1(n542), .CO(n29859));
    SB_LUT4 add_3721_7_lut (.I0(GND_net), .I1(n8208[4]), .I2(n469), .I3(n29857), 
            .O(n8193[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n24213), .I1(n7716[8]), .I2(GND_net), 
            .I3(n29464), .O(n2996[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3721_7 (.CI(n29857), .I0(n8208[4]), .I1(n469), .CO(n29858));
    SB_CARRY add_3706_6 (.CI(n29676), .I0(n7988[3]), .I1(n417), .CO(n29677));
    SB_LUT4 add_3706_5_lut (.I0(GND_net), .I1(n7988[2]), .I2(n344), .I3(n29675), 
            .O(n7980[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3706_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3706_5 (.CI(n29675), .I0(n7988[2]), .I1(n344), .CO(n29676));
    SB_LUT4 add_3706_4_lut (.I0(GND_net), .I1(n7988[1]), .I2(n271), .I3(n29674), 
            .O(n7980[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3706_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n29464), .I0(n7716[8]), .I1(GND_net), 
            .CO(n29465));
    SB_LUT4 add_3721_6_lut (.I0(GND_net), .I1(n8208[3]), .I2(n396), .I3(n29856), 
            .O(n8193[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3706_4 (.CI(n29674), .I0(n7988[1]), .I1(n271), .CO(n29675));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n28733), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n24213), .I1(n7716[7]), .I2(GND_net), 
            .I3(n29463), .O(n2996[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_16  (.CI(n28733), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n28734));
    SB_CARRY add_636_10 (.CI(n28007), .I0(n2996[8]), .I1(n3021[8]), .CO(n28008));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n28732), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_6 (.CI(n29856), .I0(n8208[3]), .I1(n396), .CO(n29857));
    SB_LUT4 add_3706_3_lut (.I0(GND_net), .I1(n7988[0]), .I2(n198_adj_3589), 
            .I3(n29673), .O(n7980[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3706_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3706_3 (.CI(n29673), .I0(n7988[0]), .I1(n198_adj_3589), 
            .CO(n29674));
    SB_CARRY mult_10_add_1225_10 (.CI(n29463), .I0(n7716[7]), .I1(GND_net), 
            .CO(n29464));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n24213), .I1(n7716[6]), .I2(GND_net), 
            .I3(n29462), .O(n2996[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_9 (.CI(n29462), .I0(n7716[6]), .I1(GND_net), 
            .CO(n29463));
    SB_LUT4 add_3721_5_lut (.I0(GND_net), .I1(n8208[2]), .I2(n323), .I3(n29855), 
            .O(n8193[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_5 (.CI(n29855), .I0(n8208[2]), .I1(n323), .CO(n29856));
    SB_LUT4 add_3721_4_lut (.I0(GND_net), .I1(n8208[1]), .I2(n250), .I3(n29854), 
            .O(n8193[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_15  (.CI(n28732), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n28733));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n28731), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[11]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3706_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n7980[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3706_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n24213), .I1(n7716[5]), .I2(n512_adj_3592), 
            .I3(n29461), .O(n2996[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_8 (.CI(n29461), .I0(n7716[5]), .I1(n512_adj_3592), 
            .CO(n29462));
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_14  (.CI(n28731), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n28732));
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[12]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[13]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n24213), .I1(n7716[4]), .I2(n439_adj_3595), 
            .I3(n29460), .O(n2996[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n28730), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_13  (.CI(n28730), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n28731));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n28729), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_12  (.CI(n28729), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n28730));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n28728), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_4 (.CI(n29854), .I0(n8208[1]), .I1(n250), .CO(n29855));
    SB_CARRY add_3706_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n29673));
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_11  (.CI(n28728), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n28729));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n28727), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_10  (.CI(n28727), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n28728));
    SB_CARRY mult_10_add_1225_7 (.CI(n29460), .I0(n7716[4]), .I1(n439_adj_3595), 
            .CO(n29461));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n28726), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_9  (.CI(n28726), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n28727));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n24213), .I1(n7716[3]), .I2(n366_adj_3596), 
            .I3(n29459), .O(n2996[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3705_8_lut (.I0(GND_net), .I1(n7980[5]), .I2(n560), .I3(n29672), 
            .O(n7971[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3705_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_3891[8]), .I3(n28140), .O(n17_adj_3597)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n28725), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_636_9_lut (.I0(GND_net), .I1(n2996[7]), .I2(n3021[7]), 
            .I3(n28006), .O(duty_23__N_3478[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n29459), .I0(n7716[3]), .I1(n366_adj_3596), 
            .CO(n29460));
    SB_LUT4 add_3721_3_lut (.I0(GND_net), .I1(n8208[0]), .I2(n177), .I3(n29853), 
            .O(n8193[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_8  (.CI(n28725), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n28726));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n28724), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3705_7_lut (.I0(GND_net), .I1(n7980[4]), .I2(n487), .I3(n29671), 
            .O(n7971[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3705_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3705_7 (.CI(n29671), .I0(n7980[4]), .I1(n487), .CO(n29672));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n24213), .I1(n7716[2]), .I2(n293_adj_3599), 
            .I3(n29458), .O(n2996[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_7  (.CI(n28724), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n28725));
    SB_LUT4 add_3705_6_lut (.I0(GND_net), .I1(n7980[3]), .I2(n414), .I3(n29670), 
            .O(n7971[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3705_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n29458), .I0(n7716[2]), .I1(n293_adj_3599), 
            .CO(n29459));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n24213), .I1(n7716[1]), .I2(n220_adj_3600), 
            .I3(n29457), .O(n2996[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3721_3 (.CI(n29853), .I0(n8208[0]), .I1(n177), .CO(n29854));
    SB_CARRY unary_minus_5_add_3_10 (.CI(n28140), .I0(GND_net), .I1(n1_adj_3891[8]), 
            .CO(n28141));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n28723), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3721_2_lut (.I0(GND_net), .I1(n35_adj_3601), .I2(n104_adj_3602), 
            .I3(GND_net), .O(n8193[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3721_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3721_2 (.CI(GND_net), .I0(n35_adj_3601), .I1(n104_adj_3602), 
            .CO(n29853));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_3891[7]), .I3(n28139), .O(n15_adj_3603)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_10_add_1225_4 (.CI(n29457), .I0(n7716[1]), .I1(n220_adj_3600), 
            .CO(n29458));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n28139), .I0(GND_net), .I1(n1_adj_3891[7]), 
            .CO(n28140));
    SB_LUT4 add_3720_15_lut (.I0(GND_net), .I1(n8193[12]), .I2(GND_net), 
            .I3(n29852), .O(n8177[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_6  (.CI(n28723), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n28724));
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_3891[6]), .I3(n28138), .O(n13_adj_3605)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3705_6 (.CI(n29670), .I0(n7980[3]), .I1(n414), .CO(n29671));
    SB_LUT4 add_3720_14_lut (.I0(GND_net), .I1(n8193[11]), .I2(GND_net), 
            .I3(n29851), .O(n8177[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n24213), .I1(n7716[0]), .I2(n147_adj_3607), 
            .I3(n29456), .O(n2996[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_636_9 (.CI(n28006), .I0(n2996[7]), .I1(n3021[7]), .CO(n28007));
    SB_LUT4 add_3705_5_lut (.I0(GND_net), .I1(n7980[2]), .I2(n341), .I3(n29669), 
            .O(n7971[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3705_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3705_5 (.CI(n29669), .I0(n7980[2]), .I1(n341), .CO(n29670));
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_3 (.CI(n29456), .I0(n7716[0]), .I1(n147_adj_3607), 
            .CO(n29457));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n24213), .I1(n5_adj_3608), .I2(n74_adj_3609), 
            .I3(GND_net), .O(n2996[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_3608), .I1(n74_adj_3609), 
            .CO(n29456));
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3705_4_lut (.I0(GND_net), .I1(n7980[1]), .I2(n268), .I3(n29668), 
            .O(n7971[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3705_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[15]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n28722), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n28138), .I0(GND_net), .I1(n1_adj_3891[6]), 
            .CO(n28139));
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_5  (.CI(n28722), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n28723));
    SB_LUT4 add_3690_23_lut (.I0(GND_net), .I1(n7740[20]), .I2(GND_net), 
            .I3(n29455), .O(n7716[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3705_4 (.CI(n29668), .I0(n7980[1]), .I1(n268), .CO(n29669));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n28721), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_4  (.CI(n28721), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n28722));
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n28720), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_22_lut (.I0(GND_net), .I1(n7740[19]), .I2(GND_net), 
            .I3(n29454), .O(n7716[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_14 (.CI(n29851), .I0(n8193[11]), .I1(GND_net), .CO(n29852));
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_3  (.CI(n28720), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n28721));
    SB_CARRY add_3690_22 (.CI(n29454), .I0(n7740[19]), .I1(GND_net), .CO(n29455));
    SB_LUT4 add_3690_21_lut (.I0(GND_net), .I1(n7740[18]), .I2(GND_net), 
            .I3(n29453), .O(n7716[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3705_3_lut (.I0(GND_net), .I1(n7980[0]), .I2(n195_adj_3610), 
            .I3(n29667), .O(n7971[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3705_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_21 (.CI(n29453), .I0(n7740[18]), .I1(GND_net), .CO(n29454));
    SB_LUT4 add_3690_20_lut (.I0(GND_net), .I1(n7740[17]), .I2(GND_net), 
            .I3(n29452), .O(n7716[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_20 (.CI(n29452), .I0(n7740[17]), .I1(GND_net), .CO(n29453));
    SB_CARRY add_3705_3 (.CI(n29667), .I0(n7980[0]), .I1(n195_adj_3610), 
            .CO(n29668));
    SB_LUT4 add_3720_13_lut (.I0(GND_net), .I1(n8193[10]), .I2(GND_net), 
            .I3(n29850), .O(n8177[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_19_lut (.I0(GND_net), .I1(n7740[16]), .I2(GND_net), 
            .I3(n29451), .O(n7716[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_19 (.CI(n29451), .I0(n7740[16]), .I1(GND_net), .CO(n29452));
    SB_LUT4 add_3690_18_lut (.I0(GND_net), .I1(n7740[15]), .I2(GND_net), 
            .I3(n29450), .O(n7716[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1179_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1179_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1179_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n28720));
    SB_CARRY add_3690_18 (.CI(n29450), .I0(n7740[15]), .I1(GND_net), .CO(n29451));
    SB_CARRY add_3720_13 (.CI(n29850), .I0(n8193[10]), .I1(GND_net), .CO(n29851));
    SB_LUT4 add_3690_17_lut (.I0(GND_net), .I1(n7740[14]), .I2(GND_net), 
            .I3(n29449), .O(n7716[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_17 (.CI(n29449), .I0(n7740[14]), .I1(GND_net), .CO(n29450));
    SB_LUT4 add_3705_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_3612), 
            .I3(GND_net), .O(n7971[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3705_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3705_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_3612), .CO(n29667));
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3704_9_lut (.I0(GND_net), .I1(n7971[6]), .I2(GND_net), 
            .I3(n29666), .O(n7961[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_12_lut (.I0(GND_net), .I1(n8193[9]), .I2(GND_net), 
            .I3(n29849), .O(n8177[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3704_8_lut (.I0(GND_net), .I1(n7971[5]), .I2(n557), .I3(n29665), 
            .O(n7961[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_16_lut (.I0(GND_net), .I1(n7740[13]), .I2(GND_net), 
            .I3(n29448), .O(n7716[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_16 (.CI(n29448), .I0(n7740[13]), .I1(GND_net), .CO(n29449));
    SB_LUT4 add_3690_15_lut (.I0(GND_net), .I1(n7740[12]), .I2(GND_net), 
            .I3(n29447), .O(n7716[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3704_8 (.CI(n29665), .I0(n7971[5]), .I1(n557), .CO(n29666));
    SB_LUT4 add_3704_7_lut (.I0(GND_net), .I1(n7971[4]), .I2(n484), .I3(n29664), 
            .O(n7961[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_15 (.CI(n29447), .I0(n7740[12]), .I1(GND_net), .CO(n29448));
    SB_LUT4 add_3690_14_lut (.I0(GND_net), .I1(n7740[11]), .I2(GND_net), 
            .I3(n29446), .O(n7716[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_14 (.CI(n29446), .I0(n7740[11]), .I1(GND_net), .CO(n29447));
    SB_CARRY add_3720_12 (.CI(n29849), .I0(n8193[9]), .I1(GND_net), .CO(n29850));
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3690_13_lut (.I0(GND_net), .I1(n7740[10]), .I2(GND_net), 
            .I3(n29445), .O(n7716[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_11_lut (.I0(GND_net), .I1(n8193[8]), .I2(GND_net), 
            .I3(n29848), .O(n8177[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3704_7 (.CI(n29664), .I0(n7971[4]), .I1(n484), .CO(n29665));
    SB_LUT4 add_636_8_lut (.I0(GND_net), .I1(n2996[6]), .I2(n3021[6]), 
            .I3(n28005), .O(duty_23__N_3478[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_11 (.CI(n29848), .I0(n8193[8]), .I1(GND_net), .CO(n29849));
    SB_CARRY add_3690_13 (.CI(n29445), .I0(n7740[10]), .I1(GND_net), .CO(n29446));
    SB_LUT4 add_3690_12_lut (.I0(GND_net), .I1(n7740[9]), .I2(GND_net), 
            .I3(n29444), .O(n7716[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_8 (.CI(n28005), .I0(n2996[6]), .I1(n3021[6]), .CO(n28006));
    SB_LUT4 add_3704_6_lut (.I0(GND_net), .I1(n7971[3]), .I2(n411), .I3(n29663), 
            .O(n7961[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_3891[5]), .I3(n28137), .O(n11_adj_3613)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3720_10_lut (.I0(GND_net), .I1(n8193[7]), .I2(GND_net), 
            .I3(n29847), .O(n8177[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_12 (.CI(n29444), .I0(n7740[9]), .I1(GND_net), .CO(n29445));
    SB_LUT4 add_3690_11_lut (.I0(GND_net), .I1(n7740[8]), .I2(GND_net), 
            .I3(n29443), .O(n7716[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_10 (.CI(n29847), .I0(n8193[7]), .I1(GND_net), .CO(n29848));
    SB_LUT4 add_636_7_lut (.I0(GND_net), .I1(n2996[5]), .I2(n3021[5]), 
            .I3(n28004), .O(duty_23__N_3478[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n28137), .I0(GND_net), .I1(n1_adj_3891[5]), 
            .CO(n28138));
    SB_CARRY add_636_7 (.CI(n28004), .I0(n2996[5]), .I1(n3021[5]), .CO(n28005));
    SB_LUT4 add_3720_9_lut (.I0(GND_net), .I1(n8193[6]), .I2(GND_net), 
            .I3(n29846), .O(n8177[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3704_6 (.CI(n29663), .I0(n7971[3]), .I1(n411), .CO(n29664));
    SB_CARRY add_3720_9 (.CI(n29846), .I0(n8193[6]), .I1(GND_net), .CO(n29847));
    SB_LUT4 add_3704_5_lut (.I0(GND_net), .I1(n7971[2]), .I2(n338), .I3(n29662), 
            .O(n7961[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_8_lut (.I0(GND_net), .I1(n8193[5]), .I2(n539), .I3(n29845), 
            .O(n8177[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3704_5 (.CI(n29662), .I0(n7971[2]), .I1(n338), .CO(n29663));
    SB_CARRY add_3690_11 (.CI(n29443), .I0(n7740[8]), .I1(GND_net), .CO(n29444));
    SB_LUT4 add_3690_10_lut (.I0(GND_net), .I1(n7740[7]), .I2(GND_net), 
            .I3(n29442), .O(n7716[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_10 (.CI(n29442), .I0(n7740[7]), .I1(GND_net), .CO(n29443));
    SB_LUT4 add_3704_4_lut (.I0(GND_net), .I1(n7971[1]), .I2(n265), .I3(n29661), 
            .O(n7961[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_9_lut (.I0(GND_net), .I1(n7740[6]), .I2(GND_net), 
            .I3(n29441), .O(n7716[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_9 (.CI(n29441), .I0(n7740[6]), .I1(GND_net), .CO(n29442));
    SB_LUT4 add_3690_8_lut (.I0(GND_net), .I1(n7740[5]), .I2(n515_adj_3615), 
            .I3(n29440), .O(n7716[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_3891[4]), .I3(n28136), .O(n9_adj_3616)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[12]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3690_8 (.CI(n29440), .I0(n7740[5]), .I1(n515_adj_3615), 
            .CO(n29441));
    SB_LUT4 add_636_6_lut (.I0(GND_net), .I1(n2996[4]), .I2(n3021[4]), 
            .I3(n28003), .O(duty_23__N_3478[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_8 (.CI(n29845), .I0(n8193[5]), .I1(n539), .CO(n29846));
    SB_CARRY add_3704_4 (.CI(n29661), .I0(n7971[1]), .I1(n265), .CO(n29662));
    SB_LUT4 add_3690_7_lut (.I0(GND_net), .I1(n7740[4]), .I2(n442_adj_3618), 
            .I3(n29439), .O(n7716[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_7 (.CI(n29439), .I0(n7740[4]), .I1(n442_adj_3618), 
            .CO(n29440));
    SB_LUT4 add_3720_7_lut (.I0(GND_net), .I1(n8193[4]), .I2(n466), .I3(n29844), 
            .O(n8177[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_6_lut (.I0(GND_net), .I1(n7740[3]), .I2(n369_adj_3619), 
            .I3(n29438), .O(n7716[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_6 (.CI(n29438), .I0(n7740[3]), .I1(n369_adj_3619), 
            .CO(n29439));
    SB_CARRY add_636_6 (.CI(n28003), .I0(n2996[4]), .I1(n3021[4]), .CO(n28004));
    SB_LUT4 add_3690_5_lut (.I0(GND_net), .I1(n7740[2]), .I2(n296_adj_3620), 
            .I3(n29437), .O(n7716[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_5 (.CI(n29437), .I0(n7740[2]), .I1(n296_adj_3620), 
            .CO(n29438));
    SB_LUT4 add_3704_3_lut (.I0(GND_net), .I1(n7971[0]), .I2(n192_adj_3621), 
            .I3(n29660), .O(n7961[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n28136), .I0(GND_net), .I1(n1_adj_3891[4]), 
            .CO(n28137));
    SB_CARRY add_3720_7 (.CI(n29844), .I0(n8193[4]), .I1(n466), .CO(n29845));
    SB_CARRY add_3704_3 (.CI(n29660), .I0(n7971[0]), .I1(n192_adj_3621), 
            .CO(n29661));
    SB_LUT4 add_3720_6_lut (.I0(GND_net), .I1(n8193[3]), .I2(n393), .I3(n29843), 
            .O(n8177[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3704_2_lut (.I0(GND_net), .I1(n50), .I2(n119_adj_3622), 
            .I3(GND_net), .O(n7961[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_4_lut (.I0(GND_net), .I1(n7740[1]), .I2(n223_adj_3623), 
            .I3(n29436), .O(n7716[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_4 (.CI(n29436), .I0(n7740[1]), .I1(n223_adj_3623), 
            .CO(n29437));
    SB_LUT4 i23021_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n7995[0]));   // verilog/motorControl.v(42[17:23])
    defparam i23021_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_3704_2 (.CI(GND_net), .I0(n50), .I1(n119_adj_3622), .CO(n29660));
    SB_LUT4 add_3703_10_lut (.I0(GND_net), .I1(n7961[7]), .I2(GND_net), 
            .I3(n29659), .O(n7950[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_3_lut (.I0(GND_net), .I1(n7740[0]), .I2(n150_adj_3624), 
            .I3(n29435), .O(n7716[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3690_3 (.CI(n29435), .I0(n7740[0]), .I1(n150_adj_3624), 
            .CO(n29436));
    SB_LUT4 add_3703_9_lut (.I0(GND_net), .I1(n7961[6]), .I2(GND_net), 
            .I3(n29658), .O(n7950[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_3891[3]), .I3(n28135), .O(n7_adj_3625)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3703_9 (.CI(n29658), .I0(n7961[6]), .I1(GND_net), .CO(n29659));
    SB_CARRY unary_minus_5_add_3_5 (.CI(n28135), .I0(GND_net), .I1(n1_adj_3891[3]), 
            .CO(n28136));
    SB_CARRY add_3720_6 (.CI(n29843), .I0(n8193[3]), .I1(n393), .CO(n29844));
    SB_LUT4 add_3703_8_lut (.I0(GND_net), .I1(n7961[5]), .I2(n554), .I3(n29657), 
            .O(n7950[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3690_2_lut (.I0(GND_net), .I1(n8_adj_3626), .I2(n77_adj_3627), 
            .I3(GND_net), .O(n7716[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3690_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_5_lut (.I0(GND_net), .I1(n8193[2]), .I2(n320), .I3(n29842), 
            .O(n8177[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3703_8 (.CI(n29657), .I0(n7961[5]), .I1(n554), .CO(n29658));
    SB_LUT4 add_3703_7_lut (.I0(GND_net), .I1(n7961[4]), .I2(n481), .I3(n29656), 
            .O(n7950[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3703_7 (.CI(n29656), .I0(n7961[4]), .I1(n481), .CO(n29657));
    SB_CARRY add_3690_2 (.CI(GND_net), .I0(n8_adj_3626), .I1(n77_adj_3627), 
            .CO(n29435));
    SB_CARRY add_3720_5 (.CI(n29842), .I0(n8193[2]), .I1(n320), .CO(n29843));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_3891[2]), .I3(n28134), .O(n5_adj_3628)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3720_4_lut (.I0(GND_net), .I1(n8193[1]), .I2(n247), .I3(n29841), 
            .O(n8177[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_4 (.CI(n29841), .I0(n8193[1]), .I1(n247), .CO(n29842));
    SB_LUT4 add_3720_3_lut (.I0(GND_net), .I1(n8193[0]), .I2(n174), .I3(n29840), 
            .O(n8177[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3703_6_lut (.I0(GND_net), .I1(n7961[3]), .I2(n408), .I3(n29655), 
            .O(n7950[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_3 (.CI(n29840), .I0(n8193[0]), .I1(n174), .CO(n29841));
    SB_CARRY add_3703_6 (.CI(n29655), .I0(n7961[3]), .I1(n408), .CO(n29656));
    SB_LUT4 add_3703_5_lut (.I0(GND_net), .I1(n7961[2]), .I2(n335), .I3(n29654), 
            .O(n7950[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3720_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8177[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3720_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3720_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n29840));
    SB_CARRY add_3703_5 (.CI(n29654), .I0(n7961[2]), .I1(n335), .CO(n29655));
    SB_LUT4 add_3703_4_lut (.I0(GND_net), .I1(n7961[1]), .I2(n262), .I3(n29653), 
            .O(n7950[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3703_4 (.CI(n29653), .I0(n7961[1]), .I1(n262), .CO(n29654));
    SB_LUT4 add_3703_3_lut (.I0(GND_net), .I1(n7961[0]), .I2(n189_adj_3630), 
            .I3(n29652), .O(n7950[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3703_3 (.CI(n29652), .I0(n7961[0]), .I1(n189_adj_3630), 
            .CO(n29653));
    SB_LUT4 add_3719_16_lut (.I0(GND_net), .I1(n8177[13]), .I2(GND_net), 
            .I3(n29839), .O(n8160[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_15_lut (.I0(GND_net), .I1(n8177[12]), .I2(GND_net), 
            .I3(n29838), .O(n8160[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3703_2_lut (.I0(GND_net), .I1(n47), .I2(n116_adj_3631), 
            .I3(GND_net), .O(n7950[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3703_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3703_2 (.CI(GND_net), .I0(n47), .I1(n116_adj_3631), .CO(n29652));
    SB_LUT4 add_3702_11_lut (.I0(GND_net), .I1(n7950[8]), .I2(GND_net), 
            .I3(n29651), .O(n7938[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3702_10_lut (.I0(GND_net), .I1(n7950[7]), .I2(GND_net), 
            .I3(n29650), .O(n7938[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[14]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[15]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3719_15 (.CI(n29838), .I0(n8177[12]), .I1(GND_net), .CO(n29839));
    SB_CARRY add_3702_10 (.CI(n29650), .I0(n7950[7]), .I1(GND_net), .CO(n29651));
    SB_LUT4 mux_634_i13_3_lut (.I0(n155[12]), .I1(PWMLimit[12]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i13_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3702_9_lut (.I0(GND_net), .I1(n7950[6]), .I2(GND_net), 
            .I3(n29649), .O(n7938[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_636_5_lut (.I0(GND_net), .I1(n2996[3]), .I2(n3021[3]), 
            .I3(n28002), .O(duty_23__N_3478[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_14_lut (.I0(GND_net), .I1(n8177[11]), .I2(GND_net), 
            .I3(n29837), .O(n8160[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3702_9 (.CI(n29649), .I0(n7950[6]), .I1(GND_net), .CO(n29650));
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3702_8_lut (.I0(GND_net), .I1(n7950[5]), .I2(n551), .I3(n29648), 
            .O(n7938[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3702_8 (.CI(n29648), .I0(n7950[5]), .I1(n551), .CO(n29649));
    SB_LUT4 add_3702_7_lut (.I0(GND_net), .I1(n7950[4]), .I2(n478), .I3(n29647), 
            .O(n7938[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_5 (.CI(n28002), .I0(n2996[3]), .I1(n3021[3]), .CO(n28003));
    SB_CARRY add_3719_14 (.CI(n29837), .I0(n8177[11]), .I1(GND_net), .CO(n29838));
    SB_LUT4 add_3719_13_lut (.I0(GND_net), .I1(n8177[10]), .I2(GND_net), 
            .I3(n29836), .O(n8160[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3719_13 (.CI(n29836), .I0(n8177[10]), .I1(GND_net), .CO(n29837));
    SB_CARRY add_3702_7 (.CI(n29647), .I0(n7950[4]), .I1(n478), .CO(n29648));
    SB_LUT4 add_3702_6_lut (.I0(GND_net), .I1(n7950[3]), .I2(n405), .I3(n29646), 
            .O(n7938[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3719_12_lut (.I0(GND_net), .I1(n8177[9]), .I2(GND_net), 
            .I3(n29835), .O(n8160[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3702_6 (.CI(n29646), .I0(n7950[3]), .I1(n405), .CO(n29647));
    SB_CARRY add_3719_12 (.CI(n29835), .I0(n8177[9]), .I1(GND_net), .CO(n29836));
    SB_LUT4 add_3702_5_lut (.I0(GND_net), .I1(n7950[2]), .I2(n332), .I3(n29645), 
            .O(n7938[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n28134), .I0(GND_net), .I1(n1_adj_3891[2]), 
            .CO(n28135));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_3891[1]), .I3(n28133), .O(n3_adj_3634)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n28133), .I0(GND_net), .I1(n1_adj_3891[1]), 
            .CO(n28134));
    SB_CARRY add_3702_5 (.CI(n29645), .I0(n7950[2]), .I1(n332), .CO(n29646));
    SB_LUT4 add_3702_4_lut (.I0(GND_net), .I1(n7950[1]), .I2(n259), .I3(n29644), 
            .O(n7938[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[13]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3702_4 (.CI(n29644), .I0(n7950[1]), .I1(n259), .CO(n29645));
    SB_LUT4 add_3702_3_lut (.I0(GND_net), .I1(n7950[0]), .I2(n186_adj_3635), 
            .I3(n29643), .O(n7938[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3891[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3454 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3478[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_3891[0]), 
            .CO(n28133));
    SB_LUT4 add_3719_11_lut (.I0(GND_net), .I1(n8177[8]), .I2(GND_net), 
            .I3(n29834), .O(n8160[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3575));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3702_3 (.CI(n29643), .I0(n7950[0]), .I1(n186_adj_3635), 
            .CO(n29644));
    SB_LUT4 add_3702_2_lut (.I0(GND_net), .I1(n44_adj_3637), .I2(n113_adj_3638), 
            .I3(GND_net), .O(n7938[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3702_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_11 (.CI(n29834), .I0(n8177[8]), .I1(GND_net), .CO(n29835));
    SB_LUT4 add_3719_10_lut (.I0(GND_net), .I1(n8177[7]), .I2(GND_net), 
            .I3(n29833), .O(n8160[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_10 (.CI(n29833), .I0(n8177[7]), .I1(GND_net), .CO(n29834));
    SB_LUT4 add_3719_9_lut (.I0(GND_net), .I1(n8177[6]), .I2(GND_net), 
            .I3(n29832), .O(n8160[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_9 (.CI(n29832), .I0(n8177[6]), .I1(GND_net), .CO(n29833));
    SB_LUT4 add_3719_8_lut (.I0(GND_net), .I1(n8177[5]), .I2(n536_adj_3639), 
            .I3(n29831), .O(n8160[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_8 (.CI(n29831), .I0(n8177[5]), .I1(n536_adj_3639), 
            .CO(n29832));
    SB_LUT4 add_3719_7_lut (.I0(GND_net), .I1(n8177[4]), .I2(n463_adj_3640), 
            .I3(n29830), .O(n8160[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3702_2 (.CI(GND_net), .I0(n44_adj_3637), .I1(n113_adj_3638), 
            .CO(n29643));
    SB_LUT4 add_3701_12_lut (.I0(GND_net), .I1(n7938[9]), .I2(GND_net), 
            .I3(n29642), .O(n7925[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3701_11_lut (.I0(GND_net), .I1(n7938[8]), .I2(GND_net), 
            .I3(n29641), .O(n7925[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_7 (.CI(n29830), .I0(n8177[4]), .I1(n463_adj_3640), 
            .CO(n29831));
    SB_CARRY add_3701_11 (.CI(n29641), .I0(n7938[8]), .I1(GND_net), .CO(n29642));
    SB_LUT4 add_3719_6_lut (.I0(GND_net), .I1(n8177[3]), .I2(n390_adj_3641), 
            .I3(n29829), .O(n8160[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3701_10_lut (.I0(GND_net), .I1(n7938[7]), .I2(GND_net), 
            .I3(n29640), .O(n7925[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3478[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3719_6 (.CI(n29829), .I0(n8177[3]), .I1(n390_adj_3641), 
            .CO(n29830));
    SB_CARRY add_3701_10 (.CI(n29640), .I0(n7938[7]), .I1(GND_net), .CO(n29641));
    SB_LUT4 add_3701_9_lut (.I0(GND_net), .I1(n7938[6]), .I2(GND_net), 
            .I3(n29639), .O(n7925[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3701_9 (.CI(n29639), .I0(n7938[6]), .I1(GND_net), .CO(n29640));
    SB_LUT4 add_3719_5_lut (.I0(GND_net), .I1(n8177[2]), .I2(n317_adj_3642), 
            .I3(n29828), .O(n8160[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3701_8_lut (.I0(GND_net), .I1(n7938[5]), .I2(n548_adj_3643), 
            .I3(n29638), .O(n7925[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_5 (.CI(n29828), .I0(n8177[2]), .I1(n317_adj_3642), 
            .CO(n29829));
    SB_LUT4 add_3719_4_lut (.I0(GND_net), .I1(n8177[1]), .I2(n244_adj_3644), 
            .I3(n29827), .O(n8160[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3478[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3478[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3478[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3719_4 (.CI(n29827), .I0(n8177[1]), .I1(n244_adj_3644), 
            .CO(n29828));
    SB_LUT4 add_3719_3_lut (.I0(GND_net), .I1(n8177[0]), .I2(n171_adj_3645), 
            .I3(n29826), .O(n8160[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3701_8 (.CI(n29638), .I0(n7938[5]), .I1(n548_adj_3643), 
            .CO(n29639));
    SB_CARRY add_3719_3 (.CI(n29826), .I0(n8177[0]), .I1(n171_adj_3645), 
            .CO(n29827));
    SB_LUT4 add_3719_2_lut (.I0(GND_net), .I1(n29_adj_3646), .I2(n98_adj_3647), 
            .I3(GND_net), .O(n8160[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3719_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3719_2 (.CI(GND_net), .I0(n29_adj_3646), .I1(n98_adj_3647), 
            .CO(n29826));
    SB_LUT4 add_3718_17_lut (.I0(GND_net), .I1(n8160[14]), .I2(GND_net), 
            .I3(n29825), .O(n8142[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3701_7_lut (.I0(GND_net), .I1(n7938[4]), .I2(n475_adj_3648), 
            .I3(n29637), .O(n7925[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3478[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3718_16_lut (.I0(GND_net), .I1(n8160[13]), .I2(GND_net), 
            .I3(n29824), .O(n8142[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3478[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3649));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3478[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3478[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_636_4_lut (.I0(GND_net), .I1(n2996[2]), .I2(n3021[2]), 
            .I3(n28001), .O(duty_23__N_3478[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3701_7 (.CI(n29637), .I0(n7938[4]), .I1(n475_adj_3648), 
            .CO(n29638));
    SB_CARRY add_3718_16 (.CI(n29824), .I0(n8160[13]), .I1(GND_net), .CO(n29825));
    SB_LUT4 add_3701_6_lut (.I0(GND_net), .I1(n7938[3]), .I2(n402_adj_3650), 
            .I3(n29636), .O(n7925[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3651));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3478[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3701_6 (.CI(n29636), .I0(n7938[3]), .I1(n402_adj_3650), 
            .CO(n29637));
    SB_LUT4 add_3718_15_lut (.I0(GND_net), .I1(n8160[12]), .I2(GND_net), 
            .I3(n29823), .O(n8142[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3701_5_lut (.I0(GND_net), .I1(n7938[2]), .I2(n329_adj_3652), 
            .I3(n29635), .O(n7925[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_15 (.CI(n29823), .I0(n8160[12]), .I1(GND_net), .CO(n29824));
    SB_CARRY add_3701_5 (.CI(n29635), .I0(n7938[2]), .I1(n329_adj_3652), 
            .CO(n29636));
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3478[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3701_4_lut (.I0(GND_net), .I1(n7938[1]), .I2(n256_adj_3653), 
            .I3(n29634), .O(n7925[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3701_4 (.CI(n29634), .I0(n7938[1]), .I1(n256_adj_3653), 
            .CO(n29635));
    SB_LUT4 add_3701_3_lut (.I0(GND_net), .I1(n7938[0]), .I2(n183_adj_3654), 
            .I3(n29633), .O(n7925[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_14_lut (.I0(GND_net), .I1(n8160[11]), .I2(GND_net), 
            .I3(n29822), .O(n8142[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3701_3 (.CI(n29633), .I0(n7938[0]), .I1(n183_adj_3654), 
            .CO(n29634));
    SB_LUT4 add_3701_2_lut (.I0(GND_net), .I1(n41_adj_3655), .I2(n110_adj_3656), 
            .I3(GND_net), .O(n7925[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3701_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3701_2 (.CI(GND_net), .I0(n41_adj_3655), .I1(n110_adj_3656), 
            .CO(n29633));
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3478[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3478[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3700_13_lut (.I0(GND_net), .I1(n7925[10]), .I2(GND_net), 
            .I3(n29632), .O(n7911[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3478[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3700_12_lut (.I0(GND_net), .I1(n7925[9]), .I2(GND_net), 
            .I3(n29631), .O(n7911[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3700_12 (.CI(n29631), .I0(n7925[9]), .I1(GND_net), .CO(n29632));
    SB_CARRY add_3718_14 (.CI(n29822), .I0(n8160[11]), .I1(GND_net), .CO(n29823));
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3478[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3718_13_lut (.I0(GND_net), .I1(n8160[10]), .I2(GND_net), 
            .I3(n29821), .O(n8142[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_13 (.CI(n29821), .I0(n8160[10]), .I1(GND_net), .CO(n29822));
    SB_LUT4 add_3700_11_lut (.I0(GND_net), .I1(n7925[8]), .I2(GND_net), 
            .I3(n29630), .O(n7911[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3478[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3478[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3700_11 (.CI(n29630), .I0(n7925[8]), .I1(GND_net), .CO(n29631));
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3478[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3478[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3478[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3478[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3478[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3657));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3718_12_lut (.I0(GND_net), .I1(n8160[9]), .I2(GND_net), 
            .I3(n29820), .O(n8142[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_12 (.CI(n29820), .I0(n8160[9]), .I1(GND_net), .CO(n29821));
    SB_LUT4 add_3700_10_lut (.I0(GND_net), .I1(n7925[7]), .I2(GND_net), 
            .I3(n29629), .O(n7911[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3700_10 (.CI(n29629), .I0(n7925[7]), .I1(GND_net), .CO(n29630));
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[16]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3700_9_lut (.I0(GND_net), .I1(n7925[6]), .I2(GND_net), 
            .I3(n29628), .O(n7911[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_11_lut (.I0(GND_net), .I1(n8160[8]), .I2(GND_net), 
            .I3(n29819), .O(n8142[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_11 (.CI(n29819), .I0(n8160[8]), .I1(GND_net), .CO(n29820));
    SB_CARRY add_3700_9 (.CI(n29628), .I0(n7925[6]), .I1(GND_net), .CO(n29629));
    SB_LUT4 add_3700_8_lut (.I0(GND_net), .I1(n7925[5]), .I2(n545_adj_3659), 
            .I3(n29627), .O(n7911[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_10_lut (.I0(GND_net), .I1(n8160[7]), .I2(GND_net), 
            .I3(n29818), .O(n8142[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3700_8 (.CI(n29627), .I0(n7925[5]), .I1(n545_adj_3659), 
            .CO(n29628));
    SB_LUT4 add_3700_7_lut (.I0(GND_net), .I1(n7925[4]), .I2(n472_adj_3660), 
            .I3(n29626), .O(n7911[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_4 (.CI(n28001), .I0(n2996[2]), .I1(n3021[2]), .CO(n28002));
    SB_CARRY add_3700_7 (.CI(n29626), .I0(n7925[4]), .I1(n472_adj_3660), 
            .CO(n29627));
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3661));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3700_6_lut (.I0(GND_net), .I1(n7925[3]), .I2(n399_adj_3662), 
            .I3(n29625), .O(n7911[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3700_6 (.CI(n29625), .I0(n7925[3]), .I1(n399_adj_3662), 
            .CO(n29626));
    SB_LUT4 add_3700_5_lut (.I0(GND_net), .I1(n7925[2]), .I2(n326_adj_3663), 
            .I3(n29624), .O(n7911[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_10 (.CI(n29818), .I0(n8160[7]), .I1(GND_net), .CO(n29819));
    SB_LUT4 add_636_3_lut (.I0(GND_net), .I1(n2996[1]), .I2(n3021[1]), 
            .I3(n28000), .O(duty_23__N_3478[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3700_5 (.CI(n29624), .I0(n7925[2]), .I1(n326_adj_3663), 
            .CO(n29625));
    SB_LUT4 add_3718_9_lut (.I0(GND_net), .I1(n8160[6]), .I2(GND_net), 
            .I3(n29817), .O(n8142[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_9 (.CI(n29817), .I0(n8160[6]), .I1(GND_net), .CO(n29818));
    SB_LUT4 add_3718_8_lut (.I0(GND_net), .I1(n8160[5]), .I2(n533), .I3(n29816), 
            .O(n8142[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_8 (.CI(n29816), .I0(n8160[5]), .I1(n533), .CO(n29817));
    SB_LUT4 add_3700_4_lut (.I0(GND_net), .I1(n7925[1]), .I2(n253_adj_3664), 
            .I3(n29623), .O(n7911[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3718_7_lut (.I0(GND_net), .I1(n8160[4]), .I2(n460), .I3(n29815), 
            .O(n8142[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_7 (.CI(n29815), .I0(n8160[4]), .I1(n460), .CO(n29816));
    SB_CARRY add_3700_4 (.CI(n29623), .I0(n7925[1]), .I1(n253_adj_3664), 
            .CO(n29624));
    SB_CARRY add_636_3 (.CI(n28000), .I0(n2996[1]), .I1(n3021[1]), .CO(n28001));
    SB_LUT4 add_3700_3_lut (.I0(GND_net), .I1(n7925[0]), .I2(n180_adj_3665), 
            .I3(n29622), .O(n7911[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3700_3 (.CI(n29622), .I0(n7925[0]), .I1(n180_adj_3665), 
            .CO(n29623));
    SB_LUT4 add_3700_2_lut (.I0(GND_net), .I1(n38_adj_3666), .I2(n107_adj_3667), 
            .I3(GND_net), .O(n7911[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3700_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3700_2 (.CI(GND_net), .I0(n38_adj_3666), .I1(n107_adj_3667), 
            .CO(n29622));
    SB_LUT4 add_3699_14_lut (.I0(GND_net), .I1(n7911[11]), .I2(GND_net), 
            .I3(n29621), .O(n7896[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3668));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3669));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_636_2_lut (.I0(GND_net), .I1(n2996[0]), .I2(n3021[0]), 
            .I3(GND_net), .O(duty_23__N_3478[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3670));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3671));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3718_6_lut (.I0(GND_net), .I1(n8160[3]), .I2(n387), .I3(n29814), 
            .O(n8142[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_6 (.CI(n29814), .I0(n8160[3]), .I1(n387), .CO(n29815));
    SB_LUT4 add_3718_5_lut (.I0(GND_net), .I1(n8160[2]), .I2(n314), .I3(n29813), 
            .O(n8142[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_2 (.CI(GND_net), .I0(n2996[0]), .I1(n3021[0]), .CO(n28000));
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3672));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3718_5 (.CI(n29813), .I0(n8160[2]), .I1(n314), .CO(n29814));
    SB_LUT4 add_3718_4_lut (.I0(GND_net), .I1(n8160[1]), .I2(n241), .I3(n29812), 
            .O(n8142[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3673));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3674));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3675));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3718_4 (.CI(n29812), .I0(n8160[1]), .I1(n241), .CO(n29813));
    SB_LUT4 add_3718_3_lut (.I0(GND_net), .I1(n8160[0]), .I2(n168), .I3(n29811), 
            .O(n8142[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3676));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3677));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3699_13_lut (.I0(GND_net), .I1(n7911[10]), .I2(GND_net), 
            .I3(n29620), .O(n7896[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_3 (.CI(n29811), .I0(n8160[0]), .I1(n168), .CO(n29812));
    SB_CARRY add_3699_13 (.CI(n29620), .I0(n7911[10]), .I1(GND_net), .CO(n29621));
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3678));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3718_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n8142[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3718_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3699_12_lut (.I0(GND_net), .I1(n7911[9]), .I2(GND_net), 
            .I3(n29619), .O(n7896[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3718_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n29811));
    SB_LUT4 add_3717_18_lut (.I0(GND_net), .I1(n8142[15]), .I2(GND_net), 
            .I3(n29810), .O(n8123[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_17_lut (.I0(GND_net), .I1(n8142[14]), .I2(GND_net), 
            .I3(n29809), .O(n8123[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_17 (.CI(n29809), .I0(n8142[14]), .I1(GND_net), .CO(n29810));
    SB_CARRY add_3699_12 (.CI(n29619), .I0(n7911[9]), .I1(GND_net), .CO(n29620));
    SB_LUT4 add_3717_16_lut (.I0(GND_net), .I1(n8142[13]), .I2(GND_net), 
            .I3(n29808), .O(n8123[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_16 (.CI(n29808), .I0(n8142[13]), .I1(GND_net), .CO(n29809));
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3679));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[17]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3681));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3717_15_lut (.I0(GND_net), .I1(n8142[12]), .I2(GND_net), 
            .I3(n29807), .O(n8123[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3682));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3699_11_lut (.I0(GND_net), .I1(n7911[8]), .I2(GND_net), 
            .I3(n29618), .O(n7896[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_15 (.CI(n29807), .I0(n8142[12]), .I1(GND_net), .CO(n29808));
    SB_LUT4 add_3717_14_lut (.I0(GND_net), .I1(n8142[11]), .I2(GND_net), 
            .I3(n29806), .O(n8123[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_14 (.CI(n29806), .I0(n8142[11]), .I1(GND_net), .CO(n29807));
    SB_CARRY add_3699_11 (.CI(n29618), .I0(n7911[8]), .I1(GND_net), .CO(n29619));
    SB_LUT4 add_3717_13_lut (.I0(GND_net), .I1(n8142[10]), .I2(GND_net), 
            .I3(n29805), .O(n8123[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_13 (.CI(n29805), .I0(n8142[10]), .I1(GND_net), .CO(n29806));
    SB_LUT4 add_3717_12_lut (.I0(GND_net), .I1(n8142[9]), .I2(GND_net), 
            .I3(n29804), .O(n8123[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3478[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3717_12 (.CI(n29804), .I0(n8142[9]), .I1(GND_net), .CO(n29805));
    SB_LUT4 add_3717_11_lut (.I0(GND_net), .I1(n8142[8]), .I2(GND_net), 
            .I3(n29803), .O(n8123[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3699_10_lut (.I0(GND_net), .I1(n7911[7]), .I2(GND_net), 
            .I3(n29617), .O(n7896[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_11 (.CI(n29803), .I0(n8142[8]), .I1(GND_net), .CO(n29804));
    SB_LUT4 add_3717_10_lut (.I0(GND_net), .I1(n8142[7]), .I2(GND_net), 
            .I3(n29802), .O(n8123[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_10 (.CI(n29802), .I0(n8142[7]), .I1(GND_net), .CO(n29803));
    SB_CARRY add_3699_10 (.CI(n29617), .I0(n7911[7]), .I1(GND_net), .CO(n29618));
    SB_LUT4 add_3717_9_lut (.I0(GND_net), .I1(n8142[6]), .I2(GND_net), 
            .I3(n29801), .O(n8123[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_9 (.CI(n29801), .I0(n8142[6]), .I1(GND_net), .CO(n29802));
    SB_LUT4 add_3699_9_lut (.I0(GND_net), .I1(n7911[6]), .I2(GND_net), 
            .I3(n29616), .O(n7896[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3717_8_lut (.I0(GND_net), .I1(n8142[5]), .I2(n530), .I3(n29800), 
            .O(n8123[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_8 (.CI(n29800), .I0(n8142[5]), .I1(n530), .CO(n29801));
    SB_LUT4 mux_634_i15_3_lut (.I0(n155[14]), .I1(PWMLimit[14]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i15_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3717_7_lut (.I0(GND_net), .I1(n8142[4]), .I2(n457), .I3(n29799), 
            .O(n8123[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_7 (.CI(n29799), .I0(n8142[4]), .I1(n457), .CO(n29800));
    SB_CARRY add_3699_9 (.CI(n29616), .I0(n7911[6]), .I1(GND_net), .CO(n29617));
    SB_LUT4 add_3717_6_lut (.I0(GND_net), .I1(n8142[3]), .I2(n384), .I3(n29798), 
            .O(n8123[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_6 (.CI(n29798), .I0(n8142[3]), .I1(n384), .CO(n29799));
    SB_LUT4 add_3717_5_lut (.I0(GND_net), .I1(n8142[2]), .I2(n311), .I3(n29797), 
            .O(n8123[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3699_8_lut (.I0(GND_net), .I1(n7911[5]), .I2(n542_adj_3683), 
            .I3(n29615), .O(n7896[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_5 (.CI(n29797), .I0(n8142[2]), .I1(n311), .CO(n29798));
    SB_LUT4 add_3717_4_lut (.I0(GND_net), .I1(n8142[1]), .I2(n238), .I3(n29796), 
            .O(n8123[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3684));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33963_4_lut (.I0(n21_adj_3678), .I1(n19_adj_3677), .I2(n17_adj_3676), 
            .I3(n9_adj_3675), .O(n40727));
    defparam i33963_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3717_4 (.CI(n29796), .I0(n8142[1]), .I1(n238), .CO(n29797));
    SB_LUT4 add_3717_3_lut (.I0(GND_net), .I1(n8142[0]), .I2(n165), .I3(n29795), 
            .O(n8123[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3717_3 (.CI(n29795), .I0(n8142[0]), .I1(n165), .CO(n29796));
    SB_LUT4 add_3717_2_lut (.I0(GND_net), .I1(n23_adj_3685), .I2(n92), 
            .I3(GND_net), .O(n8123[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3717_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33933_4_lut (.I0(n27_adj_3684), .I1(n15_adj_3682), .I2(n13_adj_3681), 
            .I3(n11_adj_3679), .O(n40697));
    defparam i33933_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[16]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[17]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \PID_CONTROLLER.integral_1179__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[0]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12_adj_3686), .I1(duty[17]), .I2(n35_adj_3673), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3717_2 (.CI(GND_net), .I0(n23_adj_3685), .I1(n92), .CO(n29795));
    SB_CARRY add_3699_8 (.CI(n29615), .I0(n7911[5]), .I1(n542_adj_3683), 
            .CO(n29616));
    SB_LUT4 add_3699_7_lut (.I0(GND_net), .I1(n7911[4]), .I2(n469_adj_3687), 
            .I3(n29614), .O(n7896[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34598_4_lut (.I0(n13_adj_3681), .I1(n11_adj_3679), .I2(n9_adj_3675), 
            .I3(n40749), .O(n41362));
    defparam i34598_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_3699_7 (.CI(n29614), .I0(n7911[4]), .I1(n469_adj_3687), 
            .CO(n29615));
    SB_LUT4 add_3699_6_lut (.I0(GND_net), .I1(n7911[3]), .I2(n396_adj_3688), 
            .I3(n29613), .O(n7896[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3699_6 (.CI(n29613), .I0(n7911[3]), .I1(n396_adj_3688), 
            .CO(n29614));
    SB_LUT4 add_3699_5_lut (.I0(GND_net), .I1(n7911[2]), .I2(n323_adj_3689), 
            .I3(n29612), .O(n7896[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_19_lut (.I0(GND_net), .I1(n8123[16]), .I2(GND_net), 
            .I3(n29794), .O(n8103[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_18_lut (.I0(GND_net), .I1(n8123[15]), .I2(GND_net), 
            .I3(n29793), .O(n8103[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_18 (.CI(n29793), .I0(n8123[15]), .I1(GND_net), .CO(n29794));
    SB_CARRY add_3699_5 (.CI(n29612), .I0(n7911[2]), .I1(n323_adj_3689), 
            .CO(n29613));
    SB_LUT4 add_3716_17_lut (.I0(GND_net), .I1(n8123[14]), .I2(GND_net), 
            .I3(n29792), .O(n8103[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34590_4_lut (.I0(n19_adj_3677), .I1(n17_adj_3676), .I2(n15_adj_3682), 
            .I3(n41362), .O(n41354));
    defparam i34590_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_3699_4_lut (.I0(GND_net), .I1(n7911[1]), .I2(n250_adj_3690), 
            .I3(n29611), .O(n7896[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3699_4 (.CI(n29611), .I0(n7911[1]), .I1(n250_adj_3690), 
            .CO(n29612));
    SB_CARRY add_3716_17 (.CI(n29792), .I0(n8123[14]), .I1(GND_net), .CO(n29793));
    SB_LUT4 add_3716_16_lut (.I0(GND_net), .I1(n8123[13]), .I2(GND_net), 
            .I3(n29791), .O(n8103[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_16 (.CI(n29791), .I0(n8123[13]), .I1(GND_net), .CO(n29792));
    SB_LUT4 add_3716_15_lut (.I0(GND_net), .I1(n8123[12]), .I2(GND_net), 
            .I3(n29790), .O(n8103[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35349_4_lut (.I0(n25_adj_3672), .I1(n23_adj_3671), .I2(n21_adj_3678), 
            .I3(n41354), .O(n42113));
    defparam i35349_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34906_4_lut (.I0(n31_adj_3669), .I1(n29_adj_3668), .I2(n27_adj_3684), 
            .I3(n42113), .O(n41670));
    defparam i34906_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35452_4_lut (.I0(n37_adj_3670), .I1(n35_adj_3673), .I2(n33_adj_3674), 
            .I3(n41670), .O(n42216));
    defparam i35452_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35145_3_lut (.I0(n6_adj_3691), .I1(duty[10]), .I2(n21_adj_3678), 
            .I3(GND_net), .O(n41909));   // verilog/motorControl.v(44[10:25])
    defparam i35145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35146_3_lut (.I0(n41909), .I1(duty[11]), .I2(n23_adj_3671), 
            .I3(GND_net), .O(n41910));   // verilog/motorControl.v(44[10:25])
    defparam i35146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[18]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16_adj_3692), .I1(duty[22]), .I2(n45_adj_3657), 
            .I3(GND_net), .O(n24_adj_3693));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33865_4_lut (.I0(n43_adj_3661), .I1(n25_adj_3672), .I2(n23_adj_3671), 
            .I3(n40727), .O(n40629));
    defparam i33865_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35056_4_lut (.I0(n24_adj_3693), .I1(n8_adj_3694), .I2(n45_adj_3657), 
            .I3(n40627), .O(n41820));   // verilog/motorControl.v(44[10:25])
    defparam i35056_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34351_3_lut (.I0(n41910), .I1(duty[12]), .I2(n25_adj_3672), 
            .I3(GND_net), .O(n41115));   // verilog/motorControl.v(44[10:25])
    defparam i34351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35143_3_lut (.I0(n4_adj_3695), .I1(duty[13]), .I2(n27_adj_3684), 
            .I3(GND_net), .O(n41907));   // verilog/motorControl.v(44[10:25])
    defparam i35143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[18]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3716_15 (.CI(n29790), .I0(n8123[12]), .I1(GND_net), .CO(n29791));
    SB_LUT4 i35144_3_lut (.I0(n41907), .I1(duty[14]), .I2(n29_adj_3668), 
            .I3(GND_net), .O(n41908));   // verilog/motorControl.v(44[10:25])
    defparam i35144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33925_4_lut (.I0(n33_adj_3674), .I1(n31_adj_3669), .I2(n29_adj_3668), 
            .I3(n40697), .O(n40689));
    defparam i33925_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3699_3_lut (.I0(GND_net), .I1(n7911[0]), .I2(n177_adj_3697), 
            .I3(n29610), .O(n7896[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3716_14_lut (.I0(GND_net), .I1(n8123[11]), .I2(GND_net), 
            .I3(n29789), .O(n8103[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_14 (.CI(n29789), .I0(n8123[11]), .I1(GND_net), .CO(n29790));
    SB_LUT4 i35387_4_lut (.I0(n30), .I1(n10_adj_3698), .I2(n35_adj_3673), 
            .I3(n40683), .O(n42151));   // verilog/motorControl.v(44[10:25])
    defparam i35387_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34353_3_lut (.I0(n41908), .I1(duty[15]), .I2(n31_adj_3669), 
            .I3(GND_net), .O(n41117));   // verilog/motorControl.v(44[10:25])
    defparam i34353_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3699_3 (.CI(n29610), .I0(n7911[0]), .I1(n177_adj_3697), 
            .CO(n29611));
    SB_LUT4 add_3699_2_lut (.I0(GND_net), .I1(n35_adj_3699), .I2(n104_adj_3700), 
            .I3(GND_net), .O(n7896[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3699_2 (.CI(GND_net), .I0(n35_adj_3699), .I1(n104_adj_3700), 
            .CO(n29610));
    SB_LUT4 i35520_4_lut (.I0(n41117), .I1(n42151), .I2(n35_adj_3673), 
            .I3(n40689), .O(n42284));   // verilog/motorControl.v(44[10:25])
    defparam i35520_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35521_3_lut (.I0(n42284), .I1(duty[18]), .I2(n37_adj_3670), 
            .I3(GND_net), .O(n42285));   // verilog/motorControl.v(44[10:25])
    defparam i35521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35507_3_lut (.I0(n42285), .I1(duty[19]), .I2(n39_adj_3651), 
            .I3(GND_net), .O(n42271));   // verilog/motorControl.v(44[10:25])
    defparam i35507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3698_15_lut (.I0(GND_net), .I1(n7896[12]), .I2(GND_net), 
            .I3(n29609), .O(n7880[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33870_4_lut (.I0(n43_adj_3661), .I1(n41_adj_3649), .I2(n39_adj_3651), 
            .I3(n42216), .O(n40634));
    defparam i33870_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3716_13_lut (.I0(GND_net), .I1(n8123[10]), .I2(GND_net), 
            .I3(n29788), .O(n8103[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35433_4_lut (.I0(n41115), .I1(n41820), .I2(n45_adj_3657), 
            .I3(n40629), .O(n42197));   // verilog/motorControl.v(44[10:25])
    defparam i35433_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34359_3_lut (.I0(n42271), .I1(duty[20]), .I2(n41_adj_3649), 
            .I3(GND_net), .O(n41123));   // verilog/motorControl.v(44[10:25])
    defparam i34359_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3716_13 (.CI(n29788), .I0(n8123[10]), .I1(GND_net), .CO(n29789));
    SB_LUT4 i35435_4_lut (.I0(n41123), .I1(n42197), .I2(n45_adj_3657), 
            .I3(n40634), .O(n42199));   // verilog/motorControl.v(44[10:25])
    defparam i35435_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3716_12_lut (.I0(GND_net), .I1(n8123[9]), .I2(GND_net), 
            .I3(n29787), .O(n8103[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_12 (.CI(n29787), .I0(n8123[9]), .I1(GND_net), .CO(n29788));
    SB_LUT4 add_3716_11_lut (.I0(GND_net), .I1(n8123[8]), .I2(GND_net), 
            .I3(n29786), .O(n8103[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35436_3_lut (.I0(n42199), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3502));   // verilog/motorControl.v(44[10:25])
    defparam i35436_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3698_14_lut (.I0(GND_net), .I1(n7896[11]), .I2(GND_net), 
            .I3(n29608), .O(n7880[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_11 (.CI(n29786), .I0(n8123[8]), .I1(GND_net), .CO(n29787));
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[19]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3478[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_634_i16_3_lut (.I0(n155[15]), .I1(PWMLimit[15]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i16_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[20]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3701));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3703));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3705));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3706));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3707));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3708));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3709));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[14]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3710));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3711));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3712));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3714));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3715));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3716));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3717));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3719));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3720));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3721));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3722));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3724));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33841_4_lut (.I0(n21_adj_3724), .I1(n19_adj_3722), .I2(n17_adj_3721), 
            .I3(n9_adj_3720), .O(n40605));
    defparam i33841_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33819_4_lut (.I0(n27_adj_3719), .I1(n15_adj_3717), .I2(n13_adj_3716), 
            .I3(n11_adj_3715), .O(n40583));
    defparam i33819_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_3714), 
            .I3(GND_net), .O(n12_adj_3725));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_3716), 
            .I3(GND_net), .O(n10_adj_3726));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_3725), .I1(n257[17]), .I2(n35_adj_3712), 
            .I3(GND_net), .O(n30_adj_3727));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34520_4_lut (.I0(n13_adj_3716), .I1(n11_adj_3715), .I2(n9_adj_3720), 
            .I3(n40623), .O(n41284));
    defparam i34520_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34516_4_lut (.I0(n19_adj_3722), .I1(n17_adj_3721), .I2(n15_adj_3717), 
            .I3(n41284), .O(n41280));
    defparam i34516_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35335_4_lut (.I0(n25_adj_3711), .I1(n23_adj_3710), .I2(n21_adj_3724), 
            .I3(n41280), .O(n42099));
    defparam i35335_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34874_4_lut (.I0(n31_adj_3709), .I1(n29_adj_3708), .I2(n27_adj_3719), 
            .I3(n42099), .O(n41638));
    defparam i34874_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35450_4_lut (.I0(n37_adj_3707), .I1(n35_adj_3712), .I2(n33_adj_3714), 
            .I3(n41638), .O(n42214));
    defparam i35450_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_3706), 
            .I3(GND_net), .O(n16_adj_3728));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35096_3_lut (.I0(n6_adj_3729), .I1(n257[10]), .I2(n21_adj_3724), 
            .I3(GND_net), .O(n41860));   // verilog/motorControl.v(46[19:35])
    defparam i35096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35097_3_lut (.I0(n41860), .I1(n257[11]), .I2(n23_adj_3710), 
            .I3(GND_net), .O(n41861));   // verilog/motorControl.v(46[19:35])
    defparam i35097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_3721), 
            .I3(GND_net), .O(n8_adj_3730));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_3728), .I1(n257[22]), .I2(n45_adj_3705), 
            .I3(GND_net), .O(n24_adj_3731));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33698_4_lut (.I0(n43_adj_3706), .I1(n25_adj_3711), .I2(n23_adj_3710), 
            .I3(n40605), .O(n40460));
    defparam i33698_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35058_4_lut (.I0(n24_adj_3731), .I1(n8_adj_3730), .I2(n45_adj_3705), 
            .I3(n40453), .O(n41822));   // verilog/motorControl.v(46[19:35])
    defparam i35058_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34361_3_lut (.I0(n41861), .I1(n257[12]), .I2(n25_adj_3711), 
            .I3(GND_net), .O(n41125));   // verilog/motorControl.v(46[19:35])
    defparam i34361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n40103), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_3732));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35072_3_lut (.I0(n4_adj_3732), .I1(n257[13]), .I2(n27_adj_3719), 
            .I3(GND_net), .O(n41836));   // verilog/motorControl.v(46[19:35])
    defparam i35072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35073_3_lut (.I0(n41836), .I1(n257[14]), .I2(n29_adj_3708), 
            .I3(GND_net), .O(n41837));   // verilog/motorControl.v(46[19:35])
    defparam i35073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33759_4_lut (.I0(n33_adj_3714), .I1(n31_adj_3709), .I2(n29_adj_3708), 
            .I3(n40583), .O(n40522));
    defparam i33759_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35403_4_lut (.I0(n30_adj_3727), .I1(n10_adj_3726), .I2(n35_adj_3712), 
            .I3(n40509), .O(n42167));   // verilog/motorControl.v(46[19:35])
    defparam i35403_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34363_3_lut (.I0(n41837), .I1(n257[15]), .I2(n31_adj_3709), 
            .I3(GND_net), .O(n41127));   // verilog/motorControl.v(46[19:35])
    defparam i34363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35528_4_lut (.I0(n41127), .I1(n42167), .I2(n35_adj_3712), 
            .I3(n40522), .O(n42292));   // verilog/motorControl.v(46[19:35])
    defparam i35528_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35529_3_lut (.I0(n42292), .I1(n257[18]), .I2(n37_adj_3707), 
            .I3(GND_net), .O(n42293));   // verilog/motorControl.v(46[19:35])
    defparam i35529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35498_3_lut (.I0(n42293), .I1(n257[19]), .I2(n39_adj_3703), 
            .I3(GND_net), .O(n42262));   // verilog/motorControl.v(46[19:35])
    defparam i35498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33706_4_lut (.I0(n43_adj_3706), .I1(n41_adj_3701), .I2(n39_adj_3703), 
            .I3(n42214), .O(n40468));
    defparam i33706_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35286_4_lut (.I0(n41125), .I1(n41822), .I2(n45_adj_3705), 
            .I3(n40460), .O(n42050));   // verilog/motorControl.v(46[19:35])
    defparam i35286_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34369_3_lut (.I0(n42262), .I1(n257[20]), .I2(n41_adj_3701), 
            .I3(GND_net), .O(n41133));   // verilog/motorControl.v(46[19:35])
    defparam i34369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35437_4_lut (.I0(n41133), .I1(n42050), .I2(n45_adj_3705), 
            .I3(n40468), .O(n42201));   // verilog/motorControl.v(46[19:35])
    defparam i35437_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35438_3_lut (.I0(n42201), .I1(duty[23]), .I2(n47_adj_3733), 
            .I3(GND_net), .O(n256_adj_3571));   // verilog/motorControl.v(46[19:35])
    defparam i35438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_634_i17_3_lut (.I0(n155[16]), .I1(PWMLimit[16]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i17_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[21]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3734));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[19]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[20]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3737));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3738));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3716_10_lut (.I0(GND_net), .I1(n8123[7]), .I2(GND_net), 
            .I3(n29785), .O(n8103[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3698_14 (.CI(n29608), .I0(n7896[11]), .I1(GND_net), .CO(n29609));
    SB_LUT4 add_3698_13_lut (.I0(GND_net), .I1(n7896[10]), .I2(GND_net), 
            .I3(n29607), .O(n7880[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_3892[23]), .I3(n28201), .O(\PID_CONTROLLER.err_23__N_3379 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_3892[22]), .I3(n28200), .O(\PID_CONTROLLER.err_23__N_3379 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_10 (.CI(n29785), .I0(n8123[7]), .I1(GND_net), .CO(n29786));
    SB_CARRY add_3698_13 (.CI(n29607), .I0(n7896[10]), .I1(GND_net), .CO(n29608));
    SB_LUT4 add_3698_12_lut (.I0(GND_net), .I1(n7896[9]), .I2(GND_net), 
            .I3(n29606), .O(n7880[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_3741));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[21]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_3743));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_3744));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3698_12 (.CI(n29606), .I0(n7896[9]), .I1(GND_net), .CO(n29607));
    SB_LUT4 add_3698_11_lut (.I0(GND_net), .I1(n7896[8]), .I2(GND_net), 
            .I3(n29605), .O(n7880[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_3745));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3716_9_lut (.I0(GND_net), .I1(n8123[6]), .I2(GND_net), 
            .I3(n29784), .O(n8103[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_3746));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3698_11 (.CI(n29605), .I0(n7896[8]), .I1(GND_net), .CO(n29606));
    SB_LUT4 add_3698_10_lut (.I0(GND_net), .I1(n7896[7]), .I2(GND_net), 
            .I3(n29604), .O(n7880[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_9 (.CI(n29784), .I0(n8123[6]), .I1(GND_net), .CO(n29785));
    SB_CARRY add_3698_10 (.CI(n29604), .I0(n7896[7]), .I1(GND_net), .CO(n29605));
    SB_LUT4 add_3698_9_lut (.I0(GND_net), .I1(n7896[6]), .I2(GND_net), 
            .I3(n29603), .O(n7880[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3698_9 (.CI(n29603), .I0(n7896[6]), .I1(GND_net), .CO(n29604));
    SB_LUT4 add_3716_8_lut (.I0(GND_net), .I1(n8123[5]), .I2(n527), .I3(n29783), 
            .O(n8103[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_8 (.CI(n29783), .I0(n8123[5]), .I1(n527), .CO(n29784));
    SB_LUT4 add_3698_8_lut (.I0(GND_net), .I1(n7896[5]), .I2(n539_adj_3747), 
            .I3(n29602), .O(n7880[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3698_8 (.CI(n29602), .I0(n7896[5]), .I1(n539_adj_3747), 
            .CO(n29603));
    SB_LUT4 add_3698_7_lut (.I0(GND_net), .I1(n7896[4]), .I2(n466_adj_3746), 
            .I3(n29601), .O(n7880[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3698_7 (.CI(n29601), .I0(n7896[4]), .I1(n466_adj_3746), 
            .CO(n29602));
    SB_LUT4 add_3716_7_lut (.I0(GND_net), .I1(n8123[4]), .I2(n454), .I3(n29782), 
            .O(n8103[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3698_6_lut (.I0(GND_net), .I1(n7896[3]), .I2(n393_adj_3745), 
            .I3(n29600), .O(n7880[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_7 (.CI(n29782), .I0(n8123[4]), .I1(n454), .CO(n29783));
    SB_LUT4 add_3716_6_lut (.I0(GND_net), .I1(n8123[3]), .I2(n381), .I3(n29781), 
            .O(n8103[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3698_6 (.CI(n29600), .I0(n7896[3]), .I1(n393_adj_3745), 
            .CO(n29601));
    SB_CARRY add_3716_6 (.CI(n29781), .I0(n8123[3]), .I1(n381), .CO(n29782));
    SB_LUT4 add_3716_5_lut (.I0(GND_net), .I1(n8123[2]), .I2(n308), .I3(n29780), 
            .O(n8103[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_3747));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3716_5 (.CI(n29780), .I0(n8123[2]), .I1(n308), .CO(n29781));
    SB_LUT4 add_3698_5_lut (.I0(GND_net), .I1(n7896[2]), .I2(n320_adj_3744), 
            .I3(n29599), .O(n7880[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n28200), .I0(motor_state[22]), 
            .I1(n1_adj_3892[22]), .CO(n28201));
    SB_CARRY add_3698_5 (.CI(n29599), .I0(n7896[2]), .I1(n320_adj_3744), 
            .CO(n29600));
    SB_LUT4 add_3716_4_lut (.I0(GND_net), .I1(n8123[1]), .I2(n235), .I3(n29779), 
            .O(n8103[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3698_4_lut (.I0(GND_net), .I1(n7896[1]), .I2(n247_adj_3743), 
            .I3(n29598), .O(n7880[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3698_4 (.CI(n29598), .I0(n7896[1]), .I1(n247_adj_3743), 
            .CO(n29599));
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_3892[21]), .I3(n28199), .O(\PID_CONTROLLER.err_23__N_3379 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3716_4 (.CI(n29779), .I0(n8123[1]), .I1(n235), .CO(n29780));
    SB_LUT4 add_3698_3_lut (.I0(GND_net), .I1(n7896[0]), .I2(n174_adj_3741), 
            .I3(n29597), .O(n7880[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n28199), .I0(motor_state[21]), 
            .I1(n1_adj_3892[21]), .CO(n28200));
    SB_CARRY add_3698_3 (.CI(n29597), .I0(n7896[0]), .I1(n174_adj_3741), 
            .CO(n29598));
    SB_LUT4 add_3716_3_lut (.I0(GND_net), .I1(n8123[0]), .I2(n162), .I3(n29778), 
            .O(n8103[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3698_2_lut (.I0(GND_net), .I1(n32_adj_3738), .I2(n101_adj_3737), 
            .I3(GND_net), .O(n7880[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3698_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3698_2 (.CI(GND_net), .I0(n32_adj_3738), .I1(n101_adj_3737), 
            .CO(n29597));
    SB_CARRY add_3716_3 (.CI(n29778), .I0(n8123[0]), .I1(n162), .CO(n29779));
    SB_LUT4 add_3697_16_lut (.I0(GND_net), .I1(n7880[13]), .I2(GND_net), 
            .I3(n29596), .O(n7863[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3697_15_lut (.I0(GND_net), .I1(n7880[12]), .I2(GND_net), 
            .I3(n29595), .O(n7863[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_3892[20]), .I3(n28198), .O(\PID_CONTROLLER.err_23__N_3379 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n28198), .I0(motor_state[20]), 
            .I1(n1_adj_3892[20]), .CO(n28199));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_3892[19]), .I3(n28197), .O(\PID_CONTROLLER.err_23__N_3379 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n28197), .I0(motor_state[19]), 
            .I1(n1_adj_3892[19]), .CO(n28198));
    SB_LUT4 add_3716_2_lut (.I0(GND_net), .I1(n20_adj_3734), .I2(n89), 
            .I3(GND_net), .O(n8103[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3716_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_15 (.CI(n29595), .I0(n7880[12]), .I1(GND_net), .CO(n29596));
    SB_LUT4 add_3697_14_lut (.I0(GND_net), .I1(n7880[11]), .I2(GND_net), 
            .I3(n29594), .O(n7863[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_14 (.CI(n29594), .I0(n7880[11]), .I1(GND_net), .CO(n29595));
    SB_CARRY add_3716_2 (.CI(GND_net), .I0(n20_adj_3734), .I1(n89), .CO(n29778));
    SB_LUT4 add_3697_13_lut (.I0(GND_net), .I1(n7880[10]), .I2(GND_net), 
            .I3(n29593), .O(n7863[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[22]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3715_20_lut (.I0(GND_net), .I1(n8103[17]), .I2(GND_net), 
            .I3(n29777), .O(n8082[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3715_19_lut (.I0(GND_net), .I1(n8103[16]), .I2(GND_net), 
            .I3(n29776), .O(n8082[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_13 (.CI(n29593), .I0(n7880[10]), .I1(GND_net), .CO(n29594));
    SB_LUT4 mux_634_i14_3_lut (.I0(n155[13]), .I1(PWMLimit[13]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i14_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_3892[18]), .I3(n28196), .O(\PID_CONTROLLER.err_23__N_3379 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3355[1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_3697_12_lut (.I0(GND_net), .I1(n7880[9]), .I2(GND_net), 
            .I3(n29592), .O(n7863[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3715_19 (.CI(n29776), .I0(n8103[16]), .I1(GND_net), .CO(n29777));
    SB_CARRY state_23__I_0_add_2_20 (.CI(n28196), .I0(motor_state[18]), 
            .I1(n1_adj_3892[18]), .CO(n28197));
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_3892[17]), .I3(n28195), .O(\PID_CONTROLLER.err_23__N_3379 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[23]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3573));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3572));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[22]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[23]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3715_18_lut (.I0(GND_net), .I1(n8103[15]), .I2(GND_net), 
            .I3(n29775), .O(n8082[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_12 (.CI(n29592), .I0(n7880[9]), .I1(GND_net), .CO(n29593));
    SB_CARRY state_23__I_0_add_2_19 (.CI(n28195), .I0(motor_state[17]), 
            .I1(n1_adj_3892[17]), .CO(n28196));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_3892[16]), .I3(n28194), .O(\PID_CONTROLLER.err_23__N_3379 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3697_11_lut (.I0(GND_net), .I1(n7880[8]), .I2(GND_net), 
            .I3(n29591), .O(n7863[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3355[2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3355[3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3355[4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3355[5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3355[6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3355[7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3355[8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3355[9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3355[10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3355[11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3355[12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3355[13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3355[14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3355[15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3355[16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3355[17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3355[18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3355[19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3355[20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3355[21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3355[22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3355[23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_3715_18 (.CI(n29775), .I0(n8103[15]), .I1(GND_net), .CO(n29776));
    SB_CARRY add_3697_11 (.CI(n29591), .I0(n7880[8]), .I1(GND_net), .CO(n29592));
    SB_LUT4 add_3697_10_lut (.I0(GND_net), .I1(n7880[7]), .I2(GND_net), 
            .I3(n29590), .O(n7863[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3715_17_lut (.I0(GND_net), .I1(n8103[14]), .I2(GND_net), 
            .I3(n29774), .O(n8082[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_10 (.CI(n29590), .I0(n7880[7]), .I1(GND_net), .CO(n29591));
    SB_LUT4 add_3697_9_lut (.I0(GND_net), .I1(n7880[6]), .I2(GND_net), 
            .I3(n29589), .O(n7863[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_17 (.CI(n29774), .I0(n8103[14]), .I1(GND_net), .CO(n29775));
    SB_CARRY add_3697_9 (.CI(n29589), .I0(n7880[6]), .I1(GND_net), .CO(n29590));
    SB_CARRY state_23__I_0_add_2_18 (.CI(n28194), .I0(motor_state[16]), 
            .I1(n1_adj_3892[16]), .CO(n28195));
    SB_LUT4 add_3697_8_lut (.I0(GND_net), .I1(n7880[5]), .I2(n536), .I3(n29588), 
            .O(n7863[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_8 (.CI(n29588), .I0(n7880[5]), .I1(n536), .CO(n29589));
    SB_LUT4 add_3715_16_lut (.I0(GND_net), .I1(n8103[13]), .I2(GND_net), 
            .I3(n29773), .O(n8082[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_3892[15]), .I3(n28193), .O(\PID_CONTROLLER.err_23__N_3379 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n28193), .I0(motor_state[15]), 
            .I1(n1_adj_3892[15]), .CO(n28194));
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_3892[14]), .I3(n28192), .O(\PID_CONTROLLER.err_23__N_3379 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3697_7_lut (.I0(GND_net), .I1(n7880[4]), .I2(n463), .I3(n29587), 
            .O(n7863[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_16 (.CI(n29773), .I0(n8103[13]), .I1(GND_net), .CO(n29774));
    SB_CARRY add_3697_7 (.CI(n29587), .I0(n7880[4]), .I1(n463), .CO(n29588));
    SB_CARRY state_23__I_0_add_2_16 (.CI(n28192), .I0(motor_state[14]), 
            .I1(n1_adj_3892[14]), .CO(n28193));
    SB_LUT4 add_3697_6_lut (.I0(GND_net), .I1(n7880[3]), .I2(n390), .I3(n29586), 
            .O(n7863[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_3892[13]), .I3(n28191), .O(\PID_CONTROLLER.err_23__N_3379 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n28191), .I0(motor_state[13]), 
            .I1(n1_adj_3892[13]), .CO(n28192));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_3892[12]), .I3(n28190), .O(\PID_CONTROLLER.err_23__N_3379 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3715_15_lut (.I0(GND_net), .I1(n8103[12]), .I2(GND_net), 
            .I3(n29772), .O(n8082[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n28190), .I0(motor_state[12]), 
            .I1(n1_adj_3892[12]), .CO(n28191));
    SB_CARRY add_3697_6 (.CI(n29586), .I0(n7880[3]), .I1(n390), .CO(n29587));
    SB_CARRY add_3715_15 (.CI(n29772), .I0(n8103[12]), .I1(GND_net), .CO(n29773));
    SB_LUT4 add_3715_14_lut (.I0(GND_net), .I1(n8103[11]), .I2(GND_net), 
            .I3(n29771), .O(n8082[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_14 (.CI(n29771), .I0(n8103[11]), .I1(GND_net), .CO(n29772));
    SB_LUT4 add_3715_13_lut (.I0(GND_net), .I1(n8103[10]), .I2(GND_net), 
            .I3(n29770), .O(n8082[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_3892[11]), .I3(n28189), .O(\PID_CONTROLLER.err_23__N_3379 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_13 (.CI(n29770), .I0(n8103[10]), .I1(GND_net), .CO(n29771));
    SB_LUT4 add_3715_12_lut (.I0(GND_net), .I1(n8103[9]), .I2(GND_net), 
            .I3(n29769), .O(n8082[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3697_5_lut (.I0(GND_net), .I1(n7880[2]), .I2(n317), .I3(n29585), 
            .O(n7863[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_5 (.CI(n29585), .I0(n7880[2]), .I1(n317), .CO(n29586));
    SB_CARRY state_23__I_0_add_2_13 (.CI(n28189), .I0(motor_state[11]), 
            .I1(n1_adj_3892[11]), .CO(n28190));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_3892[10]), .I3(n28188), .O(\PID_CONTROLLER.err_23__N_3379 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n28188), .I0(motor_state[10]), 
            .I1(n1_adj_3892[10]), .CO(n28189));
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3700));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3715_12 (.CI(n29769), .I0(n8103[9]), .I1(GND_net), .CO(n29770));
    SB_LUT4 add_3715_11_lut (.I0(GND_net), .I1(n8103[8]), .I2(GND_net), 
            .I3(n29768), .O(n8082[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_3892[9]), .I3(n28187), .O(\PID_CONTROLLER.err_23__N_3379 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n28187), .I0(motor_state[9]), .I1(n1_adj_3892[9]), 
            .CO(n28188));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_3892[8]), .I3(n28186), .O(\PID_CONTROLLER.err_23__N_3379 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n28186), .I0(motor_state[8]), .I1(n1_adj_3892[8]), 
            .CO(n28187));
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3699));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_3892[7]), .I3(n28185), .O(\PID_CONTROLLER.err_23__N_3379 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3697_4_lut (.I0(GND_net), .I1(n7880[1]), .I2(n244), .I3(n29584), 
            .O(n7863[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_11 (.CI(n29768), .I0(n8103[8]), .I1(GND_net), .CO(n29769));
    SB_LUT4 add_3715_10_lut (.I0(GND_net), .I1(n8103[7]), .I2(GND_net), 
            .I3(n29767), .O(n8082[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_9 (.CI(n28185), .I0(motor_state[7]), .I1(n1_adj_3892[7]), 
            .CO(n28186));
    SB_CARRY add_3697_4 (.CI(n29584), .I0(n7880[1]), .I1(n244), .CO(n29585));
    SB_CARRY add_3715_10 (.CI(n29767), .I0(n8103[7]), .I1(GND_net), .CO(n29768));
    SB_LUT4 add_3715_9_lut (.I0(GND_net), .I1(n8103[6]), .I2(GND_net), 
            .I3(n29766), .O(n8082[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_9 (.CI(n29766), .I0(n8103[6]), .I1(GND_net), .CO(n29767));
    SB_LUT4 add_3715_8_lut (.I0(GND_net), .I1(n8103[5]), .I2(n524), .I3(n29765), 
            .O(n8082[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_8 (.CI(n29765), .I0(n8103[5]), .I1(n524), .CO(n29766));
    SB_LUT4 add_3697_3_lut (.I0(GND_net), .I1(n7880[0]), .I2(n171), .I3(n29583), 
            .O(n7863[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_3 (.CI(n29583), .I0(n7880[0]), .I1(n171), .CO(n29584));
    SB_LUT4 add_3715_7_lut (.I0(GND_net), .I1(n8103[4]), .I2(n451), .I3(n29764), 
            .O(n8082[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_7 (.CI(n29764), .I0(n8103[4]), .I1(n451), .CO(n29765));
    SB_LUT4 add_3697_2_lut (.I0(GND_net), .I1(n29_adj_3584), .I2(n98), 
            .I3(GND_net), .O(n7863[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3697_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_3892[6]), .I3(n28184), .O(\PID_CONTROLLER.err_23__N_3379 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3697_2 (.CI(GND_net), .I0(n29_adj_3584), .I1(n98), .CO(n29583));
    SB_LUT4 add_3696_17_lut (.I0(GND_net), .I1(n7863[14]), .I2(GND_net), 
            .I3(n29582), .O(n7845[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_16_lut (.I0(GND_net), .I1(n7863[13]), .I2(GND_net), 
            .I3(n29581), .O(n7845[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3715_6_lut (.I0(GND_net), .I1(n8103[3]), .I2(n378), .I3(n29763), 
            .O(n8082[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_16 (.CI(n29581), .I0(n7863[13]), .I1(GND_net), .CO(n29582));
    SB_CARRY state_23__I_0_add_2_8 (.CI(n28184), .I0(motor_state[6]), .I1(n1_adj_3892[6]), 
            .CO(n28185));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_3892[5]), .I3(n28183), .O(\PID_CONTROLLER.err_23__N_3379 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n28183), .I0(motor_state[5]), .I1(n1_adj_3892[5]), 
            .CO(n28184));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_3892[4]), .I3(n28182), .O(\PID_CONTROLLER.err_23__N_3379 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_15_lut (.I0(GND_net), .I1(n7863[12]), .I2(GND_net), 
            .I3(n29580), .O(n7845[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3715_6 (.CI(n29763), .I0(n8103[3]), .I1(n378), .CO(n29764));
    SB_CARRY state_23__I_0_add_2_6 (.CI(n28182), .I0(motor_state[4]), .I1(n1_adj_3892[4]), 
            .CO(n28183));
    SB_LUT4 add_3715_5_lut (.I0(GND_net), .I1(n8103[2]), .I2(n305), .I3(n29762), 
            .O(n8082[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_15 (.CI(n29580), .I0(n7863[12]), .I1(GND_net), .CO(n29581));
    SB_CARRY add_3715_5 (.CI(n29762), .I0(n8103[2]), .I1(n305), .CO(n29763));
    SB_LUT4 add_3696_14_lut (.I0(GND_net), .I1(n7863[11]), .I2(GND_net), 
            .I3(n29579), .O(n7845[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_14 (.CI(n29579), .I0(n7863[11]), .I1(GND_net), .CO(n29580));
    SB_LUT4 add_3696_13_lut (.I0(GND_net), .I1(n7863[10]), .I2(GND_net), 
            .I3(n29578), .O(n7845[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_3697));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3696_13 (.CI(n29578), .I0(n7863[10]), .I1(GND_net), .CO(n29579));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_3892[3]), .I3(n28181), .O(\PID_CONTROLLER.err_23__N_3379 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n28181), .I0(motor_state[3]), .I1(n1_adj_3892[3]), 
            .CO(n28182));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_3892[2]), .I3(n28180), .O(\PID_CONTROLLER.err_23__N_3379 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_4 (.CI(n28180), .I0(motor_state[2]), .I1(n1_adj_3892[2]), 
            .CO(n28181));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_3892[1]), .I3(n28179), .O(\PID_CONTROLLER.err_23__N_3379 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3715_4_lut (.I0(GND_net), .I1(n8103[1]), .I2(n232), .I3(n29761), 
            .O(n8082[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_12_lut (.I0(GND_net), .I1(n7863[9]), .I2(GND_net), 
            .I3(n29577), .O(n7845[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n28179), .I0(motor_state[1]), .I1(n1_adj_3892[1]), 
            .CO(n28180));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_3892[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3379 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_12 (.CI(n29577), .I0(n7863[9]), .I1(GND_net), .CO(n29578));
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_3892[0]), 
            .CO(n28179));
    SB_CARRY add_3715_4 (.CI(n29761), .I0(n8103[1]), .I1(n232), .CO(n29762));
    SB_LUT4 add_3696_11_lut (.I0(GND_net), .I1(n7863[8]), .I2(GND_net), 
            .I3(n29576), .O(n7845[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_11 (.CI(n29576), .I0(n7863[8]), .I1(GND_net), .CO(n29577));
    SB_LUT4 add_3715_3_lut (.I0(GND_net), .I1(n8103[0]), .I2(n159), .I3(n29760), 
            .O(n8082[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_10_lut (.I0(GND_net), .I1(n7863[7]), .I2(GND_net), 
            .I3(n29575), .O(n7845[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1[23]), 
            .I3(n28178), .O(n47_adj_3733)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n28177), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_10 (.CI(n29575), .I0(n7863[7]), .I1(GND_net), .CO(n29576));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n28177), .I0(GND_net), .I1(n1[22]), 
            .CO(n28178));
    SB_CARRY add_3715_3 (.CI(n29760), .I0(n8103[0]), .I1(n159), .CO(n29761));
    SB_LUT4 add_3715_2_lut (.I0(GND_net), .I1(n17_adj_3754), .I2(n86), 
            .I3(GND_net), .O(n8082[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3715_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_9_lut (.I0(GND_net), .I1(n7863[6]), .I2(GND_net), 
            .I3(n29574), .O(n7845[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_9 (.CI(n29574), .I0(n7863[6]), .I1(GND_net), .CO(n29575));
    SB_CARRY add_3715_2 (.CI(GND_net), .I0(n17_adj_3754), .I1(n86), .CO(n29760));
    SB_LUT4 add_3696_8_lut (.I0(GND_net), .I1(n7863[5]), .I2(n533_adj_3755), 
            .I3(n29573), .O(n7845[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_8 (.CI(n29573), .I0(n7863[5]), .I1(n533_adj_3755), 
            .CO(n29574));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n28176), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3714_21_lut (.I0(GND_net), .I1(n8082[18]), .I2(GND_net), 
            .I3(n29759), .O(n8060[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_7_lut (.I0(GND_net), .I1(n7863[4]), .I2(n460_adj_3757), 
            .I3(n29572), .O(n7845[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_7 (.CI(n29572), .I0(n7863[4]), .I1(n460_adj_3757), 
            .CO(n29573));
    SB_LUT4 add_3714_20_lut (.I0(GND_net), .I1(n8082[17]), .I2(GND_net), 
            .I3(n29758), .O(n8060[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_6_lut (.I0(GND_net), .I1(n7863[3]), .I2(n387_adj_3758), 
            .I3(n29571), .O(n7845[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_6 (.CI(n29571), .I0(n7863[3]), .I1(n387_adj_3758), 
            .CO(n29572));
    SB_CARRY add_3714_20 (.CI(n29758), .I0(n8082[17]), .I1(GND_net), .CO(n29759));
    SB_LUT4 add_3696_5_lut (.I0(GND_net), .I1(n7863[2]), .I2(n314_adj_3759), 
            .I3(n29570), .O(n7845[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_5 (.CI(n29570), .I0(n7863[2]), .I1(n314_adj_3759), 
            .CO(n29571));
    SB_LUT4 add_3714_19_lut (.I0(GND_net), .I1(n8082[16]), .I2(GND_net), 
            .I3(n29757), .O(n8060[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3696_4_lut (.I0(GND_net), .I1(n7863[1]), .I2(n241_adj_3760), 
            .I3(n29569), .O(n7845[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_4 (.CI(n29569), .I0(n7863[1]), .I1(n241_adj_3760), 
            .CO(n29570));
    SB_CARRY unary_minus_16_add_3_23 (.CI(n28176), .I0(GND_net), .I1(n1[21]), 
            .CO(n28177));
    SB_LUT4 add_3696_3_lut (.I0(GND_net), .I1(n7863[0]), .I2(n168_adj_3761), 
            .I3(n29568), .O(n7845[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3714_19 (.CI(n29757), .I0(n8082[16]), .I1(GND_net), .CO(n29758));
    SB_LUT4 add_3714_18_lut (.I0(GND_net), .I1(n8082[15]), .I2(GND_net), 
            .I3(n29756), .O(n8060[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3696_3 (.CI(n29568), .I0(n7863[0]), .I1(n168_adj_3761), 
            .CO(n29569));
    SB_CARRY add_3714_18 (.CI(n29756), .I0(n8082[15]), .I1(GND_net), .CO(n29757));
    SB_LUT4 add_3696_2_lut (.I0(GND_net), .I1(n26_adj_3762), .I2(n95_adj_3763), 
            .I3(GND_net), .O(n7845[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3696_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_3690));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_3689));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_3688));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_3687));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3696_2 (.CI(GND_net), .I0(n26_adj_3762), .I1(n95_adj_3763), 
            .CO(n29568));
    SB_LUT4 add_3714_17_lut (.I0(GND_net), .I1(n8082[14]), .I2(GND_net), 
            .I3(n29755), .O(n8060[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_3764));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_3765));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_3766));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33754_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n40517));
    defparam i33754_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i33588_3_lut (.I0(n11_adj_3766), .I1(n9_adj_3765), .I2(n40517), 
            .I3(GND_net), .O(n40350));
    defparam i33588_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_443_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n44041));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_443_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34796_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n44041), 
            .I2(IntegralLimit[7]), .I3(n40350), .O(n41560));
    defparam i34796_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34223_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3764), 
            .I2(IntegralLimit[9]), .I3(n41560), .O(n40987));
    defparam i34223_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_425_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n44023));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_425_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34179_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3764), 
            .I2(IntegralLimit[9]), .I3(n9_adj_3765), .O(n40943));
    defparam i34179_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_3695_18_lut (.I0(GND_net), .I1(n7845[15]), .I2(GND_net), 
            .I3(n29567), .O(n7826[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34750_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n44023), 
            .I2(IntegralLimit[11]), .I3(n40943), .O(n41514));
    defparam i34750_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_419_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n44017));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_419_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34048_4_lut (.I0(n27), .I1(n15_adj_3603), .I2(n13_adj_3605), 
            .I3(n11_adj_3613), .O(n40812));
    defparam i34048_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34069_4_lut (.I0(n21_adj_3581), .I1(n19), .I2(n17_adj_3597), 
            .I3(n9_adj_3616), .O(n40833));
    defparam i34069_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_3767));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i33989_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n40753));
    defparam i33989_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_3597), .I3(GND_net), 
            .O(n8_adj_3768));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_3767), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_3769));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34109_2_lut (.I0(n7_adj_3625), .I1(n5_adj_3628), .I2(GND_net), 
            .I3(GND_net), .O(n40873));
    defparam i34109_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i34704_4_lut (.I0(n13_adj_3605), .I1(n11_adj_3613), .I2(n9_adj_3616), 
            .I3(n40873), .O(n41468));
    defparam i34704_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34688_4_lut (.I0(n19), .I1(n17_adj_3597), .I2(n15_adj_3603), 
            .I3(n41468), .O(n41452));
    defparam i34688_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35369_4_lut (.I0(n25_adj_3577), .I1(n23), .I2(n21_adj_3581), 
            .I3(n41452), .O(n42133));
    defparam i35369_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34958_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n42133), 
            .O(n41722));
    defparam i34958_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35456_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n41722), 
            .O(n42220));
    defparam i35456_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34273_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n44041), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3766), .O(n41037));
    defparam i34273_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_412_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n44010));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_412_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34738_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n44010), 
            .I2(IntegralLimit[14]), .I3(n41037), .O(n41502));
    defparam i34738_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_407_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n44005));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_407_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_3770));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34135_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n40899));
    defparam i34135_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_430_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n44028));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_430_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3771));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_3770), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_3772));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35002_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n44023), 
            .I2(IntegralLimit[11]), .I3(n40987), .O(n41766));
    defparam i35002_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34158_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n44017), 
            .I2(IntegralLimit[13]), .I3(n41766), .O(n40922));
    defparam i34158_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_410_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n44008));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_410_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34996_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n44008), 
            .I2(IntegralLimit[15]), .I3(n40922), .O(n41760));
    defparam i34996_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_436_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n44034));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_436_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35379_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n44034), 
            .I2(IntegralLimit[17]), .I3(n41760), .O(n42143));
    defparam i35379_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_401_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n43999));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_401_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35541_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n43999), 
            .I2(IntegralLimit[19]), .I3(n42143), .O(n42305));
    defparam i35541_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_398_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n43996));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_398_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_3773));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34111_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n40875));
    defparam i34111_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_3773), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_3774));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3775));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35159_3_lut (.I0(n6_adj_3775), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n41923));   // verilog/motorControl.v(39[10:34])
    defparam i35159_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35160_3_lut (.I0(n41923), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n41924));   // verilog/motorControl.v(39[10:34])
    defparam i35160_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34113_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n44017), 
            .I2(IntegralLimit[21]), .I3(n41514), .O(n40877));
    defparam i34113_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i35052_4_lut (.I0(n24_adj_3774), .I1(n8_adj_3776), .I2(n43994), 
            .I3(n40875), .O(n41816));   // verilog/motorControl.v(39[10:34])
    defparam i35052_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34331_3_lut (.I0(n41924), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n41095));   // verilog/motorControl.v(39[10:34])
    defparam i34331_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3454 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_3634), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_3777));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i35151_3_lut (.I0(n4_adj_3777), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n41915));   // verilog/motorControl.v(39[38:63])
    defparam i35151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35152_3_lut (.I0(n41915), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n41916));   // verilog/motorControl.v(39[38:63])
    defparam i35152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_3778));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n28175), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34033_2_lut (.I0(n33), .I1(n15_adj_3603), .I2(GND_net), .I3(GND_net), 
            .O(n40797));
    defparam i34033_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_3714_17 (.CI(n29755), .I0(n8082[14]), .I1(GND_net), .CO(n29756));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_3605), .I3(GND_net), 
            .O(n10_adj_3780));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_3714_16_lut (.I0(GND_net), .I1(n8082[13]), .I2(GND_net), 
            .I3(n29754), .O(n8060[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3695_17_lut (.I0(GND_net), .I1(n7845[14]), .I2(GND_net), 
            .I3(n29566), .O(n7826[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_17 (.CI(n29566), .I0(n7845[14]), .I1(GND_net), .CO(n29567));
    SB_LUT4 add_3695_16_lut (.I0(GND_net), .I1(n7845[13]), .I2(GND_net), 
            .I3(n29565), .O(n7826[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_16 (.CI(n29565), .I0(n7845[13]), .I1(GND_net), .CO(n29566));
    SB_LUT4 add_3695_15_lut (.I0(GND_net), .I1(n7845[12]), .I2(GND_net), 
            .I3(n29564), .O(n7826[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_3778), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_3781));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_3695_15 (.CI(n29564), .I0(n7845[12]), .I1(GND_net), .CO(n29565));
    SB_CARRY add_3714_16 (.CI(n29754), .I0(n8082[13]), .I1(GND_net), .CO(n29755));
    SB_LUT4 add_3695_14_lut (.I0(GND_net), .I1(n7845[11]), .I2(GND_net), 
            .I3(n29563), .O(n7826[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3714_15_lut (.I0(GND_net), .I1(n8082[12]), .I2(GND_net), 
            .I3(n29753), .O(n8060[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_14 (.CI(n29563), .I0(n7845[11]), .I1(GND_net), .CO(n29564));
    SB_LUT4 add_3695_13_lut (.I0(GND_net), .I1(n7845[10]), .I2(GND_net), 
            .I3(n29562), .O(n7826[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34039_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n40812), 
            .O(n40803));
    defparam i34039_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35385_4_lut (.I0(n30_adj_3781), .I1(n10_adj_3780), .I2(n35), 
            .I3(n40797), .O(n42149));   // verilog/motorControl.v(39[38:63])
    defparam i35385_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n28175), .I0(GND_net), .I1(n1[20]), 
            .CO(n28176));
    SB_LUT4 i34343_3_lut (.I0(n41916), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n41107));   // verilog/motorControl.v(39[38:63])
    defparam i34343_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3695_13 (.CI(n29562), .I0(n7845[10]), .I1(GND_net), .CO(n29563));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n28174), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3695_12_lut (.I0(GND_net), .I1(n7845[9]), .I2(GND_net), 
            .I3(n29561), .O(n7826[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35518_4_lut (.I0(n41107), .I1(n42149), .I2(n35), .I3(n40803), 
            .O(n42282));   // verilog/motorControl.v(39[38:63])
    defparam i35518_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3714_15 (.CI(n29753), .I0(n8082[12]), .I1(GND_net), .CO(n29754));
    SB_LUT4 add_3714_14_lut (.I0(GND_net), .I1(n8082[11]), .I2(GND_net), 
            .I3(n29752), .O(n8060[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_12 (.CI(n29561), .I0(n7845[9]), .I1(GND_net), .CO(n29562));
    SB_LUT4 add_3695_11_lut (.I0(GND_net), .I1(n7845[8]), .I2(GND_net), 
            .I3(n29560), .O(n7826[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35519_3_lut (.I0(n42282), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n42283));   // verilog/motorControl.v(39[38:63])
    defparam i35519_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3695_11 (.CI(n29560), .I0(n7845[8]), .I1(GND_net), .CO(n29561));
    SB_LUT4 i35509_3_lut (.I0(n42283), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n42273));   // verilog/motorControl.v(39[38:63])
    defparam i35509_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3714_14 (.CI(n29752), .I0(n8082[11]), .I1(GND_net), .CO(n29753));
    SB_LUT4 add_3695_10_lut (.I0(GND_net), .I1(n7845[7]), .I2(GND_net), 
            .I3(n29559), .O(n7826[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_10 (.CI(n29559), .I0(n7845[7]), .I1(GND_net), .CO(n29560));
    SB_LUT4 add_3714_13_lut (.I0(GND_net), .I1(n8082[10]), .I2(GND_net), 
            .I3(n29751), .O(n8060[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3695_9_lut (.I0(GND_net), .I1(n7845[6]), .I2(GND_net), 
            .I3(n29558), .O(n7826[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_9 (.CI(n29558), .I0(n7845[6]), .I1(GND_net), .CO(n29559));
    SB_CARRY add_3714_13 (.CI(n29751), .I0(n8082[10]), .I1(GND_net), .CO(n29752));
    SB_LUT4 add_3695_8_lut (.I0(GND_net), .I1(n7845[5]), .I2(n530_adj_3783), 
            .I3(n29557), .O(n7826[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_3625), .I3(GND_net), 
            .O(n6_adj_3784));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_3695_8 (.CI(n29557), .I0(n7845[5]), .I1(n530_adj_3783), 
            .CO(n29558));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n28174), .I0(GND_net), .I1(n1[19]), 
            .CO(n28175));
    SB_LUT4 i35153_3_lut (.I0(n6_adj_3784), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_3581), .I3(GND_net), .O(n41917));   // verilog/motorControl.v(39[38:63])
    defparam i35153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3714_12_lut (.I0(GND_net), .I1(n8082[9]), .I2(GND_net), 
            .I3(n29750), .O(n8060[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3695_7_lut (.I0(GND_net), .I1(n7845[4]), .I2(n457_adj_3785), 
            .I3(n29556), .O(n7826[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_7 (.CI(n29556), .I0(n7845[4]), .I1(n457_adj_3785), 
            .CO(n29557));
    SB_CARRY add_3714_12 (.CI(n29750), .I0(n8082[9]), .I1(GND_net), .CO(n29751));
    SB_LUT4 add_3695_6_lut (.I0(GND_net), .I1(n7845[3]), .I2(n384_adj_3786), 
            .I3(n29555), .O(n7826[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35154_3_lut (.I0(n41917), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23), .I3(GND_net), .O(n41918));   // verilog/motorControl.v(39[38:63])
    defparam i35154_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3695_6 (.CI(n29555), .I0(n7845[3]), .I1(n384_adj_3786), 
            .CO(n29556));
    SB_LUT4 add_3695_5_lut (.I0(GND_net), .I1(n7845[2]), .I2(n311_adj_3787), 
            .I3(n29554), .O(n7826[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n28173), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33993_4_lut (.I0(n43), .I1(n25_adj_3577), .I2(n23), .I3(n40833), 
            .O(n40757));
    defparam i33993_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n28173), .I0(GND_net), .I1(n1[18]), 
            .CO(n28174));
    SB_LUT4 i35054_4_lut (.I0(n24_adj_3769), .I1(n8_adj_3768), .I2(n45), 
            .I3(n40753), .O(n41818));   // verilog/motorControl.v(39[38:63])
    defparam i35054_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3714_11_lut (.I0(GND_net), .I1(n8082[8]), .I2(GND_net), 
            .I3(n29749), .O(n8060[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_5 (.CI(n29554), .I0(n7845[2]), .I1(n311_adj_3787), 
            .CO(n29555));
    SB_LUT4 add_3695_4_lut (.I0(GND_net), .I1(n7845[1]), .I2(n238_adj_3789), 
            .I3(n29553), .O(n7826[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3714_11 (.CI(n29749), .I0(n8082[8]), .I1(GND_net), .CO(n29750));
    SB_LUT4 i34341_3_lut (.I0(n41918), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_3577), .I3(GND_net), .O(n41105));   // verilog/motorControl.v(39[38:63])
    defparam i34341_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3695_4 (.CI(n29553), .I0(n7845[1]), .I1(n238_adj_3789), 
            .CO(n29554));
    SB_LUT4 add_3695_3_lut (.I0(GND_net), .I1(n7845[0]), .I2(n165_adj_3790), 
            .I3(n29552), .O(n7826[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33995_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n42220), 
            .O(n40759));
    defparam i33995_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35429_4_lut (.I0(n41105), .I1(n41818), .I2(n45), .I3(n40757), 
            .O(n42193));   // verilog/motorControl.v(39[38:63])
    defparam i35429_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34349_3_lut (.I0(n42273), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41), .I3(GND_net), .O(n41113));   // verilog/motorControl.v(39[38:63])
    defparam i34349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n28172), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35431_4_lut (.I0(n41113), .I1(n42193), .I2(n45), .I3(n40759), 
            .O(n42195));   // verilog/motorControl.v(39[38:63])
    defparam i35431_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3714_10_lut (.I0(GND_net), .I1(n8082[7]), .I2(GND_net), 
            .I3(n29748), .O(n8060[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3695_3 (.CI(n29552), .I0(n7845[0]), .I1(n165_adj_3790), 
            .CO(n29553));
    SB_CARRY add_3714_10 (.CI(n29748), .I0(n8082[7]), .I1(GND_net), .CO(n29749));
    SB_LUT4 add_3695_2_lut (.I0(GND_net), .I1(n23_adj_3792), .I2(n92_adj_3793), 
            .I3(GND_net), .O(n7826[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3695_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n28172), .I0(GND_net), .I1(n1[17]), 
            .CO(n28173));
    SB_CARRY add_3695_2 (.CI(GND_net), .I0(n23_adj_3792), .I1(n92_adj_3793), 
            .CO(n29552));
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_3794));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_3694_19_lut (.I0(GND_net), .I1(n7826[16]), .I2(GND_net), 
            .I3(n29551), .O(n7806[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n28171), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3714_9_lut (.I0(GND_net), .I1(n8082[6]), .I2(GND_net), 
            .I3(n29747), .O(n8060[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3694_18_lut (.I0(GND_net), .I1(n7826[15]), .I2(GND_net), 
            .I3(n29550), .O(n7806[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3714_9 (.CI(n29747), .I0(n8082[6]), .I1(GND_net), .CO(n29748));
    SB_CARRY add_3694_18 (.CI(n29550), .I0(n7826[15]), .I1(GND_net), .CO(n29551));
    SB_LUT4 i35157_3_lut (.I0(n4_adj_3794), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n41921));   // verilog/motorControl.v(39[10:34])
    defparam i35157_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFE \PID_CONTROLLER.integral_1179__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[1]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 add_3714_8_lut (.I0(GND_net), .I1(n8082[5]), .I2(n521_adj_3796), 
            .I3(n29746), .O(n8060[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3694_17_lut (.I0(GND_net), .I1(n7826[14]), .I2(GND_net), 
            .I3(n29549), .O(n7806[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3714_8 (.CI(n29746), .I0(n8082[5]), .I1(n521_adj_3796), 
            .CO(n29747));
    SB_CARRY add_3694_17 (.CI(n29549), .I0(n7826[14]), .I1(GND_net), .CO(n29550));
    SB_DFFE \PID_CONTROLLER.integral_1179__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[2]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[3]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[4]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[5]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[6]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[7]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[8]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[9]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[10]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[11]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[12]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[13]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[14]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[15]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[16]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[17]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[18]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[19]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[20]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[21]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[22]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1179__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n28[23]));   // verilog/motorControl.v(40[21:33])
    SB_CARRY unary_minus_16_add_3_18 (.CI(n28171), .I0(GND_net), .I1(n1[16]), 
            .CO(n28172));
    SB_LUT4 add_3694_16_lut (.I0(GND_net), .I1(n7826[13]), .I2(GND_net), 
            .I3(n29548), .O(n7806[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35158_3_lut (.I0(n41921), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n41922));   // verilog/motorControl.v(39[10:34])
    defparam i35158_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n28170), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34137_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n44005), 
            .I2(IntegralLimit[16]), .I3(n41502), .O(n40901));
    defparam i34137_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_3694_16 (.CI(n29548), .I0(n7826[13]), .I1(GND_net), .CO(n29549));
    SB_CARRY unary_minus_16_add_3_17 (.CI(n28170), .I0(GND_net), .I1(n1[15]), 
            .CO(n28171));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n28169), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n28169), .I0(GND_net), .I1(n1[14]), 
            .CO(n28170));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n28168), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3714_7_lut (.I0(GND_net), .I1(n8082[4]), .I2(n448_adj_3800), 
            .I3(n29745), .O(n8060[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3694_15_lut (.I0(GND_net), .I1(n7826[12]), .I2(GND_net), 
            .I3(n29547), .O(n7806[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n28168), .I0(GND_net), .I1(n1[13]), 
            .CO(n28169));
    SB_CARRY add_3694_15 (.CI(n29547), .I0(n7826[12]), .I1(GND_net), .CO(n29548));
    SB_CARRY add_3714_7 (.CI(n29745), .I0(n8082[4]), .I1(n448_adj_3800), 
            .CO(n29746));
    SB_LUT4 i35383_4_lut (.I0(n30_adj_3772), .I1(n10_adj_3771), .I2(n44028), 
            .I3(n40899), .O(n42147));   // verilog/motorControl.v(39[10:34])
    defparam i35383_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3714_6_lut (.I0(GND_net), .I1(n8082[3]), .I2(n375_adj_3801), 
            .I3(n29744), .O(n8060[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3694_14_lut (.I0(GND_net), .I1(n7826[11]), .I2(GND_net), 
            .I3(n29546), .O(n7806[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34333_3_lut (.I0(n41922), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n41097));   // verilog/motorControl.v(39[10:34])
    defparam i34333_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3694_14 (.CI(n29546), .I0(n7826[11]), .I1(GND_net), .CO(n29547));
    SB_CARRY add_3714_6 (.CI(n29744), .I0(n8082[3]), .I1(n375_adj_3801), 
            .CO(n29745));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n28167), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35516_4_lut (.I0(n41097), .I1(n42147), .I2(n44028), .I3(n40901), 
            .O(n42280));   // verilog/motorControl.v(39[10:34])
    defparam i35516_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3694_13_lut (.I0(GND_net), .I1(n7826[10]), .I2(GND_net), 
            .I3(n29545), .O(n7806[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_13 (.CI(n29545), .I0(n7826[10]), .I1(GND_net), .CO(n29546));
    SB_LUT4 i35517_3_lut (.I0(n42280), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n42281));   // verilog/motorControl.v(39[10:34])
    defparam i35517_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3694_12_lut (.I0(GND_net), .I1(n7826[9]), .I2(GND_net), 
            .I3(n29544), .O(n7806[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3714_5_lut (.I0(GND_net), .I1(n8082[2]), .I2(n302_adj_3803), 
            .I3(n29743), .O(n8060[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3714_5 (.CI(n29743), .I0(n8082[2]), .I1(n302_adj_3803), 
            .CO(n29744));
    SB_CARRY add_3694_12 (.CI(n29544), .I0(n7826[9]), .I1(GND_net), .CO(n29545));
    SB_LUT4 i35513_3_lut (.I0(n42281), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n42277));   // verilog/motorControl.v(39[10:34])
    defparam i35513_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34120_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n43996), 
            .I2(IntegralLimit[21]), .I3(n42305), .O(n40884));
    defparam i34120_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_396_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n43994));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_396_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35425_4_lut (.I0(n41095), .I1(n41816), .I2(n43994), .I3(n40877), 
            .O(n42189));   // verilog/motorControl.v(39[10:34])
    defparam i35425_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34339_3_lut (.I0(n42277), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n41103));   // verilog/motorControl.v(39[10:34])
    defparam i34339_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35432_3_lut (.I0(n42195), .I1(\PID_CONTROLLER.integral_23__N_3454 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3453 ));   // verilog/motorControl.v(39[38:63])
    defparam i35432_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3714_4_lut (.I0(GND_net), .I1(n8082[1]), .I2(n229_adj_3804), 
            .I3(n29742), .O(n8060[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3694_11_lut (.I0(GND_net), .I1(n7826[8]), .I2(GND_net), 
            .I3(n29543), .O(n7806[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_11 (.CI(n29543), .I0(n7826[8]), .I1(GND_net), .CO(n29544));
    SB_LUT4 i35427_4_lut (.I0(n41103), .I1(n42189), .I2(n43994), .I3(n40884), 
            .O(n42191));   // verilog/motorControl.v(39[10:34])
    defparam i35427_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3694_10_lut (.I0(GND_net), .I1(n7826[7]), .I2(GND_net), 
            .I3(n29542), .O(n7806[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3714_4 (.CI(n29742), .I0(n8082[1]), .I1(n229_adj_3804), 
            .CO(n29743));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_838_4_lut  (.I0(n42191), .I1(\PID_CONTROLLER.integral_23__N_3453 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3451 ));   // verilog/motorControl.v(39[10:63])
    defparam \PID_CONTROLLER.integral_23__I_838_4_lut .LUT_INIT = 16'h80c8;
    SB_CARRY add_3694_10 (.CI(n29542), .I0(n7826[7]), .I1(GND_net), .CO(n29543));
    SB_LUT4 add_3714_3_lut (.I0(GND_net), .I1(n8082[0]), .I2(n156_adj_3805), 
            .I3(n29741), .O(n8060[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3694_9_lut (.I0(GND_net), .I1(n7826[6]), .I2(GND_net), 
            .I3(n29541), .O(n7806[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_9 (.CI(n29541), .I0(n7826[6]), .I1(GND_net), .CO(n29542));
    SB_CARRY add_3714_3 (.CI(n29741), .I0(n8082[0]), .I1(n156_adj_3805), 
            .CO(n29742));
    SB_LUT4 add_3714_2_lut (.I0(GND_net), .I1(n14_adj_3806), .I2(n83_adj_3807), 
            .I3(GND_net), .O(n8060[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3714_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3714_2 (.CI(GND_net), .I0(n14_adj_3806), .I1(n83_adj_3807), 
            .CO(n29741));
    SB_LUT4 add_3694_8_lut (.I0(GND_net), .I1(n7826[5]), .I2(n527_adj_3808), 
            .I3(n29540), .O(n7806[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n28167), .I0(GND_net), .I1(n1[12]), 
            .CO(n28168));
    SB_LUT4 add_3713_22_lut (.I0(GND_net), .I1(n8060[19]), .I2(GND_net), 
            .I3(n29740), .O(n8037[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_8 (.CI(n29540), .I0(n7826[5]), .I1(n527_adj_3808), 
            .CO(n29541));
    SB_LUT4 add_3694_7_lut (.I0(GND_net), .I1(n7826[4]), .I2(n454_adj_3809), 
            .I3(n29539), .O(n7806[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_21_lut (.I0(GND_net), .I1(n8060[18]), .I2(GND_net), 
            .I3(n29739), .O(n8037[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_7 (.CI(n29539), .I0(n7826[4]), .I1(n454_adj_3809), 
            .CO(n29540));
    SB_CARRY add_3713_21 (.CI(n29739), .I0(n8060[18]), .I1(GND_net), .CO(n29740));
    SB_LUT4 add_3694_6_lut (.I0(GND_net), .I1(n7826[3]), .I2(n381_adj_3810), 
            .I3(n29538), .O(n7806[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n28166), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_6 (.CI(n29538), .I0(n7826[3]), .I1(n381_adj_3810), 
            .CO(n29539));
    SB_LUT4 add_3713_20_lut (.I0(GND_net), .I1(n8060[17]), .I2(GND_net), 
            .I3(n29738), .O(n8037[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3713_20 (.CI(n29738), .I0(n8060[17]), .I1(GND_net), .CO(n29739));
    SB_LUT4 add_3694_5_lut (.I0(GND_net), .I1(n7826[2]), .I2(n308_adj_3812), 
            .I3(n29537), .O(n7806[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_19_lut (.I0(GND_net), .I1(n8060[16]), .I2(GND_net), 
            .I3(n29737), .O(n8037[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_5 (.CI(n29537), .I0(n7826[2]), .I1(n308_adj_3812), 
            .CO(n29538));
    SB_CARRY add_3713_19 (.CI(n29737), .I0(n8060[16]), .I1(GND_net), .CO(n29738));
    SB_LUT4 add_3694_4_lut (.I0(GND_net), .I1(n7826[1]), .I2(n235_adj_3813), 
            .I3(n29536), .O(n7806[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_4 (.CI(n29536), .I0(n7826[1]), .I1(n235_adj_3813), 
            .CO(n29537));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n28166), .I0(GND_net), .I1(n1[11]), 
            .CO(n28167));
    SB_LUT4 add_3713_18_lut (.I0(GND_net), .I1(n8060[15]), .I2(GND_net), 
            .I3(n29736), .O(n8037[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3694_3_lut (.I0(GND_net), .I1(n7826[0]), .I2(n162_adj_3814), 
            .I3(n29535), .O(n7806[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_3 (.CI(n29535), .I0(n7826[0]), .I1(n162_adj_3814), 
            .CO(n29536));
    SB_CARRY add_3713_18 (.CI(n29736), .I0(n8060[15]), .I1(GND_net), .CO(n29737));
    SB_LUT4 add_3694_2_lut (.I0(GND_net), .I1(n20_adj_3815), .I2(n89_adj_3816), 
            .I3(GND_net), .O(n7806[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3694_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3694_2 (.CI(GND_net), .I0(n20_adj_3815), .I1(n89_adj_3816), 
            .CO(n29535));
    SB_LUT4 add_3713_17_lut (.I0(GND_net), .I1(n8060[14]), .I2(GND_net), 
            .I3(n29735), .O(n8037[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3693_20_lut (.I0(GND_net), .I1(n7806[17]), .I2(GND_net), 
            .I3(n29534), .O(n7785[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3693_19_lut (.I0(GND_net), .I1(n7806[16]), .I2(GND_net), 
            .I3(n29533), .O(n7785[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_636_25_lut (.I0(GND_net), .I1(n2996[23]), .I2(n3021[23]), 
            .I3(n28022), .O(duty_23__N_3478[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_19 (.CI(n29533), .I0(n7806[16]), .I1(GND_net), .CO(n29534));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n28165), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3713_17 (.CI(n29735), .I0(n8060[14]), .I1(GND_net), .CO(n29736));
    SB_LUT4 add_3693_18_lut (.I0(GND_net), .I1(n7806[15]), .I2(GND_net), 
            .I3(n29532), .O(n7785[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_18 (.CI(n29532), .I0(n7806[15]), .I1(GND_net), .CO(n29533));
    SB_CARRY unary_minus_16_add_3_12 (.CI(n28165), .I0(GND_net), .I1(n1[10]), 
            .CO(n28166));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n28164), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_16_lut (.I0(GND_net), .I1(n8060[13]), .I2(GND_net), 
            .I3(n29734), .O(n8037[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3693_17_lut (.I0(GND_net), .I1(n7806[14]), .I2(GND_net), 
            .I3(n29531), .O(n7785[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_17 (.CI(n29531), .I0(n7806[14]), .I1(GND_net), .CO(n29532));
    SB_CARRY add_3713_16 (.CI(n29734), .I0(n8060[13]), .I1(GND_net), .CO(n29735));
    SB_LUT4 add_3693_16_lut (.I0(GND_net), .I1(n7806[13]), .I2(GND_net), 
            .I3(n29530), .O(n7785[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_16 (.CI(n29530), .I0(n7806[13]), .I1(GND_net), .CO(n29531));
    SB_LUT4 add_3713_15_lut (.I0(GND_net), .I1(n8060[12]), .I2(GND_net), 
            .I3(n29733), .O(n8037[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3693_15_lut (.I0(GND_net), .I1(n7806[12]), .I2(GND_net), 
            .I3(n29529), .O(n7785[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_15 (.CI(n29529), .I0(n7806[12]), .I1(GND_net), .CO(n29530));
    SB_CARRY add_3713_15 (.CI(n29733), .I0(n8060[12]), .I1(GND_net), .CO(n29734));
    SB_LUT4 add_3713_14_lut (.I0(GND_net), .I1(n8060[11]), .I2(GND_net), 
            .I3(n29732), .O(n8037[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3693_14_lut (.I0(GND_net), .I1(n7806[11]), .I2(GND_net), 
            .I3(n29528), .O(n7785[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_14 (.CI(n29528), .I0(n7806[11]), .I1(GND_net), .CO(n29529));
    SB_CARRY add_3713_14 (.CI(n29732), .I0(n8060[11]), .I1(GND_net), .CO(n29733));
    SB_LUT4 add_3693_13_lut (.I0(GND_net), .I1(n7806[10]), .I2(GND_net), 
            .I3(n29527), .O(n7785[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_13 (.CI(n29527), .I0(n7806[10]), .I1(GND_net), .CO(n29528));
    SB_LUT4 add_3693_12_lut (.I0(GND_net), .I1(n7806[9]), .I2(GND_net), 
            .I3(n29526), .O(n7785[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_13_lut (.I0(GND_net), .I1(n8060[10]), .I2(GND_net), 
            .I3(n29731), .O(n8037[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_12 (.CI(n29526), .I0(n7806[9]), .I1(GND_net), .CO(n29527));
    SB_LUT4 add_3693_11_lut (.I0(GND_net), .I1(n7806[8]), .I2(GND_net), 
            .I3(n29525), .O(n7785[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_11 (.CI(n29525), .I0(n7806[8]), .I1(GND_net), .CO(n29526));
    SB_CARRY add_3713_13 (.CI(n29731), .I0(n8060[10]), .I1(GND_net), .CO(n29732));
    SB_LUT4 add_3693_10_lut (.I0(GND_net), .I1(n7806[7]), .I2(GND_net), 
            .I3(n29524), .O(n7785[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_10 (.CI(n29524), .I0(n7806[7]), .I1(GND_net), .CO(n29525));
    SB_LUT4 add_636_24_lut (.I0(GND_net), .I1(n2996[22]), .I2(n3021[22]), 
            .I3(n28021), .O(duty_23__N_3478[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_12_lut (.I0(GND_net), .I1(n8060[9]), .I2(GND_net), 
            .I3(n29730), .O(n8037[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3693_9_lut (.I0(GND_net), .I1(n7806[6]), .I2(GND_net), 
            .I3(n29523), .O(n7785[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_9 (.CI(n29523), .I0(n7806[6]), .I1(GND_net), .CO(n29524));
    SB_CARRY add_3713_12 (.CI(n29730), .I0(n8060[9]), .I1(GND_net), .CO(n29731));
    SB_LUT4 add_3693_8_lut (.I0(GND_net), .I1(n7806[5]), .I2(n524_adj_3819), 
            .I3(n29522), .O(n7785[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_11_lut (.I0(GND_net), .I1(n8060[8]), .I2(GND_net), 
            .I3(n29729), .O(n8037[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_8 (.CI(n29522), .I0(n7806[5]), .I1(n524_adj_3819), 
            .CO(n29523));
    SB_LUT4 add_3693_7_lut (.I0(GND_net), .I1(n7806[4]), .I2(n451_adj_3820), 
            .I3(n29521), .O(n7785[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_24 (.CI(n28021), .I0(n2996[22]), .I1(n3021[22]), 
            .CO(n28022));
    SB_CARRY unary_minus_16_add_3_11 (.CI(n28164), .I0(GND_net), .I1(n1[9]), 
            .CO(n28165));
    SB_LUT4 add_636_23_lut (.I0(GND_net), .I1(n2996[21]), .I2(n3021[21]), 
            .I3(n28020), .O(duty_23__N_3478[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_23 (.CI(n28020), .I0(n2996[21]), .I1(n3021[21]), 
            .CO(n28021));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n28163), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n28163), .I0(GND_net), .I1(n1[8]), 
            .CO(n28164));
    SB_CARRY add_3693_7 (.CI(n29521), .I0(n7806[4]), .I1(n451_adj_3820), 
            .CO(n29522));
    SB_CARRY add_3713_11 (.CI(n29729), .I0(n8060[8]), .I1(GND_net), .CO(n29730));
    SB_LUT4 add_3693_6_lut (.I0(GND_net), .I1(n7806[3]), .I2(n378_adj_3822), 
            .I3(n29520), .O(n7785[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_10_lut (.I0(GND_net), .I1(n8060[7]), .I2(GND_net), 
            .I3(n29728), .O(n8037[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_6 (.CI(n29520), .I0(n7806[3]), .I1(n378_adj_3822), 
            .CO(n29521));
    SB_CARRY add_3713_10 (.CI(n29728), .I0(n8060[7]), .I1(GND_net), .CO(n29729));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n28162), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3693_5_lut (.I0(GND_net), .I1(n7806[2]), .I2(n305_adj_3824), 
            .I3(n29519), .O(n7785[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_5 (.CI(n29519), .I0(n7806[2]), .I1(n305_adj_3824), 
            .CO(n29520));
    SB_LUT4 add_3693_4_lut (.I0(GND_net), .I1(n7806[1]), .I2(n232_adj_3825), 
            .I3(n29518), .O(n7785[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_9_lut (.I0(GND_net), .I1(n8060[6]), .I2(GND_net), 
            .I3(n29727), .O(n8037[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_4 (.CI(n29518), .I0(n7806[1]), .I1(n232_adj_3825), 
            .CO(n29519));
    SB_LUT4 add_3693_3_lut (.I0(GND_net), .I1(n7806[0]), .I2(n159_adj_3826), 
            .I3(n29517), .O(n7785[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_3 (.CI(n29517), .I0(n7806[0]), .I1(n159_adj_3826), 
            .CO(n29518));
    SB_LUT4 add_636_22_lut (.I0(GND_net), .I1(n2996[20]), .I2(n3021[20]), 
            .I3(n28019), .O(duty_23__N_3478[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n28162), .I0(GND_net), .I1(n1[7]), 
            .CO(n28163));
    SB_CARRY add_3713_9 (.CI(n29727), .I0(n8060[6]), .I1(GND_net), .CO(n29728));
    SB_LUT4 add_3693_2_lut (.I0(GND_net), .I1(n17_adj_3827), .I2(n86_adj_3828), 
            .I3(GND_net), .O(n7785[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3693_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3693_2 (.CI(GND_net), .I0(n17_adj_3827), .I1(n86_adj_3828), 
            .CO(n29517));
    SB_LUT4 add_3713_8_lut (.I0(GND_net), .I1(n8060[5]), .I2(n518_adj_3829), 
            .I3(n29726), .O(n8037[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_21_lut (.I0(GND_net), .I1(n7785[18]), .I2(GND_net), 
            .I3(n29516), .O(n7763[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n28161), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_20_lut (.I0(GND_net), .I1(n7785[17]), .I2(GND_net), 
            .I3(n29515), .O(n7763[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3713_8 (.CI(n29726), .I0(n8060[5]), .I1(n518_adj_3829), 
            .CO(n29727));
    SB_CARRY add_3692_20 (.CI(n29515), .I0(n7785[17]), .I1(GND_net), .CO(n29516));
    SB_LUT4 add_3713_7_lut (.I0(GND_net), .I1(n8060[4]), .I2(n445_adj_3831), 
            .I3(n29725), .O(n8037[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_19_lut (.I0(GND_net), .I1(n7785[16]), .I2(GND_net), 
            .I3(n29514), .O(n7763[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3713_7 (.CI(n29725), .I0(n8060[4]), .I1(n445_adj_3831), 
            .CO(n29726));
    SB_LUT4 mux_634_i24_3_lut_3_lut (.I0(PWMLimit[23]), .I1(n256_adj_3571), 
            .I2(n40149), .I3(GND_net), .O(n3021[23]));   // verilog/motorControl.v(47[19:28])
    defparam mux_634_i24_3_lut_3_lut.LUT_INIT = 16'h7474;
    SB_CARRY add_3692_19 (.CI(n29514), .I0(n7785[16]), .I1(GND_net), .CO(n29515));
    SB_LUT4 add_3692_18_lut (.I0(GND_net), .I1(n7785[15]), .I2(GND_net), 
            .I3(n29513), .O(n7763[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n28161), .I0(GND_net), .I1(n1[6]), 
            .CO(n28162));
    SB_LUT4 add_3713_6_lut (.I0(GND_net), .I1(n8060[3]), .I2(n372_adj_3832), 
            .I3(n29724), .O(n8037[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_18 (.CI(n29513), .I0(n7785[15]), .I1(GND_net), .CO(n29514));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n28160), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n28160), .I0(GND_net), .I1(n1[5]), 
            .CO(n28161));
    SB_LUT4 add_3692_17_lut (.I0(GND_net), .I1(n7785[14]), .I2(GND_net), 
            .I3(n29512), .O(n7763[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_22 (.CI(n28019), .I0(n2996[20]), .I1(n3021[20]), 
            .CO(n28020));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n28159), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_636_21_lut (.I0(GND_net), .I1(n2996[19]), .I2(n3021[19]), 
            .I3(n28018), .O(duty_23__N_3478[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n28159), .I0(GND_net), .I1(n1[4]), 
            .CO(n28160));
    SB_CARRY add_3713_6 (.CI(n29724), .I0(n8060[3]), .I1(n372_adj_3832), 
            .CO(n29725));
    SB_LUT4 add_3713_5_lut (.I0(GND_net), .I1(n8060[2]), .I2(n299_adj_3835), 
            .I3(n29723), .O(n8037[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_17 (.CI(n29512), .I0(n7785[14]), .I1(GND_net), .CO(n29513));
    SB_LUT4 add_3692_16_lut (.I0(GND_net), .I1(n7785[13]), .I2(GND_net), 
            .I3(n29511), .O(n7763[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n28158), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_16 (.CI(n29511), .I0(n7785[13]), .I1(GND_net), .CO(n29512));
    SB_CARRY unary_minus_16_add_3_5 (.CI(n28158), .I0(GND_net), .I1(n1[3]), 
            .CO(n28159));
    SB_CARRY add_636_21 (.CI(n28018), .I0(n2996[19]), .I1(n3021[19]), 
            .CO(n28019));
    SB_LUT4 add_636_20_lut (.I0(GND_net), .I1(n2996[18]), .I2(n3021[18]), 
            .I3(n28017), .O(duty_23__N_3478[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3713_5 (.CI(n29723), .I0(n8060[2]), .I1(n299_adj_3835), 
            .CO(n29724));
    SB_LUT4 add_3692_15_lut (.I0(GND_net), .I1(n7785[12]), .I2(GND_net), 
            .I3(n29510), .O(n7763[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n28157), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n28157), .I0(GND_net), .I1(n1[2]), 
            .CO(n28158));
    SB_LUT4 add_3713_4_lut (.I0(GND_net), .I1(n8060[1]), .I2(n226_adj_3838), 
            .I3(n29722), .O(n8037[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_15 (.CI(n29510), .I0(n7785[12]), .I1(GND_net), .CO(n29511));
    SB_LUT4 add_3692_14_lut (.I0(GND_net), .I1(n7785[11]), .I2(GND_net), 
            .I3(n29509), .O(n7763[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_7_lut (.I0(GND_net), .I1(n36243), .I2(n490_adj_3839), 
            .I3(n29920), .O(n8277[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3728_6_lut (.I0(GND_net), .I1(n8285[3]), .I2(n417_adj_3840), 
            .I3(n29919), .O(n8277[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_6 (.CI(n29919), .I0(n8285[3]), .I1(n417_adj_3840), 
            .CO(n29920));
    SB_LUT4 add_3728_5_lut (.I0(GND_net), .I1(n8285[2]), .I2(n344_adj_3841), 
            .I3(n29918), .O(n8277[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_5 (.CI(n29918), .I0(n8285[2]), .I1(n344_adj_3841), 
            .CO(n29919));
    SB_CARRY add_3713_4 (.CI(n29722), .I0(n8060[1]), .I1(n226_adj_3838), 
            .CO(n29723));
    SB_LUT4 add_3728_4_lut (.I0(GND_net), .I1(n8285[1]), .I2(n271_adj_3842), 
            .I3(n29917), .O(n8277[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_4 (.CI(n29917), .I0(n8285[1]), .I1(n271_adj_3842), 
            .CO(n29918));
    SB_LUT4 add_3728_3_lut (.I0(GND_net), .I1(n8285[0]), .I2(n198_adj_3843), 
            .I3(n29916), .O(n8277[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_3 (.CI(n29916), .I0(n8285[0]), .I1(n198_adj_3843), 
            .CO(n29917));
    SB_LUT4 add_3728_2_lut (.I0(GND_net), .I1(n56_adj_3844), .I2(n125_adj_3845), 
            .I3(GND_net), .O(n8277[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3728_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3728_2 (.CI(GND_net), .I0(n56_adj_3844), .I1(n125_adj_3845), 
            .CO(n29916));
    SB_LUT4 add_3727_8_lut (.I0(GND_net), .I1(n8277[5]), .I2(n560_adj_3846), 
            .I3(n29915), .O(n8268[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3727_7_lut (.I0(GND_net), .I1(n8277[4]), .I2(n487_adj_3847), 
            .I3(n29914), .O(n8268[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_7 (.CI(n29914), .I0(n8277[4]), .I1(n487_adj_3847), 
            .CO(n29915));
    SB_LUT4 add_3727_6_lut (.I0(GND_net), .I1(n8277[3]), .I2(n414_adj_3848), 
            .I3(n29913), .O(n8268[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_14 (.CI(n29509), .I0(n7785[11]), .I1(GND_net), .CO(n29510));
    SB_CARRY add_3727_6 (.CI(n29913), .I0(n8277[3]), .I1(n414_adj_3848), 
            .CO(n29914));
    SB_LUT4 add_3727_5_lut (.I0(GND_net), .I1(n8277[2]), .I2(n341_adj_3849), 
            .I3(n29912), .O(n8268[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_20 (.CI(n28017), .I0(n2996[18]), .I1(n3021[18]), 
            .CO(n28018));
    SB_LUT4 add_3692_13_lut (.I0(GND_net), .I1(n7785[10]), .I2(GND_net), 
            .I3(n29508), .O(n7763[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_5 (.CI(n29912), .I0(n8277[2]), .I1(n341_adj_3849), 
            .CO(n29913));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n28156), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3727_4_lut (.I0(GND_net), .I1(n8277[1]), .I2(n268_adj_3851), 
            .I3(n29911), .O(n8268[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_4 (.CI(n29911), .I0(n8277[1]), .I1(n268_adj_3851), 
            .CO(n29912));
    SB_LUT4 add_3727_3_lut (.I0(GND_net), .I1(n8277[0]), .I2(n195_adj_3852), 
            .I3(n29910), .O(n8268[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_3 (.CI(n29910), .I0(n8277[0]), .I1(n195_adj_3852), 
            .CO(n29911));
    SB_LUT4 add_3727_2_lut (.I0(GND_net), .I1(n53_adj_3853), .I2(n122_adj_3854), 
            .I3(GND_net), .O(n8268[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3727_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3727_2 (.CI(GND_net), .I0(n53_adj_3853), .I1(n122_adj_3854), 
            .CO(n29910));
    SB_LUT4 add_3726_9_lut (.I0(GND_net), .I1(n8268[6]), .I2(GND_net), 
            .I3(n29909), .O(n8258[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3726_8_lut (.I0(GND_net), .I1(n8268[5]), .I2(n557_adj_3855), 
            .I3(n29908), .O(n8258[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_3_lut (.I0(GND_net), .I1(n8060[0]), .I2(n153_adj_3856), 
            .I3(n29721), .O(n8037[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_8 (.CI(n29908), .I0(n8268[5]), .I1(n557_adj_3855), 
            .CO(n29909));
    SB_LUT4 add_3726_7_lut (.I0(GND_net), .I1(n8268[4]), .I2(n484_adj_3857), 
            .I3(n29907), .O(n8258[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_7 (.CI(n29907), .I0(n8268[4]), .I1(n484_adj_3857), 
            .CO(n29908));
    SB_LUT4 add_3726_6_lut (.I0(GND_net), .I1(n8268[3]), .I2(n411_adj_3858), 
            .I3(n29906), .O(n8258[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3692_13 (.CI(n29508), .I0(n7785[10]), .I1(GND_net), .CO(n29509));
    SB_CARRY add_3726_6 (.CI(n29906), .I0(n8268[3]), .I1(n411_adj_3858), 
            .CO(n29907));
    SB_LUT4 add_3726_5_lut (.I0(GND_net), .I1(n8268[2]), .I2(n338_adj_3859), 
            .I3(n29905), .O(n8258[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_5 (.CI(n29905), .I0(n8268[2]), .I1(n338_adj_3859), 
            .CO(n29906));
    SB_LUT4 add_3726_4_lut (.I0(GND_net), .I1(n8268[1]), .I2(n265_adj_3860), 
            .I3(n29904), .O(n8258[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_12_lut (.I0(GND_net), .I1(n7785[9]), .I2(GND_net), 
            .I3(n29507), .O(n7763[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_4 (.CI(n29904), .I0(n8268[1]), .I1(n265_adj_3860), 
            .CO(n29905));
    SB_LUT4 add_3726_3_lut (.I0(GND_net), .I1(n8268[0]), .I2(n192_adj_3861), 
            .I3(n29903), .O(n8258[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_3 (.CI(n29903), .I0(n8268[0]), .I1(n192_adj_3861), 
            .CO(n29904));
    SB_LUT4 add_3726_2_lut (.I0(GND_net), .I1(n50_adj_3862), .I2(n119_adj_3863), 
            .I3(GND_net), .O(n8258[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3726_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3726_2 (.CI(GND_net), .I0(n50_adj_3862), .I1(n119_adj_3863), 
            .CO(n29903));
    SB_LUT4 add_3725_10_lut (.I0(GND_net), .I1(n8258[7]), .I2(GND_net), 
            .I3(n29902), .O(n8247[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3725_9_lut (.I0(GND_net), .I1(n8258[6]), .I2(GND_net), 
            .I3(n29901), .O(n8247[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_9 (.CI(n29901), .I0(n8258[6]), .I1(GND_net), .CO(n29902));
    SB_LUT4 add_3725_8_lut (.I0(GND_net), .I1(n8258[5]), .I2(n554_adj_3864), 
            .I3(n29900), .O(n8247[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_8 (.CI(n29900), .I0(n8258[5]), .I1(n554_adj_3864), 
            .CO(n29901));
    SB_LUT4 add_3725_7_lut (.I0(GND_net), .I1(n8258[4]), .I2(n481_adj_3865), 
            .I3(n29899), .O(n8247[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_7 (.CI(n29899), .I0(n8258[4]), .I1(n481_adj_3865), 
            .CO(n29900));
    SB_LUT4 add_3725_6_lut (.I0(GND_net), .I1(n8258[3]), .I2(n408_adj_3866), 
            .I3(n29898), .O(n8247[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_6 (.CI(n29898), .I0(n8258[3]), .I1(n408_adj_3866), 
            .CO(n29899));
    SB_LUT4 add_3725_5_lut (.I0(GND_net), .I1(n8258[2]), .I2(n335_adj_3867), 
            .I3(n29897), .O(n8247[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_5 (.CI(n29897), .I0(n8258[2]), .I1(n335_adj_3867), 
            .CO(n29898));
    SB_LUT4 add_636_19_lut (.I0(GND_net), .I1(n2996[17]), .I2(n3021[17]), 
            .I3(n28016), .O(duty_23__N_3478[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3725_4_lut (.I0(GND_net), .I1(n8258[1]), .I2(n262_adj_3868), 
            .I3(n29896), .O(n8247[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_4 (.CI(n29896), .I0(n8258[1]), .I1(n262_adj_3868), 
            .CO(n29897));
    SB_CARRY add_3713_3 (.CI(n29721), .I0(n8060[0]), .I1(n153_adj_3856), 
            .CO(n29722));
    SB_LUT4 add_3725_3_lut (.I0(GND_net), .I1(n8258[0]), .I2(n189_adj_3869), 
            .I3(n29895), .O(n8247[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_3 (.CI(n29895), .I0(n8258[0]), .I1(n189_adj_3869), 
            .CO(n29896));
    SB_CARRY add_3692_12 (.CI(n29507), .I0(n7785[9]), .I1(GND_net), .CO(n29508));
    SB_LUT4 add_3725_2_lut (.I0(GND_net), .I1(n47_adj_3870), .I2(n116_adj_3871), 
            .I3(GND_net), .O(n8247[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3725_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3725_2 (.CI(GND_net), .I0(n47_adj_3870), .I1(n116_adj_3871), 
            .CO(n29895));
    SB_LUT4 add_3724_11_lut (.I0(GND_net), .I1(n8247[8]), .I2(GND_net), 
            .I3(n29894), .O(n8235[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_11_lut (.I0(GND_net), .I1(n7785[8]), .I2(GND_net), 
            .I3(n29506), .O(n7763[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3724_10_lut (.I0(GND_net), .I1(n8247[7]), .I2(GND_net), 
            .I3(n29893), .O(n8235[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_636_19 (.CI(n28016), .I0(n2996[17]), .I1(n3021[17]), 
            .CO(n28017));
    SB_CARRY add_3692_11 (.CI(n29506), .I0(n7785[8]), .I1(GND_net), .CO(n29507));
    SB_CARRY add_3724_10 (.CI(n29893), .I0(n8247[7]), .I1(GND_net), .CO(n29894));
    SB_LUT4 add_3724_9_lut (.I0(GND_net), .I1(n8247[6]), .I2(GND_net), 
            .I3(n29892), .O(n8235[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_9 (.CI(n29892), .I0(n8247[6]), .I1(GND_net), .CO(n29893));
    SB_LUT4 add_3724_8_lut (.I0(GND_net), .I1(n8247[5]), .I2(n551_adj_3872), 
            .I3(n29891), .O(n8235[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_8 (.CI(n29891), .I0(n8247[5]), .I1(n551_adj_3872), 
            .CO(n29892));
    SB_LUT4 add_3724_7_lut (.I0(GND_net), .I1(n8247[4]), .I2(n478_adj_3873), 
            .I3(n29890), .O(n8235[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_7 (.CI(n29890), .I0(n8247[4]), .I1(n478_adj_3873), 
            .CO(n29891));
    SB_LUT4 add_3724_6_lut (.I0(GND_net), .I1(n8247[3]), .I2(n405_adj_3874), 
            .I3(n29889), .O(n8235[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3724_6 (.CI(n29889), .I0(n8247[3]), .I1(n405_adj_3874), 
            .CO(n29890));
    SB_LUT4 add_636_18_lut (.I0(GND_net), .I1(n2996[16]), .I2(n3021[16]), 
            .I3(n28015), .O(duty_23__N_3478[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_636_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n28156), .I0(GND_net), .I1(n1[1]), 
            .CO(n28157));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n40103)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3724_5_lut (.I0(GND_net), .I1(n8247[2]), .I2(n332_adj_3876), 
            .I3(n29888), .O(n8235[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3713_2_lut (.I0(GND_net), .I1(n11_adj_3877), .I2(n80_adj_3878), 
            .I3(GND_net), .O(n8037[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3713_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_10_lut (.I0(GND_net), .I1(n7785[7]), .I2(GND_net), 
            .I3(n29505), .O(n7763[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3713_2 (.CI(GND_net), .I0(n11_adj_3877), .I1(n80_adj_3878), 
            .CO(n29721));
    SB_CARRY add_3724_5 (.CI(n29888), .I0(n8247[2]), .I1(n332_adj_3876), 
            .CO(n29889));
    SB_CARRY add_3692_10 (.CI(n29505), .I0(n7785[7]), .I1(GND_net), .CO(n29506));
    SB_LUT4 add_3724_4_lut (.I0(GND_net), .I1(n8247[1]), .I2(n259_adj_3879), 
            .I3(n29887), .O(n8235[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3724_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n8013[21]), 
            .I2(GND_net), .I3(n29720), .O(n40149)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3724_4 (.CI(n29887), .I0(n8247[1]), .I1(n259_adj_3879), 
            .CO(n29888));
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n8013[20]), .I2(GND_net), 
            .I3(n29719), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3692_9_lut (.I0(GND_net), .I1(n7785[6]), .I2(GND_net), 
            .I3(n29504), .O(n7763[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3692_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3685));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_3683));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23065_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n27655), .I3(n8006[0]), .O(n4_adj_3569));   // verilog/motorControl.v(42[17:23])
    defparam i23065_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n8006[0]), .I3(n27655), .O(n8001[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_845 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n8001[0]), .I3(n27621), .O(n7995[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_845.LUT_INIT = 16'h8778;
    SB_LUT4 i23034_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n27621), .I3(n8001[0]), .O(n4_adj_3565));   // verilog/motorControl.v(42[17:23])
    defparam i23034_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i23054_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n27655));   // verilog/motorControl.v(42[17:23])
    defparam i23054_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i23052_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n8001[0]));   // verilog/motorControl.v(42[17:23])
    defparam i23052_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i19581_2_lut_2_lut (.I0(n256_adj_3571), .I1(n6169[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2996[23]));   // verilog/motorControl.v(46[19:35])
    defparam i19581_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19317_3_lut (.I0(\Kp[0] ), .I1(n256_adj_3571), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n2996[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam i19317_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3667));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3666));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_3665));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23163_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_3880), .I3(n8292[1]), .O(n6_adj_3881));   // verilog/motorControl.v(42[26:37])
    defparam i23163_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_3664));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i2_3_lut (.I0(n155[1]), .I1(PWMLimit[1]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_3663));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_3662));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_3660));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_3659));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3656));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3655));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_846 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8292[1]), .I3(n4_adj_3880), .O(n8285[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_846.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_847 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n8298[0]), .I3(n27791), .O(n8292[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_847.LUT_INIT = 16'h8778;
    SB_LUT4 i23194_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n27791), .I3(n8298[0]), .O(n4_adj_3882));   // verilog/motorControl.v(42[26:37])
    defparam i23194_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3654));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3653));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_3652));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_3650));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_3648));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3647));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23181_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(\Ki[1] ), .O(n8292[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23181_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3646));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_3645));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3644));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_3643));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_3642));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3879));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_3878));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23183_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(\Ki[1] ), .O(n27791));   // verilog/motorControl.v(42[26:37])
    defparam i23183_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3877));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_3876));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_3874));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_3873));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_3872));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3871));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3870));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3869));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3868));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i18_3_lut (.I0(n155[17]), .I1(n1[17]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_3867));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_3866));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_3865));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_3864));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3863));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3862));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3861));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3860));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_3859));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_3858));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_3857));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_3856));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_3855));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_3641));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3854));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3853));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_3640));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_3639));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3638));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3637));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36317_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43079));   // verilog/motorControl.v(37[14] 56[8])
    defparam i36317_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[0]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3635));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[1]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3852));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i4_3_lut (.I0(n155[3]), .I1(PWMLimit[3]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i4_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3631));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3851));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23225_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n27825), .I3(n8303[0]), .O(n4_adj_3883));   // verilog/motorControl.v(42[26:37])
    defparam i23225_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_848 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n8303[0]), .I3(n27825), .O(n8298[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_848.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_3849));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_3848));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3630));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_3847));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_3846));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3845));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_3844));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3843));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3842));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_3841));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23212_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n8298[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23212_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_3840));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_849 (.I0(n6_adj_3881), .I1(\Ki[4] ), .I2(n8292[2]), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8285[3]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_849.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23235_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n8303[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23235_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_850 (.I0(n4_adj_3882), .I1(\Ki[3] ), .I2(n8298[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n8292[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_850.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_3839));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_851 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_3884));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_851.LUT_INIT = 16'h9c50;
    SB_LUT4 i23214_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n27825));   // verilog/motorControl.v(42[26:37])
    defparam i23214_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i23171_4_lut (.I0(n8292[2]), .I1(\Ki[4] ), .I2(n6_adj_3881), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_3885));   // verilog/motorControl.v(42[26:37])
    defparam i23171_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_852 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8292[0]), .I3(n27748), .O(n8285[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_852.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_853 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_3886));   // verilog/motorControl.v(42[26:37])
    defparam i1_4_lut_adj_853.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23202_4_lut (.I0(n8298[1]), .I1(\Ki[3] ), .I2(n4_adj_3882), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_3887));   // verilog/motorControl.v(42[26:37])
    defparam i23202_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i23237_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n27850));   // verilog/motorControl.v(42[26:37])
    defparam i23237_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_854 (.I0(n6_adj_3887), .I1(n11_adj_3886), .I2(n8_adj_3885), 
            .I3(n12_adj_3884), .O(n18_adj_3888));   // verilog/motorControl.v(42[26:37])
    defparam i8_4_lut_adj_854.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_855 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_3889));   // verilog/motorControl.v(42[26:37])
    defparam i3_4_lut_adj_855.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[2]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut_adj_856 (.I0(n13_adj_3889), .I1(n18_adj_3888), .I2(n27850), 
            .I3(n4_adj_3883), .O(n36243));   // verilog/motorControl.v(42[26:37])
    defparam i9_4_lut_adj_856.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_3627));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3626));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[3]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_3624));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_3838));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23155_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n27748), .I3(n8292[0]), .O(n4_adj_3880));   // verilog/motorControl.v(42[26:37])
    defparam i23155_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_3623));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3622));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3621));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_3620));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_3619));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_3618));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i5_3_lut (.I0(n155[4]), .I1(PWMLimit[4]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i5_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[4]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_3615));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23142_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n8285[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23142_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mux_634_i6_3_lut (.I0(n155[5]), .I1(PWMLimit[5]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i6_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mux_634_i19_3_lut (.I0(n155[18]), .I1(n1[18]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[5]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_3835));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i20_3_lut (.I0(n155[19]), .I1(n1[19]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_634_i7_3_lut (.I0(n155[6]), .I1(PWMLimit[6]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i7_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i23144_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n27748));   // verilog/motorControl.v(42[26:37])
    defparam i23144_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3612));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_3832));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_3831));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_3829));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3828));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3827));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i21_3_lut (.I0(n155[20]), .I1(n1[20]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3610));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3609));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3608));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_3607));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[6]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[7]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_3826));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_3825));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3602));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3601));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_3600));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_3599));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i8_3_lut (.I0(n155[7]), .I1(PWMLimit[7]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i8_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3891[8]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_3824));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_3822));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_3596));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_3595));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_3592));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3589));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_857 (.I0(n6_adj_3566), .I1(\Kp[4] ), .I2(n7995[2]), 
            .I3(\PID_CONTROLLER.err [18]), .O(n7988[3]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_857.LUT_INIT = 16'h965a;
    SB_LUT4 i23075_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n8006[0]));   // verilog/motorControl.v(42[17:23])
    defparam i23075_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_634_i22_3_lut (.I0(n155[21]), .I1(n1[21]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_3820));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_3819));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_634_i23_3_lut (.I0(n155[22]), .I1(n1[22]), .I2(n256_adj_3571), 
            .I3(GND_net), .O(n3021[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_3816));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3815));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_3814));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_3813));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_3812));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_3810));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_3809));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_3808));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_3807));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3806));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_3805));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_3804));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_3803));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_3801));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_3800));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_3796));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_3793));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3792));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_3790));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_3789));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_3787));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_3786));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_3785));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_3783));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_3763));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3762));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3761));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3760));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3759));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_3758));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_3757));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_3755));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3754));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[0]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[1]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[2]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3892[3]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33859_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n40623));   // verilog/motorControl.v(46[19:35])
    defparam i33859_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_3729));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i23003_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_3890), .I3(n7995[1]), .O(n6_adj_3566));   // verilog/motorControl.v(42[17:23])
    defparam i23003_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_858 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n7995[1]), .I3(n4_adj_3890), .O(n7988[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_858.LUT_INIT = 16'h8778;
    SB_LUT4 mux_634_i1_4_lut_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256_adj_3571), .I3(\Ki[0] ), .O(n3021[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_634_i1_4_lut_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3776));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut_4_lut_adj_859 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n7995[0]), .I3(n27578), .O(n7988[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_859.LUT_INIT = 16'h8778;
    SB_LUT4 i33691_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n40453));
    defparam i33691_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i33747_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n40509));
    defparam i33747_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i22995_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n27578), .I3(n7995[0]), .O(n4_adj_3890));   // verilog/motorControl.v(42[17:23])
    defparam i22995_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 duty_23__I_0_i4_4_lut_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_3695));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i4_4_lut_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_3694));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33863_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n40627));
    defparam i33863_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16_adj_3692));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_3698));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33919_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n40683));
    defparam i33919_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12_adj_3686));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33985_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n40749));   // verilog/motorControl.v(44[10:25])
    defparam i33985_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_3691));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i22982_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n7988[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22982_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22984_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n27578));   // verilog/motorControl.v(42[17:23])
    defparam i22984_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (PIN_19_c_0, CLK_c, \half_duty_new[0] , 
            n17573, \half_duty[0][7] , n17567, \half_duty[0][1] , n17568, 
            \half_duty[0][2] , n17569, \half_duty[0][3] , n17570, \half_duty[0][4] , 
            n17572, \half_duty[0][6] , n1169, GND_net, VCC_net, \half_duty_new[1] , 
            \half_duty[0][0] , \half_duty_new[2] , \half_duty_new[3] , 
            \half_duty_new[4] , \half_duty_new[6] , \half_duty_new[7] , 
            n16982, pwm_setpoint) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    output PIN_19_c_0;
    input CLK_c;
    output \half_duty_new[0] ;
    input n17573;
    output \half_duty[0][7] ;
    input n17567;
    output \half_duty[0][1] ;
    input n17568;
    output \half_duty[0][2] ;
    input n17569;
    output \half_duty[0][3] ;
    input n17570;
    output \half_duty[0][4] ;
    input n17572;
    output \half_duty[0][6] ;
    output n1169;
    input GND_net;
    input VCC_net;
    output \half_duty_new[1] ;
    output \half_duty[0][0] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input n16982;
    input [22:0]pwm_setpoint;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire pwm_out_0__N_582, n16587;
    wire [9:0]half_duty_new_9__N_664;
    
    wire n21848;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    wire [10:0]n49;
    
    wire pause_counter_0__N_612;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire pause_counter_0, n35433;
    wire [10:0]pwm_out_0__N_587;
    
    wire n28691, n28690, n28689, n28688, n28687, n28686, n28685, 
        n28684, n28683, n28682, n27919, pwm_out_0__N_586, n27918, 
        n10, n27917;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n42343, n27916, n42341, n4, n42339, n20, n13, n1, n22, 
        n5, n2, n3, n8, n38078, n13_adj_3561, n5_adj_3562, n18, 
        n16, n17, n15, n27915, n27914, n27913, n27912, n27911, 
        n27910, n27909;
    wire [22:0]n5532;
    
    wire n28301, n28300, n28299, n28298, n28297, n28296, n28295, 
        n28294, n28293, n28292, n28291, n28290, n28289, n28288, 
        n28287, n28286, n28285, n28284, n28283, n28282, n28281, 
        n28280, n28279, n28278, n28277, n28276, n28275, n28274, 
        n28273, n28272, n28271, n28270, n28269, n28268, n28267, 
        n28266, n28265, n28264, n28263, n28262, n28261, n28260, 
        n28259, n37985, n12, n18_adj_3563, n19;
    
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n16587), .D(pwm_out_0__N_582));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_664[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n17573));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n17567));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n17568));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n17569));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n17570));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0] [5]), .C(CLK_c), .D(n21848));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n17572));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1178__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[10]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[9]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[8]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[7]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[6]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[5]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[4]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[3]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[2]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1178__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[1]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 i36306_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_582), .I2(GND_net), 
            .I3(GND_net), .O(n35433));
    defparam i36306_2_lut.LUT_INIT = 16'h1111;
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n35433));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_612));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR count_0__1178__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[0]), .R(n1169));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 count_0__1178_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n28691), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0] [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17185_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_out_0__N_587[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i17185_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 count_0__1178_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n28690), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_11 (.CI(n28690), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n28691));
    SB_LUT4 count_0__1178_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n28689), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_10 (.CI(n28689), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n28690));
    SB_LUT4 count_0__1178_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n28688), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_9 (.CI(n28688), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n28689));
    SB_LUT4 count_0__1178_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n28687), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_8 (.CI(n28687), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n28688));
    SB_LUT4 count_0__1178_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n28686), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_7 (.CI(n28686), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n28687));
    SB_LUT4 count_0__1178_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n28685), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_6 (.CI(n28685), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n28686));
    SB_LUT4 count_0__1178_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n28684), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_5 (.CI(n28684), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n28685));
    SB_LUT4 count_0__1178_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n28683), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_4 (.CI(n28683), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n28684));
    SB_LUT4 count_0__1178_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n28682), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_3 (.CI(n28682), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n28683));
    SB_LUT4 count_0__1178_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1178_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1178_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n28682));
    SB_CARRY pwm_out_0__I_20_13 (.CI(n27919), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_586));
    SB_CARRY pwm_out_0__I_20_12 (.CI(n27918), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27919));
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n27917), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_664[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i17177_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1169), .I3(GND_net), .O(n21848));
    defparam i17177_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY pwm_out_0__I_20_11 (.CI(n27917), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27918));
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n27916), .O(n42343)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(pwm_out_0__N_586), .I1(n42341), .I2(n4), .I3(n42339), 
            .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut (.I0(n10), .I1(\count[0] [10]), .I2(GND_net), .I3(GND_net), 
            .O(n13));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i10_4_lut (.I0(n13), .I1(n20), .I2(n42343), .I3(n1), .O(n22));
    defparam i10_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i31375_4_lut (.I0(n5), .I1(n2), .I2(n3), .I3(n8), .O(n38078));
    defparam i31375_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(n38078), .I1(pause_counter_0), .I2(pwm_out_0__N_582), 
            .I3(n22), .O(n16587));
    defparam i1_4_lut.LUT_INIT = 16'h1303;
    SB_LUT4 i2_4_lut (.I0(\count[0] [5]), .I1(\half_duty[0][3] ), .I2(\half_duty[0] [5]), 
            .I3(\count[0] [3]), .O(n13_adj_3561));   // vhdl/pwm.vhd(80[8:31])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 half_duty_0__9__I_0_47_i5_2_lut (.I0(\half_duty[0][4] ), .I1(\count[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3562));   // vhdl/pwm.vhd(80[8:31])
    defparam half_duty_0__9__I_0_47_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7_3_lut (.I0(n13_adj_3561), .I1(\count[0] [8]), .I2(\count[0] [9]), 
            .I3(GND_net), .O(n18));   // vhdl/pwm.vhd(80[8:31])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut (.I0(\half_duty[0][7] ), .I1(\count[0] [0]), .I2(\count[0] [7]), 
            .I3(\half_duty[0][0] ), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i6_4_lut (.I0(\half_duty[0][2] ), .I1(n5_adj_3562), .I2(\count[0] [2]), 
            .I3(\count[0] [10]), .O(n17));   // vhdl/pwm.vhd(80[8:31])
    defparam i6_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i4_4_lut (.I0(\count[0] [6]), .I1(\half_duty[0][1] ), .I2(\half_duty[0][6] ), 
            .I3(\count[0] [1]), .O(n15));   // vhdl/pwm.vhd(80[8:31])
    defparam i4_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i10_4_lut_adj_840 (.I0(n15), .I1(n17), .I2(n16), .I3(n18), 
            .O(pwm_out_0__N_582));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut_adj_840.LUT_INIT = 16'hfffe;
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_664[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_664[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_664[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(half_duty_new[5]), .C(CLK_c), .D(half_duty_new_9__N_664[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_664[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_664[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY pwm_out_0__I_20_10 (.CI(n27916), .I0(GND_net), .I1(VCC_net), 
            .CO(n27917));
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_587[7]), 
            .I3(n27915), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_9 (.CI(n27915), .I0(GND_net), .I1(pwm_out_0__N_587[7]), 
            .CO(n27916));
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_587[6]), 
            .I3(n27914), .O(n42339)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n27914), .I0(VCC_net), .I1(pwm_out_0__N_587[6]), 
            .CO(n27915));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_587[5]), 
            .I3(n27913), .O(n42341)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_7 (.CI(n27913), .I0(GND_net), .I1(pwm_out_0__N_587[5]), 
            .CO(n27914));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_587[4]), 
            .I3(n27912), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_6 (.CI(n27912), .I0(GND_net), .I1(pwm_out_0__N_587[4]), 
            .CO(n27913));
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_587[3]), 
            .I3(n27911), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_5 (.CI(n27911), .I0(GND_net), .I1(pwm_out_0__N_587[3]), 
            .CO(n27912));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_587[2]), 
            .I3(n27910), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_4 (.CI(n27910), .I0(GND_net), .I1(pwm_out_0__N_587[2]), 
            .CO(n27911));
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_587[1]), 
            .I3(n27909), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_3 (.CI(n27909), .I0(GND_net), .I1(pwm_out_0__N_587[1]), 
            .CO(n27910));
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_587[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_587[0]), 
            .CO(n27909));
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n16982));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 add_2028_24_lut (.I0(GND_net), .I1(n5532[22]), .I2(pwm_setpoint[22]), 
            .I3(n28301), .O(half_duty_new_9__N_664[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2028_23_lut (.I0(GND_net), .I1(n5532[21]), .I2(pwm_setpoint[21]), 
            .I3(n28300), .O(half_duty_new_9__N_664[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2028_23 (.CI(n28300), .I0(n5532[21]), .I1(pwm_setpoint[21]), 
            .CO(n28301));
    SB_LUT4 add_2028_22_lut (.I0(GND_net), .I1(n5532[20]), .I2(pwm_setpoint[20]), 
            .I3(n28299), .O(half_duty_new_9__N_664[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2028_22 (.CI(n28299), .I0(n5532[20]), .I1(pwm_setpoint[20]), 
            .CO(n28300));
    SB_LUT4 add_2028_21_lut (.I0(GND_net), .I1(n5532[19]), .I2(pwm_setpoint[19]), 
            .I3(n28298), .O(half_duty_new_9__N_664[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2028_21 (.CI(n28298), .I0(n5532[19]), .I1(pwm_setpoint[19]), 
            .CO(n28299));
    SB_LUT4 add_2028_20_lut (.I0(GND_net), .I1(n5532[18]), .I2(pwm_setpoint[18]), 
            .I3(n28297), .O(half_duty_new_9__N_664[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2028_20 (.CI(n28297), .I0(n5532[18]), .I1(pwm_setpoint[18]), 
            .CO(n28298));
    SB_LUT4 add_2028_19_lut (.I0(GND_net), .I1(n5532[17]), .I2(pwm_setpoint[17]), 
            .I3(n28296), .O(half_duty_new_9__N_664[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2028_19 (.CI(n28296), .I0(n5532[17]), .I1(pwm_setpoint[17]), 
            .CO(n28297));
    SB_LUT4 add_2028_18_lut (.I0(GND_net), .I1(n5532[16]), .I2(pwm_setpoint[16]), 
            .I3(n28295), .O(half_duty_new_9__N_664[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2028_18 (.CI(n28295), .I0(n5532[16]), .I1(pwm_setpoint[16]), 
            .CO(n28296));
    SB_LUT4 add_2028_17_lut (.I0(GND_net), .I1(n5532[15]), .I2(pwm_setpoint[15]), 
            .I3(n28294), .O(half_duty_new_9__N_664[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2028_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2028_17 (.CI(n28294), .I0(n5532[15]), .I1(pwm_setpoint[15]), 
            .CO(n28295));
    SB_CARRY add_2028_16 (.CI(n28293), .I0(n5532[14]), .I1(pwm_setpoint[14]), 
            .CO(n28294));
    SB_CARRY add_2028_15 (.CI(n28292), .I0(n5532[13]), .I1(pwm_setpoint[13]), 
            .CO(n28293));
    SB_CARRY add_2028_14 (.CI(n28291), .I0(n5532[12]), .I1(pwm_setpoint[12]), 
            .CO(n28292));
    SB_CARRY add_2028_13 (.CI(n28290), .I0(n5532[11]), .I1(pwm_setpoint[11]), 
            .CO(n28291));
    SB_CARRY add_2028_12 (.CI(n28289), .I0(n5532[10]), .I1(pwm_setpoint[10]), 
            .CO(n28290));
    SB_CARRY add_2028_11 (.CI(n28288), .I0(n5532[9]), .I1(pwm_setpoint[9]), 
            .CO(n28289));
    SB_CARRY add_2028_10 (.CI(n28287), .I0(n5532[8]), .I1(pwm_setpoint[8]), 
            .CO(n28288));
    SB_CARRY add_2028_9 (.CI(n28286), .I0(n5532[7]), .I1(pwm_setpoint[7]), 
            .CO(n28287));
    SB_CARRY add_2028_8 (.CI(n28285), .I0(n5532[6]), .I1(pwm_setpoint[6]), 
            .CO(n28286));
    SB_CARRY add_2028_7 (.CI(n28284), .I0(n5532[5]), .I1(pwm_setpoint[5]), 
            .CO(n28285));
    SB_CARRY add_2028_6 (.CI(n28283), .I0(n5532[4]), .I1(pwm_setpoint[4]), 
            .CO(n28284));
    SB_CARRY add_2028_5 (.CI(n28282), .I0(n5532[3]), .I1(pwm_setpoint[3]), 
            .CO(n28283));
    SB_CARRY add_2028_4 (.CI(n28281), .I0(n5532[2]), .I1(pwm_setpoint[2]), 
            .CO(n28282));
    SB_CARRY add_2028_3 (.CI(n28280), .I0(n5532[1]), .I1(pwm_setpoint[1]), 
            .CO(n28281));
    SB_CARRY add_2028_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n28280));
    SB_LUT4 add_2036_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n28279), .O(n5532[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2036_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n28278), .O(n5532[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_22 (.CI(n28278), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n28279));
    SB_LUT4 add_2036_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n28277), .O(n5532[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_21 (.CI(n28277), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n28278));
    SB_LUT4 add_2036_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n28276), .O(n5532[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_20 (.CI(n28276), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n28277));
    SB_LUT4 add_2036_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n28275), .O(n5532[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_19 (.CI(n28275), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n28276));
    SB_LUT4 add_2036_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n28274), .O(n5532[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_18 (.CI(n28274), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n28275));
    SB_LUT4 add_2036_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n28273), .O(n5532[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_17 (.CI(n28273), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n28274));
    SB_LUT4 add_2036_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n28272), .O(n5532[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_16 (.CI(n28272), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n28273));
    SB_LUT4 add_2036_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n28271), .O(n5532[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_15 (.CI(n28271), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n28272));
    SB_LUT4 add_2036_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n28270), .O(n5532[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_14 (.CI(n28270), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n28271));
    SB_LUT4 add_2036_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n28269), .O(n5532[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_13 (.CI(n28269), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n28270));
    SB_LUT4 add_2036_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n28268), .O(n5532[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_12 (.CI(n28268), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n28269));
    SB_LUT4 add_2036_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n28267), .O(n5532[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_11 (.CI(n28267), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n28268));
    SB_LUT4 add_2036_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n28266), .O(n5532[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_10 (.CI(n28266), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n28267));
    SB_LUT4 add_2036_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n28265), .O(n5532[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_9 (.CI(n28265), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n28266));
    SB_LUT4 add_2036_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n28264), .O(n5532[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_8 (.CI(n28264), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n28265));
    SB_LUT4 add_2036_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n28263), .O(n5532[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_7 (.CI(n28263), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n28264));
    SB_LUT4 add_2036_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n28262), .O(n5532[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_6 (.CI(n28262), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n28263));
    SB_LUT4 add_2036_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n28261), .O(n5532[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_5 (.CI(n28261), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n28262));
    SB_LUT4 add_2036_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n28260), .O(n5532[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_4 (.CI(n28260), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n28261));
    SB_LUT4 add_2036_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n28259), .O(n5532[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_3 (.CI(n28259), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n28260));
    SB_LUT4 add_2036_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5532[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2036_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2036_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n28259));
    SB_LUT4 i31283_2_lut (.I0(\count[0] [8]), .I1(\count[0] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n37985));
    defparam i31283_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_841 (.I0(\count[0] [4]), .I1(\count[0] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n12));
    defparam i1_2_lut_adj_841.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut (.I0(n37985), .I1(\count[0] [3]), .I2(\count[0] [10]), 
            .I3(pause_counter_0), .O(n18_adj_3563));
    defparam i7_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i8_4_lut_adj_842 (.I0(\count[0] [9]), .I1(\count[0] [0]), .I2(\count[0] [1]), 
            .I3(\count[0] [2]), .O(n19));
    defparam i8_4_lut_adj_842.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut_adj_843 (.I0(n19), .I1(\count[0] [7]), .I2(n18_adj_3563), 
            .I3(n12), .O(n1169));
    defparam i10_4_lut_adj_843.LUT_INIT = 16'h2000;
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    
endmodule
