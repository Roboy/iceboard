-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Feb 4 2020 22:10:19

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : in std_logic;
    SCL : in std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__56344\ : std_logic;
signal \N__56343\ : std_logic;
signal \N__56342\ : std_logic;
signal \N__56335\ : std_logic;
signal \N__56334\ : std_logic;
signal \N__56333\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56324\ : std_logic;
signal \N__56317\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56315\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56307\ : std_logic;
signal \N__56306\ : std_logic;
signal \N__56299\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56297\ : std_logic;
signal \N__56290\ : std_logic;
signal \N__56289\ : std_logic;
signal \N__56288\ : std_logic;
signal \N__56281\ : std_logic;
signal \N__56280\ : std_logic;
signal \N__56279\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56270\ : std_logic;
signal \N__56263\ : std_logic;
signal \N__56262\ : std_logic;
signal \N__56261\ : std_logic;
signal \N__56254\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56252\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56243\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56235\ : std_logic;
signal \N__56234\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56226\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56218\ : std_logic;
signal \N__56217\ : std_logic;
signal \N__56216\ : std_logic;
signal \N__56209\ : std_logic;
signal \N__56208\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56200\ : std_logic;
signal \N__56199\ : std_logic;
signal \N__56198\ : std_logic;
signal \N__56191\ : std_logic;
signal \N__56190\ : std_logic;
signal \N__56189\ : std_logic;
signal \N__56182\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56180\ : std_logic;
signal \N__56163\ : std_logic;
signal \N__56160\ : std_logic;
signal \N__56157\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56151\ : std_logic;
signal \N__56148\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56145\ : std_logic;
signal \N__56144\ : std_logic;
signal \N__56143\ : std_logic;
signal \N__56140\ : std_logic;
signal \N__56137\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56127\ : std_logic;
signal \N__56126\ : std_logic;
signal \N__56125\ : std_logic;
signal \N__56124\ : std_logic;
signal \N__56119\ : std_logic;
signal \N__56118\ : std_logic;
signal \N__56113\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56111\ : std_logic;
signal \N__56110\ : std_logic;
signal \N__56107\ : std_logic;
signal \N__56102\ : std_logic;
signal \N__56101\ : std_logic;
signal \N__56100\ : std_logic;
signal \N__56099\ : std_logic;
signal \N__56096\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56090\ : std_logic;
signal \N__56083\ : std_logic;
signal \N__56080\ : std_logic;
signal \N__56077\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56069\ : std_logic;
signal \N__56064\ : std_logic;
signal \N__56055\ : std_logic;
signal \N__56046\ : std_logic;
signal \N__56045\ : std_logic;
signal \N__56044\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56036\ : std_logic;
signal \N__56031\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56024\ : std_logic;
signal \N__56021\ : std_logic;
signal \N__56018\ : std_logic;
signal \N__56017\ : std_logic;
signal \N__56014\ : std_logic;
signal \N__56013\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56003\ : std_logic;
signal \N__56002\ : std_logic;
signal \N__55999\ : std_logic;
signal \N__55996\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55987\ : std_logic;
signal \N__55982\ : std_logic;
signal \N__55977\ : std_logic;
signal \N__55968\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55963\ : std_logic;
signal \N__55962\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55957\ : std_logic;
signal \N__55952\ : std_logic;
signal \N__55951\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55947\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55936\ : std_logic;
signal \N__55933\ : std_logic;
signal \N__55930\ : std_logic;
signal \N__55927\ : std_logic;
signal \N__55922\ : std_logic;
signal \N__55921\ : std_logic;
signal \N__55920\ : std_logic;
signal \N__55915\ : std_logic;
signal \N__55912\ : std_logic;
signal \N__55907\ : std_logic;
signal \N__55902\ : std_logic;
signal \N__55899\ : std_logic;
signal \N__55890\ : std_logic;
signal \N__55889\ : std_logic;
signal \N__55884\ : std_logic;
signal \N__55883\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55881\ : std_logic;
signal \N__55878\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55864\ : std_logic;
signal \N__55861\ : std_logic;
signal \N__55854\ : std_logic;
signal \N__55851\ : std_logic;
signal \N__55848\ : std_logic;
signal \N__55845\ : std_logic;
signal \N__55842\ : std_logic;
signal \N__55839\ : std_logic;
signal \N__55836\ : std_logic;
signal \N__55835\ : std_logic;
signal \N__55834\ : std_logic;
signal \N__55833\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55831\ : std_logic;
signal \N__55830\ : std_logic;
signal \N__55829\ : std_logic;
signal \N__55828\ : std_logic;
signal \N__55827\ : std_logic;
signal \N__55826\ : std_logic;
signal \N__55825\ : std_logic;
signal \N__55824\ : std_logic;
signal \N__55823\ : std_logic;
signal \N__55822\ : std_logic;
signal \N__55821\ : std_logic;
signal \N__55820\ : std_logic;
signal \N__55819\ : std_logic;
signal \N__55818\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55816\ : std_logic;
signal \N__55815\ : std_logic;
signal \N__55814\ : std_logic;
signal \N__55813\ : std_logic;
signal \N__55812\ : std_logic;
signal \N__55811\ : std_logic;
signal \N__55810\ : std_logic;
signal \N__55809\ : std_logic;
signal \N__55808\ : std_logic;
signal \N__55807\ : std_logic;
signal \N__55806\ : std_logic;
signal \N__55805\ : std_logic;
signal \N__55804\ : std_logic;
signal \N__55803\ : std_logic;
signal \N__55802\ : std_logic;
signal \N__55801\ : std_logic;
signal \N__55800\ : std_logic;
signal \N__55799\ : std_logic;
signal \N__55798\ : std_logic;
signal \N__55797\ : std_logic;
signal \N__55796\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55794\ : std_logic;
signal \N__55793\ : std_logic;
signal \N__55792\ : std_logic;
signal \N__55791\ : std_logic;
signal \N__55790\ : std_logic;
signal \N__55789\ : std_logic;
signal \N__55788\ : std_logic;
signal \N__55787\ : std_logic;
signal \N__55786\ : std_logic;
signal \N__55785\ : std_logic;
signal \N__55784\ : std_logic;
signal \N__55783\ : std_logic;
signal \N__55782\ : std_logic;
signal \N__55781\ : std_logic;
signal \N__55780\ : std_logic;
signal \N__55779\ : std_logic;
signal \N__55778\ : std_logic;
signal \N__55777\ : std_logic;
signal \N__55776\ : std_logic;
signal \N__55775\ : std_logic;
signal \N__55774\ : std_logic;
signal \N__55773\ : std_logic;
signal \N__55644\ : std_logic;
signal \N__55641\ : std_logic;
signal \N__55638\ : std_logic;
signal \N__55637\ : std_logic;
signal \N__55634\ : std_logic;
signal \N__55633\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55629\ : std_logic;
signal \N__55626\ : std_logic;
signal \N__55623\ : std_logic;
signal \N__55620\ : std_logic;
signal \N__55617\ : std_logic;
signal \N__55612\ : std_logic;
signal \N__55609\ : std_logic;
signal \N__55606\ : std_logic;
signal \N__55603\ : std_logic;
signal \N__55596\ : std_logic;
signal \N__55593\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55591\ : std_logic;
signal \N__55590\ : std_logic;
signal \N__55587\ : std_logic;
signal \N__55584\ : std_logic;
signal \N__55581\ : std_logic;
signal \N__55578\ : std_logic;
signal \N__55573\ : std_logic;
signal \N__55568\ : std_logic;
signal \N__55565\ : std_logic;
signal \N__55560\ : std_logic;
signal \N__55557\ : std_logic;
signal \N__55554\ : std_logic;
signal \N__55551\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55545\ : std_logic;
signal \N__55542\ : std_logic;
signal \N__55539\ : std_logic;
signal \N__55536\ : std_logic;
signal \N__55533\ : std_logic;
signal \N__55530\ : std_logic;
signal \N__55527\ : std_logic;
signal \N__55524\ : std_logic;
signal \N__55521\ : std_logic;
signal \N__55518\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55505\ : std_logic;
signal \N__55504\ : std_logic;
signal \N__55501\ : std_logic;
signal \N__55496\ : std_logic;
signal \N__55491\ : std_logic;
signal \N__55488\ : std_logic;
signal \N__55485\ : std_logic;
signal \N__55482\ : std_logic;
signal \N__55479\ : std_logic;
signal \N__55476\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55467\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55463\ : std_logic;
signal \N__55460\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55452\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55440\ : std_logic;
signal \N__55437\ : std_logic;
signal \N__55436\ : std_logic;
signal \N__55433\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55427\ : std_logic;
signal \N__55422\ : std_logic;
signal \N__55419\ : std_logic;
signal \N__55416\ : std_logic;
signal \N__55415\ : std_logic;
signal \N__55412\ : std_logic;
signal \N__55409\ : std_logic;
signal \N__55404\ : std_logic;
signal \N__55403\ : std_logic;
signal \N__55402\ : std_logic;
signal \N__55401\ : std_logic;
signal \N__55400\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55393\ : std_logic;
signal \N__55390\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55386\ : std_logic;
signal \N__55383\ : std_logic;
signal \N__55380\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55374\ : std_logic;
signal \N__55371\ : std_logic;
signal \N__55368\ : std_logic;
signal \N__55365\ : std_logic;
signal \N__55362\ : std_logic;
signal \N__55359\ : std_logic;
signal \N__55354\ : std_logic;
signal \N__55347\ : std_logic;
signal \N__55344\ : std_logic;
signal \N__55335\ : std_logic;
signal \N__55334\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55332\ : std_logic;
signal \N__55331\ : std_logic;
signal \N__55330\ : std_logic;
signal \N__55329\ : std_logic;
signal \N__55328\ : std_logic;
signal \N__55327\ : std_logic;
signal \N__55326\ : std_logic;
signal \N__55325\ : std_logic;
signal \N__55324\ : std_logic;
signal \N__55323\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55316\ : std_logic;
signal \N__55311\ : std_logic;
signal \N__55310\ : std_logic;
signal \N__55309\ : std_logic;
signal \N__55308\ : std_logic;
signal \N__55307\ : std_logic;
signal \N__55306\ : std_logic;
signal \N__55301\ : std_logic;
signal \N__55298\ : std_logic;
signal \N__55291\ : std_logic;
signal \N__55284\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55278\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55271\ : std_logic;
signal \N__55264\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55262\ : std_logic;
signal \N__55261\ : std_logic;
signal \N__55260\ : std_logic;
signal \N__55255\ : std_logic;
signal \N__55252\ : std_logic;
signal \N__55245\ : std_logic;
signal \N__55242\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55232\ : std_logic;
signal \N__55229\ : std_logic;
signal \N__55224\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55207\ : std_logic;
signal \N__55202\ : std_logic;
signal \N__55191\ : std_logic;
signal \N__55188\ : std_logic;
signal \N__55185\ : std_logic;
signal \N__55182\ : std_logic;
signal \N__55179\ : std_logic;
signal \N__55176\ : std_logic;
signal \N__55175\ : std_logic;
signal \N__55172\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55161\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55146\ : std_logic;
signal \N__55145\ : std_logic;
signal \N__55142\ : std_logic;
signal \N__55139\ : std_logic;
signal \N__55134\ : std_logic;
signal \N__55131\ : std_logic;
signal \N__55130\ : std_logic;
signal \N__55127\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55119\ : std_logic;
signal \N__55116\ : std_logic;
signal \N__55115\ : std_logic;
signal \N__55112\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55104\ : std_logic;
signal \N__55101\ : std_logic;
signal \N__55100\ : std_logic;
signal \N__55097\ : std_logic;
signal \N__55094\ : std_logic;
signal \N__55089\ : std_logic;
signal \N__55086\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55071\ : std_logic;
signal \N__55068\ : std_logic;
signal \N__55067\ : std_logic;
signal \N__55064\ : std_logic;
signal \N__55061\ : std_logic;
signal \N__55056\ : std_logic;
signal \N__55053\ : std_logic;
signal \N__55052\ : std_logic;
signal \N__55049\ : std_logic;
signal \N__55046\ : std_logic;
signal \N__55041\ : std_logic;
signal \N__55038\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55034\ : std_logic;
signal \N__55031\ : std_logic;
signal \N__55030\ : std_logic;
signal \N__55029\ : std_logic;
signal \N__55028\ : std_logic;
signal \N__55027\ : std_logic;
signal \N__55022\ : std_logic;
signal \N__55019\ : std_logic;
signal \N__55016\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55008\ : std_logic;
signal \N__54999\ : std_logic;
signal \N__54996\ : std_logic;
signal \N__54993\ : std_logic;
signal \N__54990\ : std_logic;
signal \N__54987\ : std_logic;
signal \N__54986\ : std_logic;
signal \N__54983\ : std_logic;
signal \N__54980\ : std_logic;
signal \N__54975\ : std_logic;
signal \N__54974\ : std_logic;
signal \N__54971\ : std_logic;
signal \N__54968\ : std_logic;
signal \N__54963\ : std_logic;
signal \N__54960\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54956\ : std_logic;
signal \N__54953\ : std_logic;
signal \N__54948\ : std_logic;
signal \N__54945\ : std_logic;
signal \N__54944\ : std_logic;
signal \N__54941\ : std_logic;
signal \N__54938\ : std_logic;
signal \N__54933\ : std_logic;
signal \N__54930\ : std_logic;
signal \N__54929\ : std_logic;
signal \N__54926\ : std_logic;
signal \N__54923\ : std_logic;
signal \N__54920\ : std_logic;
signal \N__54915\ : std_logic;
signal \N__54912\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54905\ : std_logic;
signal \N__54900\ : std_logic;
signal \N__54897\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54882\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54878\ : std_logic;
signal \N__54875\ : std_logic;
signal \N__54874\ : std_logic;
signal \N__54873\ : std_logic;
signal \N__54870\ : std_logic;
signal \N__54867\ : std_logic;
signal \N__54864\ : std_logic;
signal \N__54861\ : std_logic;
signal \N__54852\ : std_logic;
signal \N__54849\ : std_logic;
signal \N__54848\ : std_logic;
signal \N__54847\ : std_logic;
signal \N__54844\ : std_logic;
signal \N__54841\ : std_logic;
signal \N__54838\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54834\ : std_logic;
signal \N__54831\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54825\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54819\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54805\ : std_logic;
signal \N__54802\ : std_logic;
signal \N__54801\ : std_logic;
signal \N__54798\ : std_logic;
signal \N__54795\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54786\ : std_logic;
signal \N__54783\ : std_logic;
signal \N__54780\ : std_logic;
signal \N__54777\ : std_logic;
signal \N__54774\ : std_logic;
signal \N__54765\ : std_logic;
signal \N__54764\ : std_logic;
signal \N__54763\ : std_logic;
signal \N__54762\ : std_logic;
signal \N__54759\ : std_logic;
signal \N__54756\ : std_logic;
signal \N__54755\ : std_logic;
signal \N__54752\ : std_logic;
signal \N__54749\ : std_logic;
signal \N__54748\ : std_logic;
signal \N__54745\ : std_logic;
signal \N__54742\ : std_logic;
signal \N__54739\ : std_logic;
signal \N__54736\ : std_logic;
signal \N__54733\ : std_logic;
signal \N__54730\ : std_logic;
signal \N__54725\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54708\ : std_logic;
signal \N__54705\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54699\ : std_logic;
signal \N__54698\ : std_logic;
signal \N__54697\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54693\ : std_logic;
signal \N__54690\ : std_logic;
signal \N__54689\ : std_logic;
signal \N__54688\ : std_logic;
signal \N__54685\ : std_logic;
signal \N__54684\ : std_logic;
signal \N__54679\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54671\ : std_logic;
signal \N__54670\ : std_logic;
signal \N__54667\ : std_logic;
signal \N__54664\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54642\ : std_logic;
signal \N__54639\ : std_logic;
signal \N__54638\ : std_logic;
signal \N__54637\ : std_logic;
signal \N__54636\ : std_logic;
signal \N__54635\ : std_logic;
signal \N__54634\ : std_logic;
signal \N__54631\ : std_logic;
signal \N__54628\ : std_logic;
signal \N__54625\ : std_logic;
signal \N__54624\ : std_logic;
signal \N__54623\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54617\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54605\ : std_logic;
signal \N__54602\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54591\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54579\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54570\ : std_logic;
signal \N__54567\ : std_logic;
signal \N__54566\ : std_logic;
signal \N__54565\ : std_logic;
signal \N__54564\ : std_logic;
signal \N__54561\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54553\ : std_logic;
signal \N__54546\ : std_logic;
signal \N__54545\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54543\ : std_logic;
signal \N__54540\ : std_logic;
signal \N__54539\ : std_logic;
signal \N__54536\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54530\ : std_logic;
signal \N__54529\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54527\ : std_logic;
signal \N__54526\ : std_logic;
signal \N__54523\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54521\ : std_logic;
signal \N__54520\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54518\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54516\ : std_logic;
signal \N__54515\ : std_logic;
signal \N__54514\ : std_logic;
signal \N__54513\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54510\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54506\ : std_logic;
signal \N__54505\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54503\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54491\ : std_logic;
signal \N__54484\ : std_logic;
signal \N__54477\ : std_logic;
signal \N__54466\ : std_logic;
signal \N__54465\ : std_logic;
signal \N__54462\ : std_logic;
signal \N__54461\ : std_logic;
signal \N__54460\ : std_logic;
signal \N__54459\ : std_logic;
signal \N__54458\ : std_logic;
signal \N__54457\ : std_logic;
signal \N__54456\ : std_logic;
signal \N__54455\ : std_logic;
signal \N__54452\ : std_logic;
signal \N__54449\ : std_logic;
signal \N__54446\ : std_logic;
signal \N__54443\ : std_logic;
signal \N__54440\ : std_logic;
signal \N__54437\ : std_logic;
signal \N__54434\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54428\ : std_logic;
signal \N__54425\ : std_logic;
signal \N__54424\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54418\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54415\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54413\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54407\ : std_logic;
signal \N__54406\ : std_logic;
signal \N__54405\ : std_logic;
signal \N__54404\ : std_logic;
signal \N__54403\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54400\ : std_logic;
signal \N__54399\ : std_logic;
signal \N__54396\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54392\ : std_logic;
signal \N__54391\ : std_logic;
signal \N__54390\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54386\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54376\ : std_logic;
signal \N__54371\ : std_logic;
signal \N__54366\ : std_logic;
signal \N__54365\ : std_logic;
signal \N__54362\ : std_logic;
signal \N__54361\ : std_logic;
signal \N__54360\ : std_logic;
signal \N__54359\ : std_logic;
signal \N__54358\ : std_logic;
signal \N__54355\ : std_logic;
signal \N__54354\ : std_logic;
signal \N__54353\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54350\ : std_logic;
signal \N__54347\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54345\ : std_logic;
signal \N__54342\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54334\ : std_logic;
signal \N__54325\ : std_logic;
signal \N__54316\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54296\ : std_logic;
signal \N__54295\ : std_logic;
signal \N__54294\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54292\ : std_logic;
signal \N__54291\ : std_logic;
signal \N__54290\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54287\ : std_logic;
signal \N__54286\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54284\ : std_logic;
signal \N__54283\ : std_logic;
signal \N__54282\ : std_logic;
signal \N__54281\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54279\ : std_logic;
signal \N__54278\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54276\ : std_logic;
signal \N__54275\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54273\ : std_logic;
signal \N__54272\ : std_logic;
signal \N__54271\ : std_logic;
signal \N__54270\ : std_logic;
signal \N__54269\ : std_logic;
signal \N__54268\ : std_logic;
signal \N__54267\ : std_logic;
signal \N__54266\ : std_logic;
signal \N__54265\ : std_logic;
signal \N__54264\ : std_logic;
signal \N__54263\ : std_logic;
signal \N__54262\ : std_logic;
signal \N__54259\ : std_logic;
signal \N__54252\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54242\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54232\ : std_logic;
signal \N__54219\ : std_logic;
signal \N__54216\ : std_logic;
signal \N__54207\ : std_logic;
signal \N__54202\ : std_logic;
signal \N__54201\ : std_logic;
signal \N__54198\ : std_logic;
signal \N__54197\ : std_logic;
signal \N__54194\ : std_logic;
signal \N__54191\ : std_logic;
signal \N__54190\ : std_logic;
signal \N__54189\ : std_logic;
signal \N__54188\ : std_logic;
signal \N__54187\ : std_logic;
signal \N__54186\ : std_logic;
signal \N__54185\ : std_logic;
signal \N__54184\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54182\ : std_logic;
signal \N__54181\ : std_logic;
signal \N__54180\ : std_logic;
signal \N__54179\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54176\ : std_logic;
signal \N__54169\ : std_logic;
signal \N__54164\ : std_logic;
signal \N__54151\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54135\ : std_logic;
signal \N__54134\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54128\ : std_logic;
signal \N__54125\ : std_logic;
signal \N__54122\ : std_logic;
signal \N__54121\ : std_logic;
signal \N__54118\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54112\ : std_logic;
signal \N__54109\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54103\ : std_logic;
signal \N__54102\ : std_logic;
signal \N__54099\ : std_logic;
signal \N__54098\ : std_logic;
signal \N__54097\ : std_logic;
signal \N__54096\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54094\ : std_logic;
signal \N__54093\ : std_logic;
signal \N__54092\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54082\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54080\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54078\ : std_logic;
signal \N__54075\ : std_logic;
signal \N__54072\ : std_logic;
signal \N__54069\ : std_logic;
signal \N__54066\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54062\ : std_logic;
signal \N__54059\ : std_logic;
signal \N__54056\ : std_logic;
signal \N__54053\ : std_logic;
signal \N__54052\ : std_logic;
signal \N__54049\ : std_logic;
signal \N__54046\ : std_logic;
signal \N__54043\ : std_logic;
signal \N__54040\ : std_logic;
signal \N__54037\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54019\ : std_logic;
signal \N__54018\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54012\ : std_logic;
signal \N__54011\ : std_logic;
signal \N__54010\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54008\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54005\ : std_logic;
signal \N__54004\ : std_logic;
signal \N__54003\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__54000\ : std_logic;
signal \N__53999\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53995\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53993\ : std_logic;
signal \N__53992\ : std_logic;
signal \N__53991\ : std_logic;
signal \N__53990\ : std_logic;
signal \N__53989\ : std_logic;
signal \N__53988\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53985\ : std_logic;
signal \N__53984\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53982\ : std_logic;
signal \N__53981\ : std_logic;
signal \N__53968\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53955\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53938\ : std_logic;
signal \N__53937\ : std_logic;
signal \N__53936\ : std_logic;
signal \N__53935\ : std_logic;
signal \N__53934\ : std_logic;
signal \N__53933\ : std_logic;
signal \N__53930\ : std_logic;
signal \N__53927\ : std_logic;
signal \N__53926\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53921\ : std_logic;
signal \N__53918\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53915\ : std_logic;
signal \N__53912\ : std_logic;
signal \N__53909\ : std_logic;
signal \N__53906\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53904\ : std_logic;
signal \N__53903\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53897\ : std_logic;
signal \N__53896\ : std_logic;
signal \N__53893\ : std_logic;
signal \N__53892\ : std_logic;
signal \N__53891\ : std_logic;
signal \N__53890\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53888\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53882\ : std_logic;
signal \N__53879\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53867\ : std_logic;
signal \N__53860\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53846\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53828\ : std_logic;
signal \N__53825\ : std_logic;
signal \N__53822\ : std_logic;
signal \N__53819\ : std_logic;
signal \N__53818\ : std_logic;
signal \N__53815\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53810\ : std_logic;
signal \N__53809\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53807\ : std_logic;
signal \N__53802\ : std_logic;
signal \N__53797\ : std_logic;
signal \N__53794\ : std_logic;
signal \N__53793\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53784\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53776\ : std_logic;
signal \N__53769\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53764\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53758\ : std_logic;
signal \N__53747\ : std_logic;
signal \N__53738\ : std_logic;
signal \N__53729\ : std_logic;
signal \N__53718\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53716\ : std_logic;
signal \N__53715\ : std_logic;
signal \N__53714\ : std_logic;
signal \N__53713\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53708\ : std_logic;
signal \N__53707\ : std_logic;
signal \N__53704\ : std_logic;
signal \N__53701\ : std_logic;
signal \N__53698\ : std_logic;
signal \N__53695\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53688\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53679\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53673\ : std_logic;
signal \N__53670\ : std_logic;
signal \N__53667\ : std_logic;
signal \N__53664\ : std_logic;
signal \N__53661\ : std_logic;
signal \N__53658\ : std_logic;
signal \N__53655\ : std_logic;
signal \N__53652\ : std_logic;
signal \N__53649\ : std_logic;
signal \N__53646\ : std_logic;
signal \N__53643\ : std_logic;
signal \N__53640\ : std_logic;
signal \N__53639\ : std_logic;
signal \N__53638\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53627\ : std_logic;
signal \N__53624\ : std_logic;
signal \N__53621\ : std_logic;
signal \N__53620\ : std_logic;
signal \N__53617\ : std_logic;
signal \N__53616\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53614\ : std_logic;
signal \N__53613\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53611\ : std_logic;
signal \N__53610\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53608\ : std_logic;
signal \N__53607\ : std_logic;
signal \N__53596\ : std_logic;
signal \N__53593\ : std_logic;
signal \N__53590\ : std_logic;
signal \N__53587\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53585\ : std_logic;
signal \N__53584\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53580\ : std_logic;
signal \N__53579\ : std_logic;
signal \N__53578\ : std_logic;
signal \N__53577\ : std_logic;
signal \N__53576\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53572\ : std_logic;
signal \N__53571\ : std_logic;
signal \N__53568\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53564\ : std_logic;
signal \N__53563\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53561\ : std_logic;
signal \N__53560\ : std_logic;
signal \N__53559\ : std_logic;
signal \N__53558\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53546\ : std_logic;
signal \N__53543\ : std_logic;
signal \N__53536\ : std_logic;
signal \N__53531\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53516\ : std_logic;
signal \N__53507\ : std_logic;
signal \N__53498\ : std_logic;
signal \N__53495\ : std_logic;
signal \N__53492\ : std_logic;
signal \N__53491\ : std_logic;
signal \N__53484\ : std_logic;
signal \N__53471\ : std_logic;
signal \N__53468\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53454\ : std_logic;
signal \N__53453\ : std_logic;
signal \N__53452\ : std_logic;
signal \N__53451\ : std_logic;
signal \N__53450\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53446\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53441\ : std_logic;
signal \N__53440\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53434\ : std_logic;
signal \N__53433\ : std_logic;
signal \N__53432\ : std_logic;
signal \N__53429\ : std_logic;
signal \N__53426\ : std_logic;
signal \N__53425\ : std_logic;
signal \N__53422\ : std_logic;
signal \N__53419\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53413\ : std_logic;
signal \N__53412\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53399\ : std_logic;
signal \N__53388\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53386\ : std_logic;
signal \N__53385\ : std_logic;
signal \N__53380\ : std_logic;
signal \N__53377\ : std_logic;
signal \N__53370\ : std_logic;
signal \N__53359\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53301\ : std_logic;
signal \N__53292\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53279\ : std_logic;
signal \N__53276\ : std_logic;
signal \N__53273\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53254\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53252\ : std_logic;
signal \N__53251\ : std_logic;
signal \N__53248\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53234\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53213\ : std_logic;
signal \N__53202\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53198\ : std_logic;
signal \N__53197\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53193\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53191\ : std_logic;
signal \N__53190\ : std_logic;
signal \N__53189\ : std_logic;
signal \N__53188\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53169\ : std_logic;
signal \N__53164\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53159\ : std_logic;
signal \N__53158\ : std_logic;
signal \N__53155\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53153\ : std_logic;
signal \N__53152\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53102\ : std_logic;
signal \N__53101\ : std_logic;
signal \N__53100\ : std_logic;
signal \N__53099\ : std_logic;
signal \N__53096\ : std_logic;
signal \N__53095\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53091\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53086\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53075\ : std_logic;
signal \N__53066\ : std_logic;
signal \N__53057\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53041\ : std_logic;
signal \N__53032\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53017\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53004\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__53001\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52980\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52974\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52972\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52957\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52947\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52932\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52915\ : std_logic;
signal \N__52910\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52904\ : std_logic;
signal \N__52903\ : std_logic;
signal \N__52902\ : std_logic;
signal \N__52901\ : std_logic;
signal \N__52900\ : std_logic;
signal \N__52899\ : std_logic;
signal \N__52898\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52896\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52893\ : std_logic;
signal \N__52892\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52887\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52865\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52855\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52837\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52821\ : std_logic;
signal \N__52818\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52787\ : std_logic;
signal \N__52786\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52761\ : std_logic;
signal \N__52758\ : std_logic;
signal \N__52753\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52735\ : std_logic;
signal \N__52734\ : std_logic;
signal \N__52733\ : std_logic;
signal \N__52732\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52730\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52726\ : std_logic;
signal \N__52725\ : std_logic;
signal \N__52724\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52721\ : std_logic;
signal \N__52718\ : std_logic;
signal \N__52717\ : std_logic;
signal \N__52714\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52712\ : std_logic;
signal \N__52711\ : std_logic;
signal \N__52704\ : std_logic;
signal \N__52697\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52689\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52662\ : std_logic;
signal \N__52651\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52624\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52609\ : std_logic;
signal \N__52600\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52576\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52560\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52557\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52539\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52521\ : std_logic;
signal \N__52514\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52485\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52453\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52428\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52412\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52365\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52359\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52355\ : std_logic;
signal \N__52352\ : std_logic;
signal \N__52349\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52341\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52337\ : std_logic;
signal \N__52334\ : std_logic;
signal \N__52331\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52322\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52313\ : std_logic;
signal \N__52310\ : std_logic;
signal \N__52305\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52296\ : std_logic;
signal \N__52293\ : std_logic;
signal \N__52290\ : std_logic;
signal \N__52287\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52277\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52274\ : std_logic;
signal \N__52271\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52249\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52242\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52239\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52197\ : std_logic;
signal \N__52196\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52180\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52164\ : std_logic;
signal \N__52161\ : std_logic;
signal \N__52158\ : std_logic;
signal \N__52155\ : std_logic;
signal \N__52152\ : std_logic;
signal \N__52149\ : std_logic;
signal \N__52146\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52136\ : std_logic;
signal \N__52133\ : std_logic;
signal \N__52130\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52116\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52109\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52106\ : std_logic;
signal \N__52103\ : std_logic;
signal \N__52100\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52095\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52088\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52085\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52082\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52061\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52057\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52053\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52049\ : std_logic;
signal \N__52046\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52043\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52037\ : std_logic;
signal \N__52036\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51990\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51960\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51953\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51944\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51936\ : std_logic;
signal \N__51933\ : std_logic;
signal \N__51930\ : std_logic;
signal \N__51927\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51849\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51839\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51807\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51803\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51788\ : std_logic;
signal \N__51787\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51771\ : std_logic;
signal \N__51768\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51761\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51749\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51745\ : std_logic;
signal \N__51742\ : std_logic;
signal \N__51739\ : std_logic;
signal \N__51732\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51719\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51713\ : std_logic;
signal \N__51710\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51668\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51662\ : std_logic;
signal \N__51659\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51628\ : std_logic;
signal \N__51625\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51609\ : std_logic;
signal \N__51606\ : std_logic;
signal \N__51603\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51591\ : std_logic;
signal \N__51590\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51576\ : std_logic;
signal \N__51573\ : std_logic;
signal \N__51570\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51567\ : std_logic;
signal \N__51564\ : std_logic;
signal \N__51557\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51547\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51506\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51488\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51468\ : std_logic;
signal \N__51465\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51429\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51422\ : std_logic;
signal \N__51419\ : std_logic;
signal \N__51416\ : std_logic;
signal \N__51413\ : std_logic;
signal \N__51410\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51401\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51387\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51379\ : std_logic;
signal \N__51376\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51366\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51351\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51318\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51311\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51294\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51288\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51281\ : std_logic;
signal \N__51278\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51274\ : std_logic;
signal \N__51271\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51255\ : std_logic;
signal \N__51252\ : std_logic;
signal \N__51249\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51243\ : std_logic;
signal \N__51236\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51202\ : std_logic;
signal \N__51199\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51180\ : std_logic;
signal \N__51177\ : std_logic;
signal \N__51174\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51147\ : std_logic;
signal \N__51144\ : std_logic;
signal \N__51141\ : std_logic;
signal \N__51138\ : std_logic;
signal \N__51137\ : std_logic;
signal \N__51134\ : std_logic;
signal \N__51131\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51125\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51099\ : std_logic;
signal \N__51098\ : std_logic;
signal \N__51095\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51091\ : std_logic;
signal \N__51088\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51072\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51052\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51046\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51036\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51017\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51010\ : std_logic;
signal \N__51007\ : std_logic;
signal \N__51004\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50988\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50958\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50947\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50920\ : std_logic;
signal \N__50917\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50875\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50840\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50792\ : std_logic;
signal \N__50789\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50765\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50708\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50653\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50632\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50626\ : std_logic;
signal \N__50623\ : std_logic;
signal \N__50618\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50569\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50366\ : std_logic;
signal \N__50363\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50102\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50096\ : std_logic;
signal \N__50093\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50064\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49667\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49647\ : std_logic;
signal \N__49644\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49097\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48915\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48567\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44891\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44814\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44756\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42865\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41971\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal n12703 : std_logic;
signal n12704 : std_logic;
signal n12705 : std_logic;
signal n12706 : std_logic;
signal n12707 : std_logic;
signal n12708 : std_logic;
signal n12709 : std_logic;
signal n12710 : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal n12711 : std_logic;
signal n12712 : std_logic;
signal n12713 : std_logic;
signal n12714 : std_logic;
signal n12715 : std_logic;
signal n12716 : std_logic;
signal n12717 : std_logic;
signal n12718 : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal n12719 : std_logic;
signal n12720 : std_logic;
signal n12721 : std_logic;
signal n12722 : std_logic;
signal n12723 : std_logic;
signal n12724 : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal n12725 : std_logic;
signal n12726 : std_logic;
signal n12727 : std_logic;
signal n12728 : std_logic;
signal n12729 : std_logic;
signal n12730 : std_logic;
signal n12731 : std_logic;
signal n12732 : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal n12733 : std_logic;
signal n12734 : std_logic;
signal n12735 : std_logic;
signal n12736 : std_logic;
signal n12737 : std_logic;
signal n12738 : std_logic;
signal n12739 : std_logic;
signal n12740 : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal n12741 : std_logic;
signal n12742 : std_logic;
signal n12743 : std_logic;
signal n12744 : std_logic;
signal n12745 : std_logic;
signal n12746 : std_logic;
signal n12747 : std_logic;
signal \n2719_cascade_\ : std_logic;
signal n2486 : std_logic;
signal \n2816_cascade_\ : std_logic;
signal \n2829_cascade_\ : std_logic;
signal \n13845_cascade_\ : std_logic;
signal n14702 : std_logic;
signal \bfn_1_26_0_\ : std_logic;
signal n12797 : std_logic;
signal n12798 : std_logic;
signal n12799 : std_logic;
signal n12800 : std_logic;
signal n12801 : std_logic;
signal n12802 : std_logic;
signal n12803 : std_logic;
signal n12804 : std_logic;
signal \bfn_1_27_0_\ : std_logic;
signal n12805 : std_logic;
signal n12806 : std_logic;
signal n12807 : std_logic;
signal n12808 : std_logic;
signal n12809 : std_logic;
signal n12810 : std_logic;
signal n12811 : std_logic;
signal n12812 : std_logic;
signal \bfn_1_28_0_\ : std_logic;
signal n12813 : std_logic;
signal n12814 : std_logic;
signal n12815 : std_logic;
signal n12816 : std_logic;
signal n12817 : std_logic;
signal n12818 : std_logic;
signal n12819 : std_logic;
signal n12820 : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal n2876 : std_logic;
signal n12821 : std_logic;
signal n12822 : std_logic;
signal n11956 : std_logic;
signal n2899 : std_logic;
signal n2833 : std_logic;
signal n2900 : std_logic;
signal \n2833_cascade_\ : std_logic;
signal \n2932_cascade_\ : std_logic;
signal n2901 : std_logic;
signal \n2933_cascade_\ : std_logic;
signal \bfn_1_31_0_\ : std_logic;
signal \debounce.n13016\ : std_logic;
signal \debounce.n13017\ : std_logic;
signal \debounce.n13018\ : std_logic;
signal \debounce.n13019\ : std_logic;
signal \debounce.n13020\ : std_logic;
signal \debounce.n13021\ : std_logic;
signal \debounce.n13022\ : std_logic;
signal \debounce.n13023\ : std_logic;
signal \bfn_1_32_0_\ : std_logic;
signal \debounce.n13024\ : std_logic;
signal n2501 : std_logic;
signal n2500 : std_logic;
signal \n2433_cascade_\ : std_logic;
signal \n2532_cascade_\ : std_logic;
signal n2498 : std_logic;
signal n2487 : std_logic;
signal n2497 : std_logic;
signal n2499 : std_logic;
signal n2496 : std_logic;
signal \n2418_cascade_\ : std_logic;
signal n2495 : std_logic;
signal \n2428_cascade_\ : std_logic;
signal \n2527_cascade_\ : std_logic;
signal n2488 : std_logic;
signal n2493 : std_logic;
signal n2490 : std_logic;
signal n2418 : std_logic;
signal n2485 : std_logic;
signal n2491 : std_logic;
signal n2481 : std_logic;
signal n14310 : std_logic;
signal n2494 : std_logic;
signal n2483 : std_logic;
signal n2416 : std_logic;
signal n2480 : std_logic;
signal n2482 : std_logic;
signal \n14650_cascade_\ : std_logic;
signal n2595 : std_logic;
signal n2528 : std_logic;
signal \n2627_cascade_\ : std_logic;
signal n14646 : std_logic;
signal n2520 : std_logic;
signal n2587 : std_logic;
signal n2589 : std_logic;
signal n2522 : std_logic;
signal n2596 : std_logic;
signal \n2628_cascade_\ : std_logic;
signal n14644 : std_logic;
signal n2527 : std_logic;
signal n2594 : std_logic;
signal n2579 : std_logic;
signal n2586 : std_logic;
signal n2519 : std_logic;
signal n2484 : std_logic;
signal n2583 : std_logic;
signal \n2516_cascade_\ : std_logic;
signal n2588 : std_logic;
signal n2580 : std_logic;
signal \n2612_cascade_\ : std_logic;
signal n2801 : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal n12772 : std_logic;
signal n2799 : std_logic;
signal n12773 : std_logic;
signal n2798 : std_logic;
signal n12774 : std_logic;
signal n2797 : std_logic;
signal n12775 : std_logic;
signal n12776 : std_logic;
signal n12777 : std_logic;
signal n12778 : std_logic;
signal n12779 : std_logic;
signal \bfn_2_24_0_\ : std_logic;
signal n12780 : std_logic;
signal n12781 : std_logic;
signal n12782 : std_logic;
signal n12783 : std_logic;
signal n12784 : std_logic;
signal n12785 : std_logic;
signal n2719 : std_logic;
signal n2786 : std_logic;
signal n12786 : std_logic;
signal n12787 : std_logic;
signal n2785 : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal n2784 : std_logic;
signal n12788 : std_logic;
signal n2783 : std_logic;
signal n12789 : std_logic;
signal n2782 : std_logic;
signal n12790 : std_logic;
signal n12791 : std_logic;
signal n12792 : std_logic;
signal n12793 : std_logic;
signal n12794 : std_logic;
signal n12795 : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal n12796 : std_logic;
signal \n14158_cascade_\ : std_logic;
signal n2790 : std_logic;
signal \n2742_cascade_\ : std_logic;
signal n2789 : std_logic;
signal n2711 : std_logic;
signal n2778 : std_logic;
signal n2781 : std_logic;
signal n2714 : std_logic;
signal n2800 : std_logic;
signal n2832 : std_logic;
signal n2794 : std_logic;
signal n2887 : std_logic;
signal n2779 : std_logic;
signal \n2811_cascade_\ : std_logic;
signal n14708 : std_logic;
signal n2780 : std_logic;
signal n2817 : std_logic;
signal n2884 : std_logic;
signal n2877 : std_logic;
signal n2897 : std_logic;
signal n2830 : std_logic;
signal n2811 : std_logic;
signal n2878 : std_logic;
signal \bfn_2_29_0_\ : std_logic;
signal n2933 : std_logic;
signal n3000 : std_logic;
signal n12823 : std_logic;
signal n12824 : std_logic;
signal n12825 : std_logic;
signal n12826 : std_logic;
signal n12827 : std_logic;
signal n12828 : std_logic;
signal n12829 : std_logic;
signal n12830 : std_logic;
signal \bfn_2_30_0_\ : std_logic;
signal n12831 : std_logic;
signal n12832 : std_logic;
signal n12833 : std_logic;
signal n12834 : std_logic;
signal n12835 : std_logic;
signal n12836 : std_logic;
signal n12837 : std_logic;
signal n12838 : std_logic;
signal \bfn_2_31_0_\ : std_logic;
signal n12839 : std_logic;
signal n12840 : std_logic;
signal n12841 : std_logic;
signal n12842 : std_logic;
signal n12843 : std_logic;
signal n12844 : std_logic;
signal n12845 : std_logic;
signal n12846 : std_logic;
signal \bfn_2_32_0_\ : std_logic;
signal n12847 : std_logic;
signal n12848 : std_logic;
signal n12849 : std_logic;
signal \debounce.cnt_reg_0\ : std_logic;
signal \debounce.cnt_reg_7\ : std_logic;
signal \debounce.cnt_reg_1\ : std_logic;
signal \debounce.cnt_reg_2\ : std_logic;
signal \debounce.cnt_reg_9\ : std_logic;
signal \debounce.cnt_reg_8\ : std_logic;
signal \debounce.cnt_reg_4\ : std_logic;
signal \debounce.cnt_reg_5\ : std_logic;
signal n2976 : std_logic;
signal n2432 : std_logic;
signal \n2432_cascade_\ : std_logic;
signal n2433 : std_logic;
signal n2431 : std_logic;
signal n2430 : std_logic;
signal \n11946_cascade_\ : std_logic;
signal n2429 : std_logic;
signal n2427 : std_logic;
signal n2424 : std_logic;
signal \n2427_cascade_\ : std_logic;
signal n2428 : std_logic;
signal n2529 : std_logic;
signal n11942 : std_logic;
signal n13816 : std_logic;
signal \n14622_cascade_\ : std_logic;
signal n14638 : std_logic;
signal n2420 : std_logic;
signal \n2420_cascade_\ : std_logic;
signal n14612 : std_logic;
signal n14616 : std_logic;
signal n2426 : std_logic;
signal n2421 : std_logic;
signal n2413 : std_logic;
signal n2423 : std_logic;
signal \n2425_cascade_\ : std_logic;
signal n14632 : std_logic;
signal n2419 : std_logic;
signal n2415 : std_logic;
signal \n14456_cascade_\ : std_logic;
signal \n2346_cascade_\ : std_logic;
signal n2417 : std_logic;
signal n2414 : std_logic;
signal n13790 : std_logic;
signal n14318 : std_logic;
signal \n2328_cascade_\ : std_logic;
signal \n14442_cascade_\ : std_logic;
signal \n14448_cascade_\ : std_logic;
signal n14450 : std_logic;
signal n2593 : std_logic;
signal n2422 : std_logic;
signal n2489 : std_logic;
signal n2521 : std_logic;
signal n2526 : std_logic;
signal \n2521_cascade_\ : std_logic;
signal n14312 : std_logic;
signal n14324 : std_logic;
signal n2516 : std_logic;
signal n2512 : std_logic;
signal n2513 : std_logic;
signal \n14330_cascade_\ : std_logic;
signal n2511 : std_logic;
signal n2523 : std_logic;
signal \n2544_cascade_\ : std_logic;
signal n2590 : std_logic;
signal n2591 : std_logic;
signal n2530 : std_logic;
signal n2597 : std_logic;
signal \n2629_cascade_\ : std_logic;
signal n14656 : std_logic;
signal n2601 : std_logic;
signal n2584 : std_logic;
signal n2517 : std_logic;
signal n2582 : std_logic;
signal n2515 : std_logic;
signal n2531 : std_logic;
signal n2598 : std_logic;
signal n2727 : std_logic;
signal n2585 : std_logic;
signal n2518 : std_logic;
signal n14658 : std_logic;
signal \n2617_cascade_\ : std_logic;
signal n2514 : std_logic;
signal n2581 : std_logic;
signal \n2613_cascade_\ : std_logic;
signal n14664 : std_logic;
signal \n14670_cascade_\ : std_logic;
signal \n2643_cascade_\ : std_logic;
signal n2713 : std_logic;
signal n2592 : std_logic;
signal \n14889_cascade_\ : std_logic;
signal n2525 : std_logic;
signal \n2721_cascade_\ : std_logic;
signal n2717 : std_logic;
signal n2718 : std_logic;
signal \n14140_cascade_\ : std_logic;
signal n14138 : std_logic;
signal n2716 : std_logic;
signal n2715 : std_logic;
signal \n14146_cascade_\ : std_logic;
signal n14152 : std_logic;
signal n2722 : std_logic;
signal n2787 : std_logic;
signal n2795 : std_logic;
signal n2728 : std_logic;
signal n2712 : std_logic;
signal n2725 : std_logic;
signal n2792 : std_logic;
signal n2721 : std_logic;
signal n2788 : std_logic;
signal n2793 : std_logic;
signal n2889 : std_logic;
signal \n2921_cascade_\ : std_logic;
signal n2888 : std_logic;
signal n2791 : std_logic;
signal n2822 : std_logic;
signal \n2823_cascade_\ : std_logic;
signal n2821 : std_logic;
signal n2777 : std_logic;
signal n2710 : std_logic;
signal n2809 : std_logic;
signal n2810 : std_logic;
signal n2808 : std_logic;
signal \n2809_cascade_\ : std_logic;
signal n14714 : std_logic;
signal n2823 : std_logic;
signal \n2841_cascade_\ : std_logic;
signal n2890 : std_logic;
signal n2920 : std_logic;
signal n2987 : std_logic;
signal n2898 : std_logic;
signal n2831 : std_logic;
signal n2879 : std_logic;
signal n2812 : std_logic;
signal \n2911_cascade_\ : std_logic;
signal n2829 : std_logic;
signal n2896 : std_logic;
signal n2893 : std_logic;
signal n2826 : std_logic;
signal n2882 : std_logic;
signal n2815 : std_logic;
signal n2813 : std_logic;
signal n2880 : std_logic;
signal \bfn_3_29_0_\ : std_logic;
signal n12850 : std_logic;
signal n12851 : std_logic;
signal n12852 : std_logic;
signal n12853 : std_logic;
signal n12854 : std_logic;
signal n12855 : std_logic;
signal n12856 : std_logic;
signal n12857 : std_logic;
signal \bfn_3_30_0_\ : std_logic;
signal n12858 : std_logic;
signal n12859 : std_logic;
signal n12860 : std_logic;
signal n12861 : std_logic;
signal n12862 : std_logic;
signal n12863 : std_logic;
signal n3086 : std_logic;
signal n12864 : std_logic;
signal n12865 : std_logic;
signal \bfn_3_31_0_\ : std_logic;
signal n12866 : std_logic;
signal n12867 : std_logic;
signal n12868 : std_logic;
signal n12869 : std_logic;
signal n12870 : std_logic;
signal n12871 : std_logic;
signal n12872 : std_logic;
signal n12873 : std_logic;
signal \bfn_3_32_0_\ : std_logic;
signal n12874 : std_logic;
signal n12875 : std_logic;
signal n12876 : std_logic;
signal n12877 : std_logic;
signal \debounce.cnt_reg_6\ : std_logic;
signal \debounce.n16\ : std_logic;
signal \debounce.cnt_reg_3\ : std_logic;
signal \debounce.n17\ : std_logic;
signal n2401 : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal n2400 : std_logic;
signal n12682 : std_logic;
signal n2399 : std_logic;
signal n12683 : std_logic;
signal n2398 : std_logic;
signal n12684 : std_logic;
signal n2397 : std_logic;
signal n12685 : std_logic;
signal n2329 : std_logic;
signal n2396 : std_logic;
signal n12686 : std_logic;
signal n2328 : std_logic;
signal n2395 : std_logic;
signal n12687 : std_logic;
signal n2394 : std_logic;
signal n12688 : std_logic;
signal n12689 : std_logic;
signal n2393 : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal n2392 : std_logic;
signal n12690 : std_logic;
signal n2391 : std_logic;
signal n12691 : std_logic;
signal n2390 : std_logic;
signal n12692 : std_logic;
signal n2389 : std_logic;
signal n12693 : std_logic;
signal n2388 : std_logic;
signal n12694 : std_logic;
signal n2387 : std_logic;
signal n12695 : std_logic;
signal n2386 : std_logic;
signal n12696 : std_logic;
signal n12697 : std_logic;
signal n2385 : std_logic;
signal \bfn_4_19_0_\ : std_logic;
signal n2384 : std_logic;
signal n12698 : std_logic;
signal n2383 : std_logic;
signal n12699 : std_logic;
signal n2382 : std_logic;
signal n12700 : std_logic;
signal n2381 : std_logic;
signal n12701 : std_logic;
signal n12702 : std_logic;
signal n2412 : std_logic;
signal n2314_adj_622 : std_logic;
signal n2327 : std_logic;
signal \n2327_cascade_\ : std_logic;
signal n2326 : std_logic;
signal n14440 : std_logic;
signal n2492 : std_logic;
signal n2425 : std_logic;
signal n2524 : std_logic;
signal n2318 : std_logic;
signal n2320 : std_logic;
signal n2319 : std_logic;
signal \bfn_4_21_0_\ : std_logic;
signal n2700 : std_logic;
signal n12748 : std_logic;
signal n12749 : std_logic;
signal n12750 : std_logic;
signal n12751 : std_logic;
signal n2629 : std_logic;
signal n2696 : std_logic;
signal n12752 : std_logic;
signal n2628 : std_logic;
signal n2695 : std_logic;
signal n12753 : std_logic;
signal n2627 : std_logic;
signal n2694 : std_logic;
signal n12754 : std_logic;
signal n12755 : std_logic;
signal n2626 : std_logic;
signal n2693 : std_logic;
signal \bfn_4_22_0_\ : std_logic;
signal n2625 : std_logic;
signal n2692 : std_logic;
signal n12756 : std_logic;
signal n2624 : std_logic;
signal n2691 : std_logic;
signal n12757 : std_logic;
signal n2623 : std_logic;
signal n2690 : std_logic;
signal n12758 : std_logic;
signal n2622 : std_logic;
signal n2689 : std_logic;
signal n12759 : std_logic;
signal n12760 : std_logic;
signal n2620 : std_logic;
signal n2687 : std_logic;
signal n12761 : std_logic;
signal n2619 : std_logic;
signal n2686 : std_logic;
signal n12762 : std_logic;
signal n12763 : std_logic;
signal n2618 : std_logic;
signal n2685 : std_logic;
signal \bfn_4_23_0_\ : std_logic;
signal n2617 : std_logic;
signal n2684 : std_logic;
signal n12764 : std_logic;
signal n2616 : std_logic;
signal n2683 : std_logic;
signal n12765 : std_logic;
signal n2615 : std_logic;
signal n2682 : std_logic;
signal n12766 : std_logic;
signal n2614 : std_logic;
signal n2681 : std_logic;
signal n12767 : std_logic;
signal n2613 : std_logic;
signal n2680 : std_logic;
signal n12768 : std_logic;
signal n2612 : std_logic;
signal n2679 : std_logic;
signal n12769 : std_logic;
signal n2611 : std_logic;
signal n2678 : std_logic;
signal n12770 : std_logic;
signal n12771 : std_logic;
signal n2610 : std_logic;
signal \bfn_4_24_0_\ : std_logic;
signal n2709 : std_logic;
signal n2816 : std_logic;
signal n2883 : std_logic;
signal n2621 : std_logic;
signal n2688 : std_logic;
signal n2720 : std_logic;
signal n2726 : std_logic;
signal n2724 : std_logic;
signal \n2720_cascade_\ : std_logic;
signal n2723 : std_logic;
signal n14136 : std_logic;
signal n2699 : std_logic;
signal n2698 : std_logic;
signal n2820 : std_logic;
signal \n14688_cascade_\ : std_logic;
signal n14690 : std_logic;
signal n14696 : std_logic;
signal \ENCODER0_B_N\ : std_logic;
signal n2697 : std_logic;
signal n2630 : std_logic;
signal n2731 : std_logic;
signal n2730 : std_logic;
signal \n2729_cascade_\ : std_logic;
signal n13796 : std_logic;
signal n3094 : std_logic;
signal n2701 : std_logic;
signal n2733 : std_logic;
signal \n2733_cascade_\ : std_logic;
signal n2732 : std_logic;
signal n11936 : std_logic;
signal n2729 : std_logic;
signal n2796 : std_logic;
signal n2819 : std_logic;
signal n2886 : std_logic;
signal \n2918_cascade_\ : std_logic;
signal n2827 : std_logic;
signal n2894 : std_logic;
signal \n2926_cascade_\ : std_logic;
signal n14346 : std_logic;
signal \n14336_cascade_\ : std_logic;
signal \n14352_cascade_\ : std_logic;
signal n14350 : std_logic;
signal n2828 : std_logic;
signal n2895 : std_logic;
signal n2885 : std_logic;
signal n2818 : std_logic;
signal n2881 : std_logic;
signal n2814 : std_logic;
signal n12038 : std_logic;
signal n14358 : std_logic;
signal \n14360_cascade_\ : std_logic;
signal n14366 : std_logic;
signal n2927 : std_logic;
signal n2994 : std_logic;
signal n2909 : std_logic;
signal n2907 : std_logic;
signal n14372 : std_logic;
signal n2929 : std_logic;
signal \n2940_cascade_\ : std_logic;
signal n2996 : std_logic;
signal n2921 : std_logic;
signal n2988 : std_logic;
signal n3083 : std_logic;
signal n2995 : std_logic;
signal n2928 : std_logic;
signal n2997 : std_logic;
signal n2930 : std_logic;
signal n3096 : std_logic;
signal \n3029_cascade_\ : std_logic;
signal n2991 : std_logic;
signal n3019 : std_logic;
signal \n3023_cascade_\ : std_logic;
signal n2922 : std_logic;
signal n2989 : std_logic;
signal n3078 : std_logic;
signal n3075 : std_logic;
signal n2984 : std_logic;
signal n2917 : std_logic;
signal n2931 : std_logic;
signal n2998 : std_logic;
signal n3097 : std_logic;
signal \n3030_cascade_\ : std_logic;
signal n3020 : std_logic;
signal n3087 : std_logic;
signal n2985 : std_logic;
signal n2918 : std_logic;
signal n2911 : std_logic;
signal n2978 : std_logic;
signal n2825 : std_logic;
signal n2892 : std_logic;
signal n2924 : std_logic;
signal n2913 : std_logic;
signal n2980 : std_logic;
signal n2915 : std_logic;
signal n2982 : std_logic;
signal n2912 : std_logic;
signal n2979 : std_logic;
signal n2919 : std_logic;
signal n2986 : std_logic;
signal n3016 : std_logic;
signal \n3018_cascade_\ : std_logic;
signal n2914 : std_logic;
signal n2981 : std_logic;
signal n2908 : std_logic;
signal n2975 : std_logic;
signal n3074 : std_logic;
signal \n3007_cascade_\ : std_logic;
signal n2910 : std_logic;
signal n2977 : std_logic;
signal \debounce.reg_A_2\ : std_logic;
signal \debounce.cnt_next_9__N_424\ : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal n12643 : std_logic;
signal n12644 : std_logic;
signal n12645 : std_logic;
signal n12646 : std_logic;
signal n12647 : std_logic;
signal n12648 : std_logic;
signal n12649 : std_logic;
signal n12650 : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal n12651 : std_logic;
signal n12652 : std_logic;
signal n12653 : std_logic;
signal n12654 : std_logic;
signal n12655 : std_logic;
signal n12656 : std_logic;
signal n12657 : std_logic;
signal n12658 : std_logic;
signal \bfn_5_19_0_\ : std_logic;
signal n12659 : std_logic;
signal n12660 : std_logic;
signal n12661 : std_logic;
signal n2315 : std_logic;
signal n2325 : std_logic;
signal n2195 : std_logic;
signal \bfn_5_20_0_\ : std_logic;
signal n12662 : std_logic;
signal n12663 : std_logic;
signal n12664 : std_logic;
signal n2297 : std_logic;
signal n12665 : std_logic;
signal n2296 : std_logic;
signal n12666 : std_logic;
signal n2295 : std_logic;
signal n12667 : std_logic;
signal n2294 : std_logic;
signal n12668 : std_logic;
signal n12669 : std_logic;
signal n2293 : std_logic;
signal \bfn_5_21_0_\ : std_logic;
signal n12670 : std_logic;
signal n12671 : std_logic;
signal n12672 : std_logic;
signal n12673 : std_logic;
signal n2288 : std_logic;
signal n12674 : std_logic;
signal n2287 : std_logic;
signal n12675 : std_logic;
signal n2286 : std_logic;
signal n12676 : std_logic;
signal n12677 : std_logic;
signal \bfn_5_22_0_\ : std_logic;
signal n12678 : std_logic;
signal n2283 : std_logic;
signal n12679 : std_logic;
signal n2282 : std_logic;
signal n12680 : std_logic;
signal n12681 : std_logic;
signal n2313 : std_logic;
signal n2299 : std_logic;
signal n2196 : std_logic;
signal n2198 : std_logic;
signal n2230 : std_logic;
signal \n2230_cascade_\ : std_logic;
signal n2289 : std_logic;
signal n2321 : std_logic;
signal n2331 : std_logic;
signal n11954 : std_logic;
signal n311 : std_logic;
signal n2533 : std_logic;
signal n2600 : std_logic;
signal n2532 : std_logic;
signal n2599 : std_logic;
signal n2631 : std_logic;
signal n2633 : std_logic;
signal \n2631_cascade_\ : std_logic;
signal n2632 : std_logic;
signal n12044 : std_logic;
signal n2301 : std_logic;
signal n2333 : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal n12878 : std_logic;
signal n12879 : std_logic;
signal n12880 : std_logic;
signal n12881 : std_logic;
signal n12882 : std_logic;
signal n12883 : std_logic;
signal n12884 : std_logic;
signal n12885 : std_logic;
signal \bfn_5_26_0_\ : std_logic;
signal n12886 : std_logic;
signal n12887 : std_logic;
signal n12888 : std_logic;
signal n12889 : std_logic;
signal n12890 : std_logic;
signal n12891 : std_logic;
signal n12892 : std_logic;
signal n12893 : std_logic;
signal \bfn_5_27_0_\ : std_logic;
signal n12894 : std_logic;
signal n12895 : std_logic;
signal n12896 : std_logic;
signal n12897 : std_logic;
signal n12898 : std_logic;
signal n12899 : std_logic;
signal n12900 : std_logic;
signal n12901 : std_logic;
signal \bfn_5_28_0_\ : std_logic;
signal n12902 : std_logic;
signal n12903 : std_logic;
signal n12904 : std_logic;
signal n12905 : std_logic;
signal n12906 : std_logic;
signal n3180 : std_logic;
signal n2925 : std_logic;
signal n2992 : std_logic;
signal n3099 : std_logic;
signal n3076 : std_logic;
signal n2926 : std_logic;
signal n2993 : std_logic;
signal n3027 : std_logic;
signal \n3025_cascade_\ : std_logic;
signal n14736 : std_logic;
signal n3014 : std_logic;
signal n3081 : std_logic;
signal n3100 : std_logic;
signal n3001 : std_logic;
signal n3033 : std_logic;
signal \n3033_cascade_\ : std_logic;
signal n3032 : std_logic;
signal n2990 : std_logic;
signal \n3022_cascade_\ : std_logic;
signal n14732 : std_logic;
signal n3030 : std_logic;
signal n3029 : std_logic;
signal n11932 : std_logic;
signal \n13859_cascade_\ : std_logic;
signal n14738 : std_logic;
signal n2999 : std_logic;
signal n2932 : std_logic;
signal n3031 : std_logic;
signal n3098 : std_logic;
signal \n3031_cascade_\ : std_logic;
signal n2916 : std_logic;
signal n2983 : std_logic;
signal n3015 : std_logic;
signal n3082 : std_logic;
signal \n3015_cascade_\ : std_logic;
signal n3089 : std_logic;
signal n3022 : std_logic;
signal n3095 : std_logic;
signal n3028 : std_logic;
signal \n3127_cascade_\ : std_logic;
signal n3011 : std_logic;
signal n14744 : std_logic;
signal n14816 : std_logic;
signal \n14750_cascade_\ : std_logic;
signal n3009 : std_logic;
signal n3007 : std_logic;
signal n3008 : std_logic;
signal \n14754_cascade_\ : std_logic;
signal n3006 : std_logic;
signal n3079 : std_logic;
signal \n3039_cascade_\ : std_logic;
signal n3012 : std_logic;
signal \n14194_cascade_\ : std_logic;
signal n14196 : std_logic;
signal n3018 : std_logic;
signal n3085 : std_logic;
signal \n3117_cascade_\ : std_logic;
signal n14198 : std_logic;
signal n3017 : std_logic;
signal n3084 : std_logic;
signal n3025 : std_logic;
signal n3092 : std_logic;
signal n3010 : std_logic;
signal n3077 : std_logic;
signal n2192 : std_logic;
signal n2291 : std_logic;
signal \n2224_cascade_\ : std_logic;
signal n2323 : std_logic;
signal n2193 : std_logic;
signal \n2126_cascade_\ : std_logic;
signal n2292 : std_logic;
signal \n2225_cascade_\ : std_logic;
signal n2324 : std_logic;
signal \n2116_cascade_\ : std_logic;
signal n2183 : std_logic;
signal \n2049_cascade_\ : std_logic;
signal n2186 : std_logic;
signal n2290 : std_logic;
signal n2322 : std_logic;
signal n2116 : std_logic;
signal \n2117_cascade_\ : std_logic;
signal \n2148_cascade_\ : std_logic;
signal n2197 : std_logic;
signal n2229 : std_logic;
signal n2189 : std_logic;
signal n2184 : std_logic;
signal n2117 : std_logic;
signal n2216 : std_logic;
signal n2215 : std_logic;
signal n2214 : std_logic;
signal \n2216_cascade_\ : std_logic;
signal n2298 : std_logic;
signal \n2247_cascade_\ : std_logic;
signal n2330 : std_logic;
signal n2187 : std_logic;
signal n2199 : std_logic;
signal n2285 : std_logic;
signal n2317 : std_logic;
signal n2200 : std_logic;
signal n2191 : std_logic;
signal n2185 : std_logic;
signal n2218 : std_logic;
signal n2219 : std_logic;
signal \n2217_cascade_\ : std_logic;
signal n14598 : std_logic;
signal n2188 : std_logic;
signal n2300 : std_logic;
signal n2332 : std_logic;
signal n2190 : std_logic;
signal n2228 : std_logic;
signal n2224 : std_logic;
signal n2227 : std_logic;
signal \n14578_cascade_\ : std_logic;
signal n2225 : std_logic;
signal n2223 : std_logic;
signal n2222 : std_logic;
signal \n14582_cascade_\ : std_logic;
signal n2221 : std_logic;
signal n2220 : std_logic;
signal \n14588_cascade_\ : std_logic;
signal n14812 : std_logic;
signal n14592 : std_logic;
signal n309 : std_logic;
signal \n17_adj_710_cascade_\ : std_logic;
signal \n19_adj_711_cascade_\ : std_logic;
signal n14236 : std_logic;
signal \n14230_cascade_\ : std_logic;
signal n61 : std_logic;
signal \n14268_cascade_\ : std_logic;
signal \n14806_cascade_\ : std_logic;
signal \n3237_cascade_\ : std_logic;
signal n14228 : std_logic;
signal n14270 : std_logic;
signal n14272 : std_logic;
signal n3173 : std_logic;
signal n3182 : std_logic;
signal \n3214_cascade_\ : std_logic;
signal n3190 : std_logic;
signal \n3222_cascade_\ : std_logic;
signal n27_adj_713 : std_logic;
signal n3183 : std_logic;
signal n3116 : std_logic;
signal n14794 : std_logic;
signal n14800 : std_logic;
signal n2891 : std_logic;
signal n2824 : std_logic;
signal n2923 : std_logic;
signal n3187 : std_logic;
signal n3189 : std_logic;
signal \n3221_cascade_\ : std_logic;
signal n3175 : std_logic;
signal n3121 : std_logic;
signal n3188 : std_logic;
signal n3191 : std_logic;
signal n3124 : std_logic;
signal n3179 : std_logic;
signal n3113 : std_logic;
signal n3108 : std_logic;
signal \n14216_cascade_\ : std_logic;
signal n3105 : std_logic;
signal \n14222_cascade_\ : std_logic;
signal n3106 : std_logic;
signal \n3138_cascade_\ : std_logic;
signal n3107 : std_logic;
signal n3174 : std_logic;
signal n3201 : std_logic;
signal n11861 : std_logic;
signal \n3233_cascade_\ : std_logic;
signal n3111 : std_logic;
signal n3178 : std_logic;
signal n3023 : std_logic;
signal n3090 : std_logic;
signal n3122 : std_logic;
signal n3181 : std_logic;
signal n3199 : std_logic;
signal n3198 : std_logic;
signal n3115 : std_logic;
signal n3114 : std_logic;
signal n14204 : std_logic;
signal n14210 : std_logic;
signal n3101 : std_logic;
signal n3200 : std_logic;
signal \n3133_cascade_\ : std_logic;
signal \n3232_cascade_\ : std_logic;
signal \n25_adj_712_cascade_\ : std_logic;
signal n37_adj_715 : std_logic;
signal n14234 : std_logic;
signal \n14238_cascade_\ : std_logic;
signal n14248 : std_logic;
signal \n14250_cascade_\ : std_logic;
signal n3026 : std_logic;
signal n3093 : std_logic;
signal n59 : std_logic;
signal n14252 : std_logic;
signal n5_adj_703 : std_logic;
signal \n14254_cascade_\ : std_logic;
signal n11926 : std_logic;
signal \n14256_cascade_\ : std_logic;
signal n7_adj_708 : std_logic;
signal \n14264_cascade_\ : std_logic;
signal n14266 : std_logic;
signal n14258 : std_logic;
signal \n14260_cascade_\ : std_logic;
signal n14262 : std_logic;
signal n3021 : std_logic;
signal n3088 : std_logic;
signal n3120 : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal n12625 : std_logic;
signal n2099 : std_logic;
signal n12626 : std_logic;
signal n12627 : std_logic;
signal n2097 : std_logic;
signal n12628 : std_logic;
signal n2096 : std_logic;
signal n12629 : std_logic;
signal n12630 : std_logic;
signal n2094 : std_logic;
signal n12631 : std_logic;
signal n12632 : std_logic;
signal n2093 : std_logic;
signal \bfn_7_18_0_\ : std_logic;
signal n12633 : std_logic;
signal n2091 : std_logic;
signal n12634 : std_logic;
signal n12635 : std_logic;
signal n12636 : std_logic;
signal n2088 : std_logic;
signal n12637 : std_logic;
signal n2087 : std_logic;
signal n12638 : std_logic;
signal n12639 : std_logic;
signal n12640 : std_logic;
signal n2085 : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal n2084 : std_logic;
signal n12641 : std_logic;
signal n12642 : std_logic;
signal n2115 : std_logic;
signal n2095 : std_logic;
signal n2123 : std_logic;
signal \n2127_cascade_\ : std_logic;
signal n2126 : std_logic;
signal n2018 : std_logic;
signal n2092 : std_logic;
signal n2124 : std_logic;
signal n2098 : std_logic;
signal n2130 : std_logic;
signal n2131 : std_logic;
signal n2129 : std_logic;
signal \n2130_cascade_\ : std_logic;
signal n2119 : std_logic;
signal \n13775_cascade_\ : std_logic;
signal n14398 : std_logic;
signal n2090 : std_logic;
signal n2122 : std_logic;
signal n2125 : std_logic;
signal \n2122_cascade_\ : std_logic;
signal n2128 : std_logic;
signal n2120 : std_logic;
signal \n14386_cascade_\ : std_logic;
signal n14384 : std_logic;
signal n14392 : std_logic;
signal n2089 : std_logic;
signal n2121 : std_logic;
signal n2127 : std_logic;
signal n2194 : std_logic;
signal n2226 : std_logic;
signal n2101 : std_logic;
signal n2133 : std_logic;
signal \n2133_cascade_\ : std_logic;
signal n11892 : std_logic;
signal n307 : std_logic;
signal n2201 : std_logic;
signal n2233 : std_logic;
signal n2231 : std_logic;
signal \n2233_cascade_\ : std_logic;
signal n2232 : std_logic;
signal n11950 : std_logic;
signal n2086 : std_logic;
signal n2118 : std_logic;
signal n308 : std_logic;
signal n2284 : std_logic;
signal n2217 : std_logic;
signal n2316 : std_logic;
signal n2100 : std_logic;
signal n2132 : std_logic;
signal n315 : std_logic;
signal n15484 : std_logic;
signal n12034 : std_logic;
signal \bfn_7_23_0_\ : std_logic;
signal n12938 : std_logic;
signal n15445 : std_logic;
signal n12939 : std_logic;
signal n15412 : std_logic;
signal n12940 : std_logic;
signal n15378 : std_logic;
signal n2940 : std_logic;
signal n12941 : std_logic;
signal n15346 : std_logic;
signal n2841 : std_logic;
signal n12942 : std_logic;
signal n15310 : std_logic;
signal n2742 : std_logic;
signal n12943 : std_logic;
signal n15852 : std_logic;
signal n2643 : std_logic;
signal n12944 : std_logic;
signal n12945 : std_logic;
signal n15821 : std_logic;
signal n2544 : std_logic;
signal \bfn_7_24_0_\ : std_logic;
signal n15791 : std_logic;
signal n2445 : std_logic;
signal n12946 : std_logic;
signal n15765 : std_logic;
signal n2346 : std_logic;
signal n12947 : std_logic;
signal n15739 : std_logic;
signal n2247 : std_logic;
signal n12948 : std_logic;
signal n15714 : std_logic;
signal n2148 : std_logic;
signal n12949 : std_logic;
signal n15689 : std_logic;
signal n2049 : std_logic;
signal n12950 : std_logic;
signal n12951 : std_logic;
signal n12952 : std_logic;
signal n12953 : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal n12954 : std_logic;
signal n12955 : std_logic;
signal n12956 : std_logic;
signal n12957 : std_logic;
signal n12958 : std_logic;
signal n12959 : std_logic;
signal n12960 : std_logic;
signal n3177 : std_logic;
signal n3110 : std_logic;
signal \n31_adj_714_cascade_\ : std_logic;
signal n14232 : std_logic;
signal n3126 : std_logic;
signal n3193 : std_logic;
signal \n3225_cascade_\ : std_logic;
signal \n14776_cascade_\ : std_logic;
signal n14764 : std_logic;
signal \n14780_cascade_\ : std_logic;
signal n3128 : std_logic;
signal n3195 : std_logic;
signal n3117 : std_logic;
signal n3184 : std_logic;
signal n3119 : std_logic;
signal n3186 : std_logic;
signal \n3218_cascade_\ : std_logic;
signal n14778 : std_logic;
signal n12030 : std_logic;
signal n14786 : std_logic;
signal n14788 : std_logic;
signal encoder0_position_scaled_12 : std_logic;
signal n3194 : std_logic;
signal n3127 : std_logic;
signal n3013 : std_logic;
signal n3080 : std_logic;
signal n3112 : std_logic;
signal n3192 : std_logic;
signal n3125 : std_logic;
signal n3196 : std_logic;
signal \debounce.reg_A_0\ : std_logic;
signal \reg_B_0\ : std_logic;
signal \debounce.reg_A_1\ : std_logic;
signal \debounce.n6\ : std_logic;
signal n3185 : std_logic;
signal n3118 : std_logic;
signal n3197 : std_logic;
signal \n3229_cascade_\ : std_logic;
signal n3237 : std_logic;
signal n13_adj_709 : std_logic;
signal n319 : std_logic;
signal \bfn_7_29_0_\ : std_logic;
signal n3301 : std_logic;
signal n12907 : std_logic;
signal n3233 : std_logic;
signal n3300 : std_logic;
signal n12908 : std_logic;
signal n3232 : std_logic;
signal n3299 : std_logic;
signal n12909 : std_logic;
signal n3231 : std_logic;
signal n12910 : std_logic;
signal n3298 : std_logic;
signal n3230 : std_logic;
signal n15097 : std_logic;
signal n12911 : std_logic;
signal n3229 : std_logic;
signal n3296 : std_logic;
signal n12912 : std_logic;
signal n3228 : std_logic;
signal n3295 : std_logic;
signal n12913 : std_logic;
signal n12914 : std_logic;
signal n3227 : std_logic;
signal n3294 : std_logic;
signal \bfn_7_30_0_\ : std_logic;
signal n3226 : std_logic;
signal n3293 : std_logic;
signal n12915 : std_logic;
signal n3225 : std_logic;
signal n3292 : std_logic;
signal n12916 : std_logic;
signal n3224 : std_logic;
signal n3291 : std_logic;
signal n12917 : std_logic;
signal n3223 : std_logic;
signal n3290 : std_logic;
signal n12918 : std_logic;
signal n3222 : std_logic;
signal n3289 : std_logic;
signal n12919 : std_logic;
signal n3221 : std_logic;
signal n3288 : std_logic;
signal n12920 : std_logic;
signal n3220 : std_logic;
signal n3287 : std_logic;
signal n12921 : std_logic;
signal n12922 : std_logic;
signal n3219 : std_logic;
signal n3286 : std_logic;
signal \bfn_7_31_0_\ : std_logic;
signal n3218 : std_logic;
signal n3285 : std_logic;
signal n12923 : std_logic;
signal n3217 : std_logic;
signal n3284 : std_logic;
signal n12924 : std_logic;
signal n3216 : std_logic;
signal n3283 : std_logic;
signal n12925 : std_logic;
signal n3215 : std_logic;
signal n3282 : std_logic;
signal n12926 : std_logic;
signal n3214 : std_logic;
signal n3281 : std_logic;
signal n12927 : std_logic;
signal n3213 : std_logic;
signal n3280 : std_logic;
signal n12928 : std_logic;
signal n3212 : std_logic;
signal n3279 : std_logic;
signal n12929 : std_logic;
signal n12930 : std_logic;
signal n3211 : std_logic;
signal n3278 : std_logic;
signal \bfn_7_32_0_\ : std_logic;
signal n3210 : std_logic;
signal n3277 : std_logic;
signal n12931 : std_logic;
signal n3209 : std_logic;
signal n3276 : std_logic;
signal n12932 : std_logic;
signal n3275 : std_logic;
signal n12933 : std_logic;
signal n3207 : std_logic;
signal n3274 : std_logic;
signal n12934 : std_logic;
signal n3206 : std_logic;
signal n3273 : std_logic;
signal n12935 : std_logic;
signal n3205 : std_logic;
signal n3272 : std_logic;
signal n12936 : std_logic;
signal n15450 : std_logic;
signal n3204 : std_logic;
signal n12937 : std_logic;
signal n14873 : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal n12608 : std_logic;
signal n12609 : std_logic;
signal n12610 : std_logic;
signal n12611 : std_logic;
signal n12612 : std_logic;
signal n12613 : std_logic;
signal n12614 : std_logic;
signal n12615 : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal n12616 : std_logic;
signal n12617 : std_logic;
signal n12618 : std_logic;
signal n12619 : std_logic;
signal n12620 : std_logic;
signal n12621 : std_logic;
signal n1986 : std_logic;
signal n12622 : std_logic;
signal n12623 : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal n12624 : std_logic;
signal n2016 : std_logic;
signal n1993 : std_logic;
signal n1990 : std_logic;
signal n1985 : std_logic;
signal n2017 : std_logic;
signal n1992 : std_logic;
signal n1997 : std_logic;
signal n1987 : std_logic;
signal n2025 : std_logic;
signal n2022 : std_logic;
signal n2024 : std_logic;
signal \n14550_cascade_\ : std_logic;
signal n2029 : std_logic;
signal \n14556_cascade_\ : std_logic;
signal \n14558_cascade_\ : std_logic;
signal n2019 : std_logic;
signal n14564 : std_logic;
signal n1991 : std_logic;
signal n2023 : std_logic;
signal n1994 : std_logic;
signal n2026 : std_logic;
signal encoder0_position_0 : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \quad_counter0.n13025\ : std_logic;
signal \quad_counter0.n13026\ : std_logic;
signal \quad_counter0.n13027\ : std_logic;
signal encoder0_position_4 : std_logic;
signal \quad_counter0.n13028\ : std_logic;
signal \quad_counter0.n13029\ : std_logic;
signal \quad_counter0.n13030\ : std_logic;
signal \quad_counter0.n13031\ : std_logic;
signal \quad_counter0.n13032\ : std_logic;
signal encoder0_position_8 : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \quad_counter0.n13033\ : std_logic;
signal \quad_counter0.n13034\ : std_logic;
signal encoder0_position_11 : std_logic;
signal \quad_counter0.n13035\ : std_logic;
signal encoder0_position_12 : std_logic;
signal \quad_counter0.n13036\ : std_logic;
signal encoder0_position_13 : std_logic;
signal \quad_counter0.n13037\ : std_logic;
signal \quad_counter0.n13038\ : std_logic;
signal \quad_counter0.n13039\ : std_logic;
signal \quad_counter0.n13040\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \quad_counter0.n13041\ : std_logic;
signal \quad_counter0.n13042\ : std_logic;
signal \quad_counter0.n13043\ : std_logic;
signal \quad_counter0.n13044\ : std_logic;
signal \quad_counter0.n13045\ : std_logic;
signal \quad_counter0.n13046\ : std_logic;
signal \quad_counter0.n13047\ : std_logic;
signal \quad_counter0.n13048\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \quad_counter0.n13049\ : std_logic;
signal \quad_counter0.n13050\ : std_logic;
signal \quad_counter0.n13051\ : std_logic;
signal \quad_counter0.n13052\ : std_logic;
signal \quad_counter0.n13053\ : std_logic;
signal \quad_counter0.n13054\ : std_logic;
signal \quad_counter0.n13055\ : std_logic;
signal encoder0_position_scaled_17 : std_logic;
signal encoder0_position_14 : std_logic;
signal encoder0_position_scaled_4 : std_logic;
signal encoder0_position_scaled_5 : std_logic;
signal encoder0_position_scaled_22 : std_logic;
signal n3133 : std_logic;
signal n3132 : std_logic;
signal n3129 : std_logic;
signal n3130 : std_logic;
signal \n11930_cascade_\ : std_logic;
signal n3131 : std_logic;
signal n13819 : std_logic;
signal \quad_counter0.a_prev_N_543_cascade_\ : std_logic;
signal \quad_counter0.direction_N_536\ : std_logic;
signal n3024 : std_logic;
signal n3091 : std_logic;
signal n3039 : std_logic;
signal n3123 : std_logic;
signal \ENCODER0_A_N\ : std_logic;
signal \quad_counter0.a_new_0\ : std_logic;
signal encoder0_position_scaled_21 : std_logic;
signal encoder0_position_scaled_19 : std_logic;
signal n25_adj_605 : std_logic;
signal \pwm_setpoint_23_N_171_0\ : std_logic;
signal \bfn_9_30_0_\ : std_logic;
signal n24_adj_604 : std_logic;
signal \pwm_setpoint_23_N_171_1\ : std_logic;
signal n12412 : std_logic;
signal n23_adj_603 : std_logic;
signal n12413 : std_logic;
signal n22_adj_602 : std_logic;
signal n12414 : std_logic;
signal n12415 : std_logic;
signal n12416 : std_logic;
signal n12417 : std_logic;
signal n18_adj_598 : std_logic;
signal n12418 : std_logic;
signal n12419 : std_logic;
signal n17_adj_597 : std_logic;
signal \bfn_9_31_0_\ : std_logic;
signal n12420 : std_logic;
signal n12421 : std_logic;
signal n14_adj_594 : std_logic;
signal n12422 : std_logic;
signal n13_adj_593 : std_logic;
signal n12423 : std_logic;
signal n12424 : std_logic;
signal n12425 : std_logic;
signal n10_adj_590 : std_logic;
signal n12426 : std_logic;
signal n12427 : std_logic;
signal \bfn_9_32_0_\ : std_logic;
signal n12428 : std_logic;
signal n12429 : std_logic;
signal n6_adj_586 : std_logic;
signal n12430 : std_logic;
signal n12431 : std_logic;
signal n12432 : std_logic;
signal n12433 : std_logic;
signal n12434 : std_logic;
signal encoder0_position_9 : std_logic;
signal n310 : std_logic;
signal n1927 : std_logic;
signal n1923 : std_logic;
signal n1926 : std_logic;
signal \n1923_cascade_\ : std_logic;
signal n1924 : std_logic;
signal n14408 : std_logic;
signal \n1921_cascade_\ : std_logic;
signal n14410 : std_logic;
signal n1995 : std_logic;
signal n2027 : std_logic;
signal n1925 : std_logic;
signal n1922 : std_logic;
signal n1989 : std_logic;
signal \n1922_cascade_\ : std_logic;
signal n2021 : std_logic;
signal n14416 : std_logic;
signal \n14420_cascade_\ : std_logic;
signal \n1950_cascade_\ : std_logic;
signal n1998 : std_logic;
signal n2030 : std_logic;
signal n15666 : std_logic;
signal n1917 : std_logic;
signal n1988 : std_logic;
signal n1921 : std_logic;
signal n2020 : std_logic;
signal n11966 : std_logic;
signal n1932 : std_logic;
signal \n1932_cascade_\ : std_logic;
signal n1999 : std_logic;
signal n2031 : std_logic;
signal n306 : std_logic;
signal \n2031_cascade_\ : std_logic;
signal n11964 : std_logic;
signal n305 : std_logic;
signal n2001 : std_logic;
signal n2033 : std_logic;
signal n1996 : std_logic;
signal n2028 : std_logic;
signal n2000 : std_logic;
signal n1933 : std_logic;
signal n1950 : std_logic;
signal n2032 : std_logic;
signal n33_adj_654 : std_logic;
signal n33 : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal n32_adj_653 : std_logic;
signal n12968 : std_logic;
signal n31_adj_652 : std_logic;
signal n12969 : std_logic;
signal n12970 : std_logic;
signal n29_adj_650 : std_logic;
signal n29 : std_logic;
signal n12971 : std_logic;
signal n28_adj_649 : std_logic;
signal n12972 : std_logic;
signal n27_adj_648 : std_logic;
signal n12973 : std_logic;
signal n26_adj_647 : std_logic;
signal n12974 : std_logic;
signal n12975 : std_logic;
signal n25_adj_646 : std_logic;
signal n25_adj_551 : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal n24_adj_645 : std_logic;
signal n24 : std_logic;
signal n12976 : std_logic;
signal n23 : std_logic;
signal n12977 : std_logic;
signal n22_adj_643 : std_logic;
signal n22 : std_logic;
signal n12978 : std_logic;
signal n21_adj_642 : std_logic;
signal n21 : std_logic;
signal n12979 : std_logic;
signal n20_adj_641 : std_logic;
signal n20 : std_logic;
signal n12980 : std_logic;
signal n19_adj_640 : std_logic;
signal n19 : std_logic;
signal n12981 : std_logic;
signal n12982 : std_logic;
signal n12983 : std_logic;
signal n17_adj_638 : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal n12984 : std_logic;
signal n15_adj_636 : std_logic;
signal n12985 : std_logic;
signal n12986 : std_logic;
signal n13_adj_634 : std_logic;
signal n12987 : std_logic;
signal n12988 : std_logic;
signal n12989 : std_logic;
signal n12990 : std_logic;
signal n12991 : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal n12992 : std_logic;
signal n12993 : std_logic;
signal n12994 : std_logic;
signal n12995 : std_logic;
signal n12996 : std_logic;
signal n12997 : std_logic;
signal n12998 : std_logic;
signal n5_adj_626 : std_logic;
signal n6_adj_627 : std_logic;
signal n8_adj_629 : std_logic;
signal n7_adj_628 : std_logic;
signal n4_adj_625 : std_logic;
signal pwm_setpoint_1 : std_logic;
signal pwm_setpoint_0 : std_logic;
signal n28 : std_logic;
signal encoder0_position_5 : std_logic;
signal n314 : std_logic;
signal \quad_counter0.b_new_0\ : std_logic;
signal encoder0_position_scaled_0 : std_logic;
signal encoder0_position_scaled_15 : std_logic;
signal encoder0_position_scaled_13 : std_logic;
signal n3_adj_624 : std_logic;
signal encoder0_position_scaled_2 : std_logic;
signal n4_adj_655 : std_logic;
signal \quad_counter0.a_prev_N_543\ : std_logic;
signal \quad_counter0.b_new_1\ : std_logic;
signal \quad_counter0.a_prev\ : std_logic;
signal \quad_counter0.debounce_cnt\ : std_logic;
signal \quad_counter0.direction_N_540_cascade_\ : std_logic;
signal \direction_N_537\ : std_logic;
signal a_new_1 : std_logic;
signal \direction_N_537_cascade_\ : std_logic;
signal b_prev : std_logic;
signal n1302 : std_logic;
signal \n29_adj_672_cascade_\ : std_logic;
signal n15233 : std_logic;
signal n15234 : std_logic;
signal encoder0_position_scaled_16 : std_logic;
signal \n33_adj_675_cascade_\ : std_logic;
signal n12_adj_592 : std_logic;
signal \pwm_setpoint_23_N_171_16\ : std_logic;
signal \pwm_setpoint_23_N_171_2\ : std_logic;
signal \pwm_setpoint_23_N_171_14\ : std_logic;
signal pwm_setpoint_14 : std_logic;
signal n15121 : std_logic;
signal n15182 : std_logic;
signal n29_adj_672 : std_logic;
signal \n30_adj_673_cascade_\ : std_logic;
signal n10_adj_659 : std_logic;
signal n15267 : std_logic;
signal n20_adj_600 : std_logic;
signal n16_adj_596 : std_logic;
signal n15_adj_595 : std_logic;
signal n21_adj_601 : std_logic;
signal \pwm_setpoint_23_N_171_5\ : std_logic;
signal n19_adj_599 : std_logic;
signal \pwm_setpoint_23_N_171_6\ : std_logic;
signal \pwm_setpoint_23_N_171_10\ : std_logic;
signal \pwm_setpoint_23_N_171_9\ : std_logic;
signal \pwm_setpoint_23_N_171_4\ : std_logic;
signal n7_adj_587 : std_logic;
signal \pwm_setpoint_23_N_171_15\ : std_logic;
signal \reg_B_1\ : std_logic;
signal pwm_setpoint_15 : std_logic;
signal n31_adj_674 : std_logic;
signal n11_adj_591 : std_logic;
signal \pwm_setpoint_23_N_171_18\ : std_logic;
signal n3_adj_583 : std_logic;
signal n9_adj_589 : std_logic;
signal \reg_B_2\ : std_logic;
signal n14125 : std_logic;
signal n14937 : std_logic;
signal \n14936_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal \pwm_setpoint_23_N_171_22\ : std_logic;
signal \n1826_cascade_\ : std_logic;
signal n1928 : std_logic;
signal n14526 : std_logic;
signal \n14530_cascade_\ : std_logic;
signal \n1819_cascade_\ : std_logic;
signal n14532 : std_logic;
signal \n1851_cascade_\ : std_logic;
signal n1920 : std_logic;
signal n1919 : std_logic;
signal n1930 : std_logic;
signal \n1930_cascade_\ : std_logic;
signal n1929 : std_logic;
signal n14540 : std_logic;
signal n1931 : std_logic;
signal n1918 : std_logic;
signal n14520 : std_logic;
signal \n14176_cascade_\ : std_logic;
signal \n1752_cascade_\ : std_logic;
signal n1851 : std_logic;
signal n15644 : std_logic;
signal \n1832_cascade_\ : std_logic;
signal n11968 : std_logic;
signal \n1820_cascade_\ : std_logic;
signal n14538 : std_logic;
signal n30_adj_651 : std_logic;
signal n26 : std_logic;
signal encoder0_position_7 : std_logic;
signal n312 : std_logic;
signal n31 : std_logic;
signal encoder0_position_2 : std_logic;
signal n317 : std_logic;
signal encoder0_position_10 : std_logic;
signal n23_adj_644 : std_logic;
signal encoder0_position_scaled_1 : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal n12487 : std_logic;
signal n12488 : std_logic;
signal n12489 : std_logic;
signal n12490 : std_logic;
signal n12491 : std_logic;
signal n12492 : std_logic;
signal n901 : std_logic;
signal n896 : std_logic;
signal n900 : std_logic;
signal n899 : std_logic;
signal \n931_cascade_\ : std_logic;
signal n10 : std_logic;
signal n897 : std_logic;
signal encoder0_position_25 : std_logic;
signal n8 : std_logic;
signal n294 : std_logic;
signal n14574 : std_logic;
signal n828 : std_logic;
signal \n828_cascade_\ : std_logic;
signal n12012 : std_logic;
signal n861 : std_logic;
signal \n861_cascade_\ : std_logic;
signal n898 : std_logic;
signal \n13644_cascade_\ : std_logic;
signal n830 : std_logic;
signal n7 : std_logic;
signal n5_adj_676 : std_logic;
signal \n5_adj_676_cascade_\ : std_logic;
signal \n13641_cascade_\ : std_logic;
signal \n13646_cascade_\ : std_logic;
signal n831 : std_logic;
signal encoder0_position_28 : std_logic;
signal n5 : std_logic;
signal encoder0_position_29 : std_logic;
signal n4 : std_logic;
signal n3 : std_logic;
signal encoder0_position_30 : std_logic;
signal \n13642_cascade_\ : std_logic;
signal n829 : std_logic;
signal n32 : std_logic;
signal encoder0_position_1 : std_logic;
signal n318 : std_logic;
signal encoder0_position_scaled_14 : std_logic;
signal \n10_adj_606_cascade_\ : std_logic;
signal \n15_adj_565_cascade_\ : std_logic;
signal n16_adj_564 : std_logic;
signal encoder0_position_scaled_10 : std_logic;
signal \pwm_setpoint_23_N_171_3\ : std_logic;
signal encoder0_position_scaled_11 : std_logic;
signal \pwm_setpoint_23_N_171_13\ : std_logic;
signal \n15_adj_663_cascade_\ : std_logic;
signal n15125 : std_logic;
signal encoder0_position_scaled_18 : std_logic;
signal encoder0_position_scaled_20 : std_logic;
signal encoder0_position_scaled_23 : std_logic;
signal n12_adj_661 : std_logic;
signal \pwm_setpoint_23_N_171_7\ : std_logic;
signal pwm_setpoint_16 : std_logic;
signal pwm_setpoint_7 : std_logic;
signal n15119 : std_logic;
signal encoder0_position_scaled_9 : std_logic;
signal n26_adj_697 : std_logic;
signal \bfn_11_29_0_\ : std_logic;
signal n25_adj_696 : std_logic;
signal n13087 : std_logic;
signal n24_adj_695 : std_logic;
signal n13088 : std_logic;
signal n23_adj_694 : std_logic;
signal n13089 : std_logic;
signal n22_adj_693 : std_logic;
signal n13090 : std_logic;
signal n21_adj_692 : std_logic;
signal n13091 : std_logic;
signal n20_adj_691 : std_logic;
signal n13092 : std_logic;
signal n19_adj_690 : std_logic;
signal n13093 : std_logic;
signal n13094 : std_logic;
signal n18_adj_689 : std_logic;
signal \bfn_11_30_0_\ : std_logic;
signal n17_adj_688 : std_logic;
signal n13095 : std_logic;
signal n16_adj_687 : std_logic;
signal n13096 : std_logic;
signal n15_adj_686 : std_logic;
signal n13097 : std_logic;
signal n14_adj_685 : std_logic;
signal n13098 : std_logic;
signal n13_adj_684 : std_logic;
signal n13099 : std_logic;
signal n12_adj_683 : std_logic;
signal n13100 : std_logic;
signal n11_adj_682 : std_logic;
signal n13101 : std_logic;
signal n13102 : std_logic;
signal n10_adj_681 : std_logic;
signal \bfn_11_31_0_\ : std_logic;
signal n9_adj_680 : std_logic;
signal n13103 : std_logic;
signal n8_adj_679 : std_logic;
signal n13104 : std_logic;
signal n7_adj_678 : std_logic;
signal n13105 : std_logic;
signal n6_adj_677 : std_logic;
signal n13106 : std_logic;
signal blink_counter_21 : std_logic;
signal n13107 : std_logic;
signal blink_counter_22 : std_logic;
signal n13108 : std_logic;
signal blink_counter_23 : std_logic;
signal n13109 : std_logic;
signal n13110 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_11_32_0_\ : std_logic;
signal n13111 : std_logic;
signal blink_counter_25 : std_logic;
signal \pwm_setpoint_23_N_171_19\ : std_logic;
signal n8_adj_588 : std_logic;
signal n5_adj_585 : std_logic;
signal n1901 : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal n1833 : std_logic;
signal n1900 : std_logic;
signal n12592 : std_logic;
signal n1832 : std_logic;
signal n1899 : std_logic;
signal n12593 : std_logic;
signal n1831 : std_logic;
signal n1898 : std_logic;
signal n12594 : std_logic;
signal n1830 : std_logic;
signal n1897 : std_logic;
signal n12595 : std_logic;
signal n1829 : std_logic;
signal n1896 : std_logic;
signal n12596 : std_logic;
signal n1828 : std_logic;
signal n1895 : std_logic;
signal n12597 : std_logic;
signal n1894 : std_logic;
signal n12598 : std_logic;
signal n12599 : std_logic;
signal n1826 : std_logic;
signal n1893 : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal n1825 : std_logic;
signal n1892 : std_logic;
signal n12600 : std_logic;
signal n1824 : std_logic;
signal n1891 : std_logic;
signal n12601 : std_logic;
signal n1823 : std_logic;
signal n1890 : std_logic;
signal n12602 : std_logic;
signal n1822 : std_logic;
signal n1889 : std_logic;
signal n12603 : std_logic;
signal n1888 : std_logic;
signal n12604 : std_logic;
signal n1820 : std_logic;
signal n1887 : std_logic;
signal n12605 : std_logic;
signal n1819 : std_logic;
signal n1886 : std_logic;
signal n12606 : std_logic;
signal n12607 : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal n1885 : std_logic;
signal \n1722_cascade_\ : std_logic;
signal n1821 : std_logic;
signal n1827 : std_logic;
signal n1752 : std_logic;
signal n16_adj_637 : std_logic;
signal n2 : std_logic;
signal n16 : std_logic;
signal encoder0_position_17 : std_logic;
signal n30 : std_logic;
signal encoder0_position_3 : std_logic;
signal n316 : std_logic;
signal n2_adj_623 : std_logic;
signal encoder0_position_scaled_7 : std_logic;
signal encoder0_position_23 : std_logic;
signal n10_adj_631 : std_logic;
signal n18_adj_639 : std_logic;
signal n17 : std_logic;
signal encoder0_position_16 : std_logic;
signal n18 : std_logic;
signal encoder0_position_15 : std_logic;
signal n304 : std_logic;
signal n15 : std_logic;
signal encoder0_position_18 : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal n12493 : std_logic;
signal n12494 : std_logic;
signal n12495 : std_logic;
signal n12496 : std_logic;
signal n12497 : std_logic;
signal n12498 : std_logic;
signal n12499 : std_logic;
signal n1001 : std_logic;
signal n927 : std_logic;
signal \n14466_cascade_\ : std_logic;
signal n11940 : std_logic;
signal n930 : std_logic;
signal \n960_cascade_\ : std_logic;
signal n997 : std_logic;
signal n929 : std_logic;
signal n996 : std_logic;
signal \n1028_cascade_\ : std_logic;
signal n998 : std_logic;
signal n931 : std_logic;
signal encoder0_position_scaled_8 : std_logic;
signal n6 : std_logic;
signal n13641 : std_logic;
signal \n13648_cascade_\ : std_logic;
signal encoder0_position_27 : std_logic;
signal n832 : std_logic;
signal n999 : std_logic;
signal n932 : std_logic;
signal encoder0_position_26 : std_logic;
signal n13650 : std_logic;
signal n833 : std_logic;
signal encoder0_position_scaled_3 : std_logic;
signal n293 : std_logic;
signal n2542 : std_logic;
signal \bfn_12_25_0_\ : std_logic;
signal n292 : std_logic;
signal n2541 : std_logic;
signal n12482 : std_logic;
signal n174 : std_logic;
signal n2540 : std_logic;
signal n12483 : std_logic;
signal n404 : std_logic;
signal n2539 : std_logic;
signal n12484 : std_logic;
signal n403 : std_logic;
signal n2538 : std_logic;
signal n12485 : std_logic;
signal n402 : std_logic;
signal n12486 : std_logic;
signal n2537 : std_logic;
signal encoder0_position_scaled_6 : std_logic;
signal n3109 : std_logic;
signal n3176 : std_logic;
signal n3138 : std_logic;
signal n3208 : std_logic;
signal n25_adj_552 : std_logic;
signal duty_0 : std_logic;
signal \bfn_12_26_0_\ : std_logic;
signal n24_adj_553 : std_logic;
signal duty_1 : std_logic;
signal n12459 : std_logic;
signal n23_adj_554 : std_logic;
signal duty_2 : std_logic;
signal n12460 : std_logic;
signal n22_adj_555 : std_logic;
signal duty_3 : std_logic;
signal n12461 : std_logic;
signal n21_adj_556 : std_logic;
signal duty_4 : std_logic;
signal n12462 : std_logic;
signal n20_adj_557 : std_logic;
signal duty_5 : std_logic;
signal n12463 : std_logic;
signal n19_adj_558 : std_logic;
signal duty_6 : std_logic;
signal n12464 : std_logic;
signal n18_adj_559 : std_logic;
signal duty_7 : std_logic;
signal n12465 : std_logic;
signal n12466 : std_logic;
signal n17_adj_560 : std_logic;
signal \bfn_12_27_0_\ : std_logic;
signal n16_adj_563 : std_logic;
signal duty_9 : std_logic;
signal n12467 : std_logic;
signal n15_adj_568 : std_logic;
signal duty_10 : std_logic;
signal n12468 : std_logic;
signal n14_adj_569 : std_logic;
signal n12469 : std_logic;
signal n13_adj_570 : std_logic;
signal n12470 : std_logic;
signal n12_adj_571 : std_logic;
signal duty_13 : std_logic;
signal n12471 : std_logic;
signal n11_adj_572 : std_logic;
signal duty_14 : std_logic;
signal n12472 : std_logic;
signal n10_adj_573 : std_logic;
signal duty_15 : std_logic;
signal n12473 : std_logic;
signal n12474 : std_logic;
signal n9_adj_574 : std_logic;
signal duty_16 : std_logic;
signal \bfn_12_28_0_\ : std_logic;
signal n8_adj_575 : std_logic;
signal n12475 : std_logic;
signal n7_adj_576 : std_logic;
signal duty_18 : std_logic;
signal n12476 : std_logic;
signal n6_adj_577 : std_logic;
signal duty_19 : std_logic;
signal n12477 : std_logic;
signal n5_adj_578 : std_logic;
signal n12478 : std_logic;
signal n4_adj_579 : std_logic;
signal n12479 : std_logic;
signal n3_adj_580 : std_logic;
signal duty_22 : std_logic;
signal n12480 : std_logic;
signal n2_adj_581 : std_logic;
signal n12481 : std_logic;
signal n35 : std_logic;
signal n33_adj_675 : std_logic;
signal \n35_cascade_\ : std_logic;
signal n15225 : std_logic;
signal pwm_setpoint_13 : std_logic;
signal n27_adj_671 : std_logic;
signal duty_12 : std_logic;
signal \pwm_setpoint_23_N_171_12\ : std_logic;
signal n37 : std_logic;
signal pwm_setpoint_18 : std_logic;
signal n15277 : std_logic;
signal n6_adj_656 : std_logic;
signal \n15235_cascade_\ : std_logic;
signal \n15236_cascade_\ : std_logic;
signal duty_11 : std_logic;
signal \pwm_setpoint_23_N_171_11\ : std_logic;
signal duty_17 : std_logic;
signal \pwm_setpoint_23_N_171_17\ : std_logic;
signal pwm_setpoint_17 : std_logic;
signal n15278 : std_logic;
signal \n8_adj_657_cascade_\ : std_logic;
signal n15180 : std_logic;
signal \n15219_cascade_\ : std_logic;
signal n24_adj_669 : std_logic;
signal pwm_setpoint_22 : std_logic;
signal n15274 : std_logic;
signal n45 : std_logic;
signal n15255 : std_logic;
signal \n40_cascade_\ : std_logic;
signal duty_20 : std_logic;
signal \pwm_setpoint_23_N_171_20\ : std_logic;
signal n4_adj_584 : std_logic;
signal n16_adj_664 : std_logic;
signal \pwm_setpoint_23__N_195\ : std_logic;
signal \pwm_setpoint_23_N_171_21\ : std_logic;
signal duty_21 : std_logic;
signal n1801 : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal n1800 : std_logic;
signal n12577 : std_logic;
signal n1799 : std_logic;
signal n12578 : std_logic;
signal n1798 : std_logic;
signal n12579 : std_logic;
signal n1797 : std_logic;
signal n12580 : std_logic;
signal n1796 : std_logic;
signal n12581 : std_logic;
signal n1795 : std_logic;
signal n12582 : std_logic;
signal n1794 : std_logic;
signal n12583 : std_logic;
signal n12584 : std_logic;
signal n1793 : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal n1792 : std_logic;
signal n12585 : std_logic;
signal n1791 : std_logic;
signal n12586 : std_logic;
signal n1790 : std_logic;
signal n12587 : std_logic;
signal n1722 : std_logic;
signal n1789 : std_logic;
signal n12588 : std_logic;
signal n1721 : std_logic;
signal n1788 : std_logic;
signal n12589 : std_logic;
signal n1720 : std_logic;
signal n1787 : std_logic;
signal n12590 : std_logic;
signal n15622 : std_logic;
signal n12591 : std_logic;
signal n1818 : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal n12550 : std_logic;
signal n12551 : std_logic;
signal n12552 : std_logic;
signal n12553 : std_logic;
signal n12554 : std_logic;
signal n12555 : std_logic;
signal n12556 : std_logic;
signal n12557 : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal n12558 : std_logic;
signal n1591 : std_logic;
signal n12559 : std_logic;
signal n12560 : std_logic;
signal n12561 : std_logic;
signal n12562 : std_logic;
signal n13 : std_logic;
signal encoder0_position_20 : std_logic;
signal n27 : std_logic;
signal encoder0_position_6 : std_logic;
signal n313 : std_logic;
signal n11 : std_logic;
signal encoder0_position_22 : std_logic;
signal n11_adj_632 : std_logic;
signal n9 : std_logic;
signal n295 : std_logic;
signal encoder0_position_24 : std_logic;
signal n9_adj_630 : std_logic;
signal n933 : std_logic;
signal n1000 : std_logic;
signal \n1032_cascade_\ : std_logic;
signal \n11914_cascade_\ : std_logic;
signal \n13716_cascade_\ : std_logic;
signal \n1059_cascade_\ : std_logic;
signal \n1126_cascade_\ : std_logic;
signal n928 : std_logic;
signal n960 : std_logic;
signal n995 : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal n12500 : std_logic;
signal n12501 : std_logic;
signal n12502 : std_logic;
signal n12503 : std_logic;
signal n1029 : std_logic;
signal n1096 : std_logic;
signal n12504 : std_logic;
signal n1028 : std_logic;
signal n1095 : std_logic;
signal n12505 : std_logic;
signal n1027 : std_logic;
signal n1094 : std_logic;
signal n12506 : std_logic;
signal n12507 : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal n1026 : std_logic;
signal n1093 : std_logic;
signal n1030 : std_logic;
signal n1097 : std_logic;
signal pwm_counter_0 : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal pwm_counter_1 : std_logic;
signal \PWM.n13056\ : std_logic;
signal \PWM.n13057\ : std_logic;
signal \PWM.n13058\ : std_logic;
signal \PWM.n13059\ : std_logic;
signal \PWM.n13060\ : std_logic;
signal \PWM.n13061\ : std_logic;
signal \PWM.n13062\ : std_logic;
signal \PWM.n13063\ : std_logic;
signal \bfn_13_27_0_\ : std_logic;
signal \PWM.n13064\ : std_logic;
signal \PWM.n13065\ : std_logic;
signal \PWM.n13066\ : std_logic;
signal \PWM.n13067\ : std_logic;
signal \PWM.n13068\ : std_logic;
signal \PWM.n13069\ : std_logic;
signal \PWM.n13070\ : std_logic;
signal \PWM.n13071\ : std_logic;
signal \bfn_13_28_0_\ : std_logic;
signal \PWM.n13072\ : std_logic;
signal \PWM.n13073\ : std_logic;
signal \PWM.n13074\ : std_logic;
signal \PWM.n13075\ : std_logic;
signal \PWM.n13076\ : std_logic;
signal \PWM.n13077\ : std_logic;
signal \PWM.n13078\ : std_logic;
signal \PWM.n13079\ : std_logic;
signal \bfn_13_29_0_\ : std_logic;
signal \PWM.n13080\ : std_logic;
signal \PWM.n13081\ : std_logic;
signal \PWM.n13082\ : std_logic;
signal \PWM.n13083\ : std_logic;
signal \PWM.n13084\ : std_logic;
signal \PWM.n13085\ : std_logic;
signal \PWM.n13086\ : std_logic;
signal n6_adj_717 : std_logic;
signal pwm_setpoint_5 : std_logic;
signal pwm_setpoint_6 : std_logic;
signal pwm_setpoint_10 : std_logic;
signal pwm_setpoint_11 : std_logic;
signal pwm_setpoint_12 : std_logic;
signal pwm_setpoint_20 : std_logic;
signal n41 : std_logic;
signal \n41_cascade_\ : std_logic;
signal n15265 : std_logic;
signal n15112 : std_logic;
signal pwm_setpoint_23 : std_logic;
signal n15257 : std_logic;
signal n15108 : std_logic;
signal pwm_setpoint_21 : std_logic;
signal pwm_setpoint_19 : std_logic;
signal n39 : std_logic;
signal \n14910_cascade_\ : std_logic;
signal n1730 : std_logic;
signal \n14514_cascade_\ : std_logic;
signal \n1653_cascade_\ : std_logic;
signal n1598 : std_logic;
signal \n1630_adj_617_cascade_\ : std_logic;
signal n1729 : std_logic;
signal \n11902_cascade_\ : std_logic;
signal n13736 : std_logic;
signal n1599 : std_logic;
signal n1731 : std_logic;
signal n1733 : std_logic;
signal n303 : std_logic;
signal \n1731_cascade_\ : std_logic;
signal n11970 : std_logic;
signal n1732 : std_logic;
signal n1590 : std_logic;
signal n1589 : std_logic;
signal n1531 : std_logic;
signal \n1531_cascade_\ : std_logic;
signal n1592 : std_logic;
signal n1533 : std_logic;
signal n1600 : std_logic;
signal \n1533_cascade_\ : std_logic;
signal n15582 : std_logic;
signal \n14294_cascade_\ : std_logic;
signal n11974 : std_logic;
signal \n1527_cascade_\ : std_logic;
signal n14288 : std_logic;
signal n14 : std_logic;
signal \n1324_cascade_\ : std_logic;
signal encoder0_position_19 : std_logic;
signal n14_adj_635 : std_logic;
signal n1032 : std_logic;
signal n1099 : std_logic;
signal \n11908_cascade_\ : std_logic;
signal \n13708_cascade_\ : std_logic;
signal \n1356_cascade_\ : std_logic;
signal \n1433_cascade_\ : std_logic;
signal n1031 : std_logic;
signal n1098 : std_logic;
signal n296 : std_logic;
signal n1101 : std_logic;
signal \n1133_cascade_\ : std_logic;
signal n14428 : std_logic;
signal \n12000_cascade_\ : std_logic;
signal \n1158_cascade_\ : std_logic;
signal \n1232_cascade_\ : std_logic;
signal n12 : std_logic;
signal encoder0_position_31 : std_logic;
signal n1100 : std_logic;
signal n1033 : std_logic;
signal \n1132_cascade_\ : std_logic;
signal n1059 : std_logic;
signal n15499 : std_logic;
signal n14470 : std_logic;
signal encoder0_position_21 : std_logic;
signal n12_adj_633 : std_logic;
signal \n16_adj_701_cascade_\ : std_logic;
signal n24_adj_561 : std_logic;
signal n25 : std_logic;
signal \n13932_cascade_\ : std_logic;
signal \n14110_cascade_\ : std_logic;
signal n10_adj_567 : std_logic;
signal n15_adj_702 : std_logic;
signal n11853 : std_logic;
signal n23_adj_562 : std_logic;
signal pwm_setpoint_2 : std_logic;
signal pwm_setpoint_3 : std_logic;
signal pwm_counter_2 : std_logic;
signal pwm_counter_3 : std_logic;
signal pwm_counter_5 : std_logic;
signal pwm_counter_7 : std_logic;
signal pwm_counter_6 : std_logic;
signal pwm_counter_11 : std_logic;
signal pwm_counter_10 : std_logic;
signal pwm_counter_14 : std_logic;
signal pwm_counter_20 : std_logic;
signal pwm_counter_16 : std_logic;
signal pwm_counter_17 : std_logic;
signal pwm_counter_13 : std_logic;
signal pwm_counter_23 : std_logic;
signal pwm_counter_22 : std_logic;
signal pwm_counter_18 : std_logic;
signal pwm_counter_15 : std_logic;
signal pwm_counter_21 : std_logic;
signal pwm_counter_12 : std_logic;
signal \PWM.n26_cascade_\ : std_logic;
signal \PWM.n28\ : std_logic;
signal \PWM.n29_cascade_\ : std_logic;
signal \PWM.n27\ : std_logic;
signal \PWM.pwm_counter_31__N_407\ : std_logic;
signal pwm_counter_19 : std_logic;
signal \PWM.n13995\ : std_logic;
signal \PWM.n17\ : std_logic;
signal pwm_counter_24 : std_logic;
signal pwm_counter_29 : std_logic;
signal pwm_counter_27 : std_logic;
signal pwm_counter_26 : std_logic;
signal pwm_counter_30 : std_logic;
signal pwm_counter_25 : std_logic;
signal \n12_adj_566_cascade_\ : std_logic;
signal pwm_counter_28 : std_logic;
signal n5162 : std_logic;
signal \n5162_cascade_\ : std_logic;
signal pwm_counter_31 : std_logic;
signal n5164 : std_logic;
signal \pwm_setpoint_23_N_171_8\ : std_logic;
signal duty_8 : std_logic;
signal pwm_setpoint_4 : std_logic;
signal pwm_counter_4 : std_logic;
signal n15150 : std_logic;
signal n11_adj_660 : std_logic;
signal \n9_adj_658_cascade_\ : std_logic;
signal n13_adj_662 : std_logic;
signal n15_adj_663 : std_logic;
signal n15205 : std_logic;
signal \n15201_cascade_\ : std_logic;
signal n15261 : std_logic;
signal pwm_setpoint_8 : std_logic;
signal pwm_counter_8 : std_logic;
signal pwm_setpoint_9 : std_logic;
signal pwm_counter_9 : std_logic;
signal n21_adj_667 : std_logic;
signal n19_adj_666 : std_logic;
signal n17_adj_665 : std_logic;
signal n9_adj_658 : std_logic;
signal n43 : std_logic;
signal n23_adj_668 : std_logic;
signal \n15132_cascade_\ : std_logic;
signal n25_adj_670 : std_logic;
signal n15110 : std_logic;
signal \commutation_state_7__N_261\ : std_logic;
signal h3 : std_logic;
signal h1 : std_logic;
signal h2 : std_logic;
signal n302 : std_logic;
signal n1701 : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal n1700 : std_logic;
signal n12563 : std_logic;
signal n1632_adj_619 : std_logic;
signal n1699 : std_logic;
signal n12564 : std_logic;
signal n1631_adj_618 : std_logic;
signal n1698 : std_logic;
signal n12565 : std_logic;
signal n1630_adj_617 : std_logic;
signal n1697 : std_logic;
signal n12566 : std_logic;
signal n12567 : std_logic;
signal n12568 : std_logic;
signal n1694 : std_logic;
signal n12569 : std_logic;
signal n12570 : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal n12571 : std_logic;
signal n1624_adj_611 : std_logic;
signal n1691 : std_logic;
signal n12572 : std_logic;
signal n1623_adj_610 : std_logic;
signal n1690 : std_logic;
signal n12573 : std_logic;
signal n1622_adj_609 : std_logic;
signal n1689 : std_logic;
signal n12574 : std_logic;
signal n1621_adj_608 : std_logic;
signal n1688 : std_logic;
signal n12575 : std_logic;
signal n15603 : std_logic;
signal n1620_adj_607 : std_logic;
signal n12576 : std_logic;
signal n1719 : std_logic;
signal n1692 : std_logic;
signal n1523 : std_logic;
signal n1522 : std_logic;
signal \n1523_cascade_\ : std_logic;
signal n14296 : std_logic;
signal n1601 : std_logic;
signal \n1554_cascade_\ : std_logic;
signal n301 : std_logic;
signal n1633_adj_620 : std_logic;
signal n1532 : std_logic;
signal n11906 : std_logic;
signal \n14490_cascade_\ : std_logic;
signal n13727 : std_logic;
signal \n14496_cascade_\ : std_logic;
signal \n1455_cascade_\ : std_logic;
signal n1525 : std_logic;
signal n1524 : std_logic;
signal n299 : std_logic;
signal n1401 : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal n1400 : std_logic;
signal n12527 : std_logic;
signal n1399 : std_logic;
signal n12528 : std_logic;
signal n1331 : std_logic;
signal n1398 : std_logic;
signal n12529 : std_logic;
signal n1330 : std_logic;
signal n1397 : std_logic;
signal n12530 : std_logic;
signal n1396 : std_logic;
signal n12531 : std_logic;
signal n12532 : std_logic;
signal n1394 : std_logic;
signal n12533 : std_logic;
signal n12534 : std_logic;
signal n1393 : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal n12535 : std_logic;
signal n1324 : std_logic;
signal n1391 : std_logic;
signal n12536 : std_logic;
signal n15544 : std_logic;
signal n12537 : std_logic;
signal n1332 : std_logic;
signal n1329 : std_logic;
signal n1333 : std_logic;
signal n298 : std_logic;
signal n1301 : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal n1233 : std_logic;
signal n1300 : std_logic;
signal n12517 : std_logic;
signal n1232 : std_logic;
signal n1299 : std_logic;
signal n12518 : std_logic;
signal n1298 : std_logic;
signal n12519 : std_logic;
signal n1297 : std_logic;
signal n12520 : std_logic;
signal n12521 : std_logic;
signal n12522 : std_logic;
signal n12523 : std_logic;
signal n12524 : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal n1292 : std_logic;
signal n12525 : std_logic;
signal n12526 : std_logic;
signal n1323 : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal encoder0_position_target_0 : std_logic;
signal n12435 : std_logic;
signal encoder0_position_target_1 : std_logic;
signal n12436 : std_logic;
signal encoder0_position_target_2 : std_logic;
signal n12437 : std_logic;
signal encoder0_position_target_3 : std_logic;
signal n12438 : std_logic;
signal encoder0_position_target_4 : std_logic;
signal n12439 : std_logic;
signal encoder0_position_target_5 : std_logic;
signal n12440 : std_logic;
signal encoder0_position_target_6 : std_logic;
signal n12441 : std_logic;
signal n12442 : std_logic;
signal encoder0_position_target_7 : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal encoder0_position_target_8 : std_logic;
signal n12443 : std_logic;
signal encoder0_position_target_9 : std_logic;
signal n12444 : std_logic;
signal encoder0_position_target_10 : std_logic;
signal n12445 : std_logic;
signal encoder0_position_target_11 : std_logic;
signal n12446 : std_logic;
signal encoder0_position_target_12 : std_logic;
signal n12447 : std_logic;
signal encoder0_position_target_13 : std_logic;
signal n12448 : std_logic;
signal encoder0_position_target_14 : std_logic;
signal n12449 : std_logic;
signal n12450 : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal encoder0_position_target_16 : std_logic;
signal n12451 : std_logic;
signal encoder0_position_target_17 : std_logic;
signal n12452 : std_logic;
signal encoder0_position_target_18 : std_logic;
signal n12453 : std_logic;
signal n12454 : std_logic;
signal encoder0_position_target_20 : std_logic;
signal n12455 : std_logic;
signal n12456 : std_logic;
signal encoder0_position_target_22 : std_logic;
signal n12457 : std_logic;
signal n12458 : std_logic;
signal \bfn_15_28_0_\ : std_logic;
signal \n14_adj_718_cascade_\ : std_logic;
signal n10_adj_719 : std_logic;
signal \n5119_cascade_\ : std_logic;
signal n15088 : std_logic;
signal dti_counter_0 : std_logic;
signal \bfn_15_31_0_\ : std_logic;
signal n15095 : std_logic;
signal dti_counter_1 : std_logic;
signal n12961 : std_logic;
signal n15094 : std_logic;
signal dti_counter_2 : std_logic;
signal n12962 : std_logic;
signal n15093 : std_logic;
signal dti_counter_3 : std_logic;
signal n12963 : std_logic;
signal n15092 : std_logic;
signal dti_counter_4 : std_logic;
signal n12964 : std_logic;
signal n15091 : std_logic;
signal dti_counter_5 : std_logic;
signal n12965 : std_logic;
signal n12966 : std_logic;
signal n11514 : std_logic;
signal n15089 : std_logic;
signal n12967 : std_logic;
signal dti_counter_7 : std_logic;
signal \n4_adj_716_cascade_\ : std_logic;
signal dti_counter_6 : std_logic;
signal n15090 : std_logic;
signal commutation_state_prev_1 : std_logic;
signal commutation_state_prev_2 : std_logic;
signal n1693_adj_621 : std_logic;
signal n1695 : std_logic;
signal n1727 : std_logic;
signal \n1727_cascade_\ : std_logic;
signal n1726 : std_logic;
signal n1724 : std_logic;
signal n1725 : std_logic;
signal \n14166_cascade_\ : std_logic;
signal n1723 : std_logic;
signal n14172 : std_logic;
signal n1696 : std_logic;
signal n1653 : std_logic;
signal n1728 : std_logic;
signal n14508 : std_logic;
signal n1395 : std_logic;
signal \n1427_cascade_\ : std_logic;
signal n1526 : std_logic;
signal \n1526_cascade_\ : std_logic;
signal n1593 : std_logic;
signal n1625_adj_612 : std_logic;
signal n1528 : std_logic;
signal n1595 : std_logic;
signal n1627_adj_614 : std_logic;
signal n1527 : std_logic;
signal n1594 : std_logic;
signal n1626_adj_613 : std_logic;
signal n1529 : std_logic;
signal n1596 : std_logic;
signal n1628_adj_615 : std_logic;
signal n1597 : std_logic;
signal n1554 : std_logic;
signal n1530 : std_logic;
signal n1629_adj_616 : std_logic;
signal n300 : std_logic;
signal n1501 : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal n1433 : std_logic;
signal n1500 : std_logic;
signal n12538 : std_logic;
signal n1432 : std_logic;
signal n1499 : std_logic;
signal n12539 : std_logic;
signal n1431 : std_logic;
signal n1498 : std_logic;
signal n12540 : std_logic;
signal n1430 : std_logic;
signal n1497 : std_logic;
signal n12541 : std_logic;
signal n1429 : std_logic;
signal n1496 : std_logic;
signal n12542 : std_logic;
signal n1428 : std_logic;
signal n1495 : std_logic;
signal n12543 : std_logic;
signal n1427 : std_logic;
signal n1494 : std_logic;
signal n12544 : std_logic;
signal n12545 : std_logic;
signal n1426 : std_logic;
signal n1493 : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal n1425 : std_logic;
signal n1492 : std_logic;
signal n12546 : std_logic;
signal n1491 : std_logic;
signal n12547 : std_logic;
signal n1423 : std_logic;
signal n1490 : std_logic;
signal n12548 : std_logic;
signal n1422 : std_logic;
signal n12549 : std_logic;
signal n1521 : std_logic;
signal n1455 : std_logic;
signal n15562 : std_logic;
signal n1392 : std_logic;
signal n1356 : std_logic;
signal n1424 : std_logic;
signal n1294 : std_logic;
signal n1295 : std_logic;
signal n1227 : std_logic;
signal \n14482_cascade_\ : std_logic;
signal n1296 : std_logic;
signal \n1257_cascade_\ : std_logic;
signal n1328 : std_logic;
signal n1327 : std_logic;
signal \n1328_cascade_\ : std_logic;
signal n1326 : std_logic;
signal n14282 : std_logic;
signal n1226 : std_logic;
signal \n1226_cascade_\ : std_logic;
signal n1293 : std_logic;
signal n1325 : std_logic;
signal n1229 : std_logic;
signal n11910 : std_logic;
signal \n1229_cascade_\ : std_logic;
signal n1231 : std_logic;
signal n13711 : std_logic;
signal n1257 : std_logic;
signal n15528 : std_logic;
signal n1228 : std_logic;
signal n1230 : std_logic;
signal n297 : std_logic;
signal n1201 : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal n1133 : std_logic;
signal n1200 : std_logic;
signal n12508 : std_logic;
signal n1132 : std_logic;
signal n1199 : std_logic;
signal n12509 : std_logic;
signal n1131 : std_logic;
signal n1198 : std_logic;
signal n12510 : std_logic;
signal n1130 : std_logic;
signal n1197 : std_logic;
signal n12511 : std_logic;
signal n1129 : std_logic;
signal n1196 : std_logic;
signal n12512 : std_logic;
signal n1128 : std_logic;
signal n1195 : std_logic;
signal n12513 : std_logic;
signal n1127 : std_logic;
signal n1194 : std_logic;
signal n12514 : std_logic;
signal n12515 : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n15513 : std_logic;
signal n1125 : std_logic;
signal n12516 : std_logic;
signal n1224 : std_logic;
signal n1126 : std_logic;
signal n1193 : std_logic;
signal n1158 : std_logic;
signal n1225 : std_logic;
signal n23_adj_700 : std_logic;
signal n25_adj_698 : std_logic;
signal \direction_N_342_cascade_\ : std_logic;
signal n1693 : std_logic;
signal \direction_N_340\ : std_logic;
signal \direction_N_342\ : std_logic;
signal \n13661_cascade_\ : std_logic;
signal direction_c : std_logic;
signal \n22_adj_705_cascade_\ : std_logic;
signal \n6_adj_582_cascade_\ : std_logic;
signal n14108 : std_logic;
signal encoder0_position_target_15 : std_logic;
signal encoder0_position_target_21 : std_logic;
signal encoder0_position_target_19 : std_logic;
signal encoder0_position_target_23 : std_logic;
signal n24_adj_699 : std_logic;
signal n16_adj_707 : std_logic;
signal commutation_state_prev_0 : std_logic;
signal \dti_N_333_cascade_\ : std_logic;
signal n4_adj_716 : std_logic;
signal n5169 : std_logic;
signal n1377 : std_logic;
signal n5119 : std_logic;
signal \n5183_cascade_\ : std_logic;
signal dti : std_logic;
signal \n20_adj_706_cascade_\ : std_logic;
signal n24_adj_704 : std_logic;
signal n13187 : std_logic;
signal sweep_counter_0 : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal sweep_counter_1 : std_logic;
signal n12999 : std_logic;
signal sweep_counter_2 : std_logic;
signal n13000 : std_logic;
signal sweep_counter_3 : std_logic;
signal n13001 : std_logic;
signal sweep_counter_4 : std_logic;
signal n13002 : std_logic;
signal sweep_counter_5 : std_logic;
signal n13003 : std_logic;
signal sweep_counter_6 : std_logic;
signal n13004 : std_logic;
signal sweep_counter_7 : std_logic;
signal n13005 : std_logic;
signal n13006 : std_logic;
signal sweep_counter_8 : std_logic;
signal \bfn_17_27_0_\ : std_logic;
signal sweep_counter_9 : std_logic;
signal n13007 : std_logic;
signal sweep_counter_10 : std_logic;
signal n13008 : std_logic;
signal sweep_counter_11 : std_logic;
signal n13009 : std_logic;
signal sweep_counter_12 : std_logic;
signal n13010 : std_logic;
signal sweep_counter_13 : std_logic;
signal n13011 : std_logic;
signal sweep_counter_14 : std_logic;
signal n13012 : std_logic;
signal sweep_counter_15 : std_logic;
signal n13013 : std_logic;
signal n13014 : std_logic;
signal sweep_counter_16 : std_logic;
signal \bfn_17_28_0_\ : std_logic;
signal n13015 : std_logic;
signal sweep_counter_17 : std_logic;
signal n5197 : std_logic;
signal duty_23 : std_logic;
signal \INLB_c_0\ : std_logic;
signal \INLA_c_0\ : std_logic;
signal commutation_state_0 : std_logic;
signal commutation_state_1 : std_logic;
signal commutation_state_2 : std_logic;
signal dir : std_logic;
signal \INLC_c_0\ : std_logic;
signal \CLK_N\ : std_logic;
signal n5183 : std_logic;
signal n5235 : std_logic;
signal \GHB\ : std_logic;
signal \INHB_c_0\ : std_logic;
signal \GHC\ : std_logic;
signal \INHC_c_0\ : std_logic;
signal pwm_out : std_logic;
signal \GHA\ : std_logic;
signal \INHA_c_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \ENCODER0_A_wire\ : std_logic;
signal \ENCODER0_B_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \HALL1_wire\ : std_logic;
signal \HALL2_wire\ : std_logic;
signal \HALL3_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    \ENCODER0_A_wire\ <= ENCODER0_A;
    \ENCODER0_B_wire\ <= ENCODER0_B;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \HALL1_wire\ <= HALL1;
    \HALL2_wire\ <= HALL2;
    \HALL3_wire\ <= HALL3;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56344\,
            DIN => \N__56343\,
            DOUT => \N__56342\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56344\,
            PADOUT => \N__56343\,
            PADIN => \N__56342\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56335\,
            DIN => \N__56334\,
            DOUT => \N__56333\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56335\,
            PADOUT => \N__56334\,
            PADIN => \N__56333\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56326\,
            DIN => \N__56325\,
            DOUT => \N__56324\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56326\,
            PADOUT => \N__56325\,
            PADIN => \N__56324\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ENCODER0_A_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56317\,
            DIN => \N__56316\,
            DOUT => \N__56315\,
            PACKAGEPIN => \ENCODER0_A_wire\
        );

    \ENCODER0_A_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56317\,
            PADOUT => \N__56316\,
            PADIN => \N__56315\,
            CLOCKENABLE => 'H',
            DIN0 => \ENCODER0_A_N\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ENCODER0_B_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56308\,
            DIN => \N__56307\,
            DOUT => \N__56306\,
            PACKAGEPIN => \ENCODER0_B_wire\
        );

    \ENCODER0_B_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56308\,
            PADOUT => \N__56307\,
            PADIN => \N__56306\,
            CLOCKENABLE => 'H',
            DIN0 => \ENCODER0_B_N\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56299\,
            DIN => \N__56298\,
            DOUT => \N__56297\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56299\,
            PADOUT => \N__56298\,
            PADIN => \N__56297\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55479\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56290\,
            DIN => \N__56289\,
            DOUT => \N__56288\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56290\,
            PADOUT => \N__56289\,
            PADIN => \N__56288\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55548\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56281\,
            DIN => \N__56280\,
            DOUT => \N__56279\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56281\,
            PADOUT => \N__56280\,
            PADIN => \N__56279\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55527\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56272\,
            DIN => \N__56271\,
            DOUT => \N__56270\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56272\,
            PADOUT => \N__56271\,
            PADIN => \N__56270\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__56163\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56263\,
            DIN => \N__56262\,
            DOUT => \N__56261\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56263\,
            PADOUT => \N__56262\,
            PADIN => \N__56261\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55191\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56254\,
            DIN => \N__56253\,
            DOUT => \N__56252\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56254\,
            PADOUT => \N__56253\,
            PADIN => \N__56252\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55854\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56245\,
            DIN => \N__56244\,
            DOUT => \N__56243\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56245\,
            PADOUT => \N__56244\,
            PADIN => \N__56243\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__39489\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56236\,
            DIN => \N__56235\,
            DOUT => \N__56234\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56236\,
            PADOUT => \N__56235\,
            PADIN => \N__56234\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56227\,
            DIN => \N__56226\,
            DOUT => \N__56225\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56227\,
            PADOUT => \N__56226\,
            PADIN => \N__56225\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56218\,
            DIN => \N__56217\,
            DOUT => \N__56216\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56218\,
            PADOUT => \N__56217\,
            PADIN => \N__56216\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall1_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56209\,
            DIN => \N__56208\,
            DOUT => \N__56207\,
            PACKAGEPIN => \HALL1_wire\
        );

    \hall1_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56209\,
            PADOUT => \N__56208\,
            PADIN => \N__56207\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_2\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__55776\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall2_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56200\,
            DIN => \N__56199\,
            DOUT => \N__56198\,
            PACKAGEPIN => \HALL2_wire\
        );

    \hall2_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56200\,
            PADOUT => \N__56199\,
            PADIN => \N__56198\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_1\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__55774\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall3_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56191\,
            DIN => \N__56190\,
            DOUT => \N__56189\,
            PACKAGEPIN => \HALL3_wire\
        );

    \hall3_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56191\,
            PADOUT => \N__56190\,
            PADIN => \N__56189\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_0\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__55774\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56182\,
            DIN => \N__56181\,
            DOUT => \N__56180\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56182\,
            PADOUT => \N__56181\,
            PADIN => \N__56180\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__13316\ : IoInMux
    port map (
            O => \N__56163\,
            I => \N__56160\
        );

    \I__13315\ : LocalMux
    port map (
            O => \N__56160\,
            I => \N__56157\
        );

    \I__13314\ : IoSpan4Mux
    port map (
            O => \N__56157\,
            I => \N__56154\
        );

    \I__13313\ : Span4Mux_s0_v
    port map (
            O => \N__56154\,
            I => \N__56151\
        );

    \I__13312\ : Odrv4
    port map (
            O => \N__56151\,
            I => \INLA_c_0\
        );

    \I__13311\ : InMux
    port map (
            O => \N__56148\,
            I => \N__56140\
        );

    \I__13310\ : InMux
    port map (
            O => \N__56147\,
            I => \N__56137\
        );

    \I__13309\ : InMux
    port map (
            O => \N__56146\,
            I => \N__56132\
        );

    \I__13308\ : InMux
    port map (
            O => \N__56145\,
            I => \N__56132\
        );

    \I__13307\ : InMux
    port map (
            O => \N__56144\,
            I => \N__56127\
        );

    \I__13306\ : InMux
    port map (
            O => \N__56143\,
            I => \N__56127\
        );

    \I__13305\ : LocalMux
    port map (
            O => \N__56140\,
            I => \N__56119\
        );

    \I__13304\ : LocalMux
    port map (
            O => \N__56137\,
            I => \N__56119\
        );

    \I__13303\ : LocalMux
    port map (
            O => \N__56132\,
            I => \N__56113\
        );

    \I__13302\ : LocalMux
    port map (
            O => \N__56127\,
            I => \N__56113\
        );

    \I__13301\ : InMux
    port map (
            O => \N__56126\,
            I => \N__56107\
        );

    \I__13300\ : InMux
    port map (
            O => \N__56125\,
            I => \N__56102\
        );

    \I__13299\ : InMux
    port map (
            O => \N__56124\,
            I => \N__56102\
        );

    \I__13298\ : Span4Mux_v
    port map (
            O => \N__56119\,
            I => \N__56096\
        );

    \I__13297\ : InMux
    port map (
            O => \N__56118\,
            I => \N__56093\
        );

    \I__13296\ : Span4Mux_s2_v
    port map (
            O => \N__56113\,
            I => \N__56090\
        );

    \I__13295\ : InMux
    port map (
            O => \N__56112\,
            I => \N__56083\
        );

    \I__13294\ : InMux
    port map (
            O => \N__56111\,
            I => \N__56083\
        );

    \I__13293\ : InMux
    port map (
            O => \N__56110\,
            I => \N__56083\
        );

    \I__13292\ : LocalMux
    port map (
            O => \N__56107\,
            I => \N__56080\
        );

    \I__13291\ : LocalMux
    port map (
            O => \N__56102\,
            I => \N__56077\
        );

    \I__13290\ : InMux
    port map (
            O => \N__56101\,
            I => \N__56074\
        );

    \I__13289\ : InMux
    port map (
            O => \N__56100\,
            I => \N__56069\
        );

    \I__13288\ : InMux
    port map (
            O => \N__56099\,
            I => \N__56069\
        );

    \I__13287\ : Span4Mux_h
    port map (
            O => \N__56096\,
            I => \N__56064\
        );

    \I__13286\ : LocalMux
    port map (
            O => \N__56093\,
            I => \N__56064\
        );

    \I__13285\ : Span4Mux_h
    port map (
            O => \N__56090\,
            I => \N__56055\
        );

    \I__13284\ : LocalMux
    port map (
            O => \N__56083\,
            I => \N__56055\
        );

    \I__13283\ : Span4Mux_h
    port map (
            O => \N__56080\,
            I => \N__56055\
        );

    \I__13282\ : Span4Mux_s2_v
    port map (
            O => \N__56077\,
            I => \N__56055\
        );

    \I__13281\ : LocalMux
    port map (
            O => \N__56074\,
            I => commutation_state_0
        );

    \I__13280\ : LocalMux
    port map (
            O => \N__56069\,
            I => commutation_state_0
        );

    \I__13279\ : Odrv4
    port map (
            O => \N__56064\,
            I => commutation_state_0
        );

    \I__13278\ : Odrv4
    port map (
            O => \N__56055\,
            I => commutation_state_0
        );

    \I__13277\ : CascadeMux
    port map (
            O => \N__56046\,
            I => \N__56040\
        );

    \I__13276\ : CascadeMux
    port map (
            O => \N__56045\,
            I => \N__56037\
        );

    \I__13275\ : InMux
    port map (
            O => \N__56044\,
            I => \N__56031\
        );

    \I__13274\ : InMux
    port map (
            O => \N__56043\,
            I => \N__56031\
        );

    \I__13273\ : InMux
    port map (
            O => \N__56040\,
            I => \N__56024\
        );

    \I__13272\ : InMux
    port map (
            O => \N__56037\,
            I => \N__56024\
        );

    \I__13271\ : InMux
    port map (
            O => \N__56036\,
            I => \N__56021\
        );

    \I__13270\ : LocalMux
    port map (
            O => \N__56031\,
            I => \N__56018\
        );

    \I__13269\ : InMux
    port map (
            O => \N__56030\,
            I => \N__56014\
        );

    \I__13268\ : CascadeMux
    port map (
            O => \N__56029\,
            I => \N__56010\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__56024\,
            I => \N__56003\
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__56021\,
            I => \N__56003\
        );

    \I__13265\ : Span4Mux_s1_v
    port map (
            O => \N__56018\,
            I => \N__56003\
        );

    \I__13264\ : CascadeMux
    port map (
            O => \N__56017\,
            I => \N__55999\
        );

    \I__13263\ : LocalMux
    port map (
            O => \N__56014\,
            I => \N__55996\
        );

    \I__13262\ : InMux
    port map (
            O => \N__56013\,
            I => \N__55993\
        );

    \I__13261\ : InMux
    port map (
            O => \N__56010\,
            I => \N__55990\
        );

    \I__13260\ : Span4Mux_h
    port map (
            O => \N__56003\,
            I => \N__55987\
        );

    \I__13259\ : InMux
    port map (
            O => \N__56002\,
            I => \N__55982\
        );

    \I__13258\ : InMux
    port map (
            O => \N__55999\,
            I => \N__55982\
        );

    \I__13257\ : Span4Mux_s1_v
    port map (
            O => \N__55996\,
            I => \N__55977\
        );

    \I__13256\ : LocalMux
    port map (
            O => \N__55993\,
            I => \N__55977\
        );

    \I__13255\ : LocalMux
    port map (
            O => \N__55990\,
            I => commutation_state_1
        );

    \I__13254\ : Odrv4
    port map (
            O => \N__55987\,
            I => commutation_state_1
        );

    \I__13253\ : LocalMux
    port map (
            O => \N__55982\,
            I => commutation_state_1
        );

    \I__13252\ : Odrv4
    port map (
            O => \N__55977\,
            I => commutation_state_1
        );

    \I__13251\ : CascadeMux
    port map (
            O => \N__55968\,
            I => \N__55965\
        );

    \I__13250\ : InMux
    port map (
            O => \N__55965\,
            I => \N__55957\
        );

    \I__13249\ : InMux
    port map (
            O => \N__55964\,
            I => \N__55952\
        );

    \I__13248\ : InMux
    port map (
            O => \N__55963\,
            I => \N__55952\
        );

    \I__13247\ : CascadeMux
    port map (
            O => \N__55962\,
            I => \N__55947\
        );

    \I__13246\ : CascadeMux
    port map (
            O => \N__55961\,
            I => \N__55944\
        );

    \I__13245\ : CascadeMux
    port map (
            O => \N__55960\,
            I => \N__55941\
        );

    \I__13244\ : LocalMux
    port map (
            O => \N__55957\,
            I => \N__55936\
        );

    \I__13243\ : LocalMux
    port map (
            O => \N__55952\,
            I => \N__55936\
        );

    \I__13242\ : InMux
    port map (
            O => \N__55951\,
            I => \N__55933\
        );

    \I__13241\ : CascadeMux
    port map (
            O => \N__55950\,
            I => \N__55930\
        );

    \I__13240\ : InMux
    port map (
            O => \N__55947\,
            I => \N__55927\
        );

    \I__13239\ : InMux
    port map (
            O => \N__55944\,
            I => \N__55922\
        );

    \I__13238\ : InMux
    port map (
            O => \N__55941\,
            I => \N__55922\
        );

    \I__13237\ : Span4Mux_h
    port map (
            O => \N__55936\,
            I => \N__55915\
        );

    \I__13236\ : LocalMux
    port map (
            O => \N__55933\,
            I => \N__55915\
        );

    \I__13235\ : InMux
    port map (
            O => \N__55930\,
            I => \N__55912\
        );

    \I__13234\ : LocalMux
    port map (
            O => \N__55927\,
            I => \N__55907\
        );

    \I__13233\ : LocalMux
    port map (
            O => \N__55922\,
            I => \N__55907\
        );

    \I__13232\ : InMux
    port map (
            O => \N__55921\,
            I => \N__55902\
        );

    \I__13231\ : InMux
    port map (
            O => \N__55920\,
            I => \N__55902\
        );

    \I__13230\ : Span4Mux_h
    port map (
            O => \N__55915\,
            I => \N__55899\
        );

    \I__13229\ : LocalMux
    port map (
            O => \N__55912\,
            I => commutation_state_2
        );

    \I__13228\ : Odrv12
    port map (
            O => \N__55907\,
            I => commutation_state_2
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__55902\,
            I => commutation_state_2
        );

    \I__13226\ : Odrv4
    port map (
            O => \N__55899\,
            I => commutation_state_2
        );

    \I__13225\ : InMux
    port map (
            O => \N__55890\,
            I => \N__55884\
        );

    \I__13224\ : InMux
    port map (
            O => \N__55889\,
            I => \N__55884\
        );

    \I__13223\ : LocalMux
    port map (
            O => \N__55884\,
            I => \N__55878\
        );

    \I__13222\ : InMux
    port map (
            O => \N__55883\,
            I => \N__55873\
        );

    \I__13221\ : InMux
    port map (
            O => \N__55882\,
            I => \N__55873\
        );

    \I__13220\ : InMux
    port map (
            O => \N__55881\,
            I => \N__55869\
        );

    \I__13219\ : Span4Mux_v
    port map (
            O => \N__55878\,
            I => \N__55864\
        );

    \I__13218\ : LocalMux
    port map (
            O => \N__55873\,
            I => \N__55864\
        );

    \I__13217\ : InMux
    port map (
            O => \N__55872\,
            I => \N__55861\
        );

    \I__13216\ : LocalMux
    port map (
            O => \N__55869\,
            I => dir
        );

    \I__13215\ : Odrv4
    port map (
            O => \N__55864\,
            I => dir
        );

    \I__13214\ : LocalMux
    port map (
            O => \N__55861\,
            I => dir
        );

    \I__13213\ : IoInMux
    port map (
            O => \N__55854\,
            I => \N__55851\
        );

    \I__13212\ : LocalMux
    port map (
            O => \N__55851\,
            I => \N__55848\
        );

    \I__13211\ : Span4Mux_s0_v
    port map (
            O => \N__55848\,
            I => \N__55845\
        );

    \I__13210\ : Span4Mux_h
    port map (
            O => \N__55845\,
            I => \N__55842\
        );

    \I__13209\ : Span4Mux_h
    port map (
            O => \N__55842\,
            I => \N__55839\
        );

    \I__13208\ : Odrv4
    port map (
            O => \N__55839\,
            I => \INLC_c_0\
        );

    \I__13207\ : ClkMux
    port map (
            O => \N__55836\,
            I => \N__55644\
        );

    \I__13206\ : ClkMux
    port map (
            O => \N__55835\,
            I => \N__55644\
        );

    \I__13205\ : ClkMux
    port map (
            O => \N__55834\,
            I => \N__55644\
        );

    \I__13204\ : ClkMux
    port map (
            O => \N__55833\,
            I => \N__55644\
        );

    \I__13203\ : ClkMux
    port map (
            O => \N__55832\,
            I => \N__55644\
        );

    \I__13202\ : ClkMux
    port map (
            O => \N__55831\,
            I => \N__55644\
        );

    \I__13201\ : ClkMux
    port map (
            O => \N__55830\,
            I => \N__55644\
        );

    \I__13200\ : ClkMux
    port map (
            O => \N__55829\,
            I => \N__55644\
        );

    \I__13199\ : ClkMux
    port map (
            O => \N__55828\,
            I => \N__55644\
        );

    \I__13198\ : ClkMux
    port map (
            O => \N__55827\,
            I => \N__55644\
        );

    \I__13197\ : ClkMux
    port map (
            O => \N__55826\,
            I => \N__55644\
        );

    \I__13196\ : ClkMux
    port map (
            O => \N__55825\,
            I => \N__55644\
        );

    \I__13195\ : ClkMux
    port map (
            O => \N__55824\,
            I => \N__55644\
        );

    \I__13194\ : ClkMux
    port map (
            O => \N__55823\,
            I => \N__55644\
        );

    \I__13193\ : ClkMux
    port map (
            O => \N__55822\,
            I => \N__55644\
        );

    \I__13192\ : ClkMux
    port map (
            O => \N__55821\,
            I => \N__55644\
        );

    \I__13191\ : ClkMux
    port map (
            O => \N__55820\,
            I => \N__55644\
        );

    \I__13190\ : ClkMux
    port map (
            O => \N__55819\,
            I => \N__55644\
        );

    \I__13189\ : ClkMux
    port map (
            O => \N__55818\,
            I => \N__55644\
        );

    \I__13188\ : ClkMux
    port map (
            O => \N__55817\,
            I => \N__55644\
        );

    \I__13187\ : ClkMux
    port map (
            O => \N__55816\,
            I => \N__55644\
        );

    \I__13186\ : ClkMux
    port map (
            O => \N__55815\,
            I => \N__55644\
        );

    \I__13185\ : ClkMux
    port map (
            O => \N__55814\,
            I => \N__55644\
        );

    \I__13184\ : ClkMux
    port map (
            O => \N__55813\,
            I => \N__55644\
        );

    \I__13183\ : ClkMux
    port map (
            O => \N__55812\,
            I => \N__55644\
        );

    \I__13182\ : ClkMux
    port map (
            O => \N__55811\,
            I => \N__55644\
        );

    \I__13181\ : ClkMux
    port map (
            O => \N__55810\,
            I => \N__55644\
        );

    \I__13180\ : ClkMux
    port map (
            O => \N__55809\,
            I => \N__55644\
        );

    \I__13179\ : ClkMux
    port map (
            O => \N__55808\,
            I => \N__55644\
        );

    \I__13178\ : ClkMux
    port map (
            O => \N__55807\,
            I => \N__55644\
        );

    \I__13177\ : ClkMux
    port map (
            O => \N__55806\,
            I => \N__55644\
        );

    \I__13176\ : ClkMux
    port map (
            O => \N__55805\,
            I => \N__55644\
        );

    \I__13175\ : ClkMux
    port map (
            O => \N__55804\,
            I => \N__55644\
        );

    \I__13174\ : ClkMux
    port map (
            O => \N__55803\,
            I => \N__55644\
        );

    \I__13173\ : ClkMux
    port map (
            O => \N__55802\,
            I => \N__55644\
        );

    \I__13172\ : ClkMux
    port map (
            O => \N__55801\,
            I => \N__55644\
        );

    \I__13171\ : ClkMux
    port map (
            O => \N__55800\,
            I => \N__55644\
        );

    \I__13170\ : ClkMux
    port map (
            O => \N__55799\,
            I => \N__55644\
        );

    \I__13169\ : ClkMux
    port map (
            O => \N__55798\,
            I => \N__55644\
        );

    \I__13168\ : ClkMux
    port map (
            O => \N__55797\,
            I => \N__55644\
        );

    \I__13167\ : ClkMux
    port map (
            O => \N__55796\,
            I => \N__55644\
        );

    \I__13166\ : ClkMux
    port map (
            O => \N__55795\,
            I => \N__55644\
        );

    \I__13165\ : ClkMux
    port map (
            O => \N__55794\,
            I => \N__55644\
        );

    \I__13164\ : ClkMux
    port map (
            O => \N__55793\,
            I => \N__55644\
        );

    \I__13163\ : ClkMux
    port map (
            O => \N__55792\,
            I => \N__55644\
        );

    \I__13162\ : ClkMux
    port map (
            O => \N__55791\,
            I => \N__55644\
        );

    \I__13161\ : ClkMux
    port map (
            O => \N__55790\,
            I => \N__55644\
        );

    \I__13160\ : ClkMux
    port map (
            O => \N__55789\,
            I => \N__55644\
        );

    \I__13159\ : ClkMux
    port map (
            O => \N__55788\,
            I => \N__55644\
        );

    \I__13158\ : ClkMux
    port map (
            O => \N__55787\,
            I => \N__55644\
        );

    \I__13157\ : ClkMux
    port map (
            O => \N__55786\,
            I => \N__55644\
        );

    \I__13156\ : ClkMux
    port map (
            O => \N__55785\,
            I => \N__55644\
        );

    \I__13155\ : ClkMux
    port map (
            O => \N__55784\,
            I => \N__55644\
        );

    \I__13154\ : ClkMux
    port map (
            O => \N__55783\,
            I => \N__55644\
        );

    \I__13153\ : ClkMux
    port map (
            O => \N__55782\,
            I => \N__55644\
        );

    \I__13152\ : ClkMux
    port map (
            O => \N__55781\,
            I => \N__55644\
        );

    \I__13151\ : ClkMux
    port map (
            O => \N__55780\,
            I => \N__55644\
        );

    \I__13150\ : ClkMux
    port map (
            O => \N__55779\,
            I => \N__55644\
        );

    \I__13149\ : ClkMux
    port map (
            O => \N__55778\,
            I => \N__55644\
        );

    \I__13148\ : ClkMux
    port map (
            O => \N__55777\,
            I => \N__55644\
        );

    \I__13147\ : ClkMux
    port map (
            O => \N__55776\,
            I => \N__55644\
        );

    \I__13146\ : ClkMux
    port map (
            O => \N__55775\,
            I => \N__55644\
        );

    \I__13145\ : ClkMux
    port map (
            O => \N__55774\,
            I => \N__55644\
        );

    \I__13144\ : ClkMux
    port map (
            O => \N__55773\,
            I => \N__55644\
        );

    \I__13143\ : GlobalMux
    port map (
            O => \N__55644\,
            I => \N__55641\
        );

    \I__13142\ : gio2CtrlBuf
    port map (
            O => \N__55641\,
            I => \CLK_N\
        );

    \I__13141\ : CEMux
    port map (
            O => \N__55638\,
            I => \N__55634\
        );

    \I__13140\ : CEMux
    port map (
            O => \N__55637\,
            I => \N__55630\
        );

    \I__13139\ : LocalMux
    port map (
            O => \N__55634\,
            I => \N__55626\
        );

    \I__13138\ : CEMux
    port map (
            O => \N__55633\,
            I => \N__55623\
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__55630\,
            I => \N__55620\
        );

    \I__13136\ : CEMux
    port map (
            O => \N__55629\,
            I => \N__55617\
        );

    \I__13135\ : Span4Mux_s1_v
    port map (
            O => \N__55626\,
            I => \N__55612\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__55623\,
            I => \N__55612\
        );

    \I__13133\ : Span4Mux_s1_v
    port map (
            O => \N__55620\,
            I => \N__55609\
        );

    \I__13132\ : LocalMux
    port map (
            O => \N__55617\,
            I => \N__55606\
        );

    \I__13131\ : Span4Mux_v
    port map (
            O => \N__55612\,
            I => \N__55603\
        );

    \I__13130\ : Odrv4
    port map (
            O => \N__55609\,
            I => n5183
        );

    \I__13129\ : Odrv12
    port map (
            O => \N__55606\,
            I => n5183
        );

    \I__13128\ : Odrv4
    port map (
            O => \N__55603\,
            I => n5183
        );

    \I__13127\ : SRMux
    port map (
            O => \N__55596\,
            I => \N__55593\
        );

    \I__13126\ : LocalMux
    port map (
            O => \N__55593\,
            I => \N__55587\
        );

    \I__13125\ : SRMux
    port map (
            O => \N__55592\,
            I => \N__55584\
        );

    \I__13124\ : SRMux
    port map (
            O => \N__55591\,
            I => \N__55581\
        );

    \I__13123\ : SRMux
    port map (
            O => \N__55590\,
            I => \N__55578\
        );

    \I__13122\ : Span4Mux_h
    port map (
            O => \N__55587\,
            I => \N__55573\
        );

    \I__13121\ : LocalMux
    port map (
            O => \N__55584\,
            I => \N__55573\
        );

    \I__13120\ : LocalMux
    port map (
            O => \N__55581\,
            I => \N__55568\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__55578\,
            I => \N__55568\
        );

    \I__13118\ : Span4Mux_h
    port map (
            O => \N__55573\,
            I => \N__55565\
        );

    \I__13117\ : Span4Mux_s1_v
    port map (
            O => \N__55568\,
            I => \N__55560\
        );

    \I__13116\ : Span4Mux_s1_v
    port map (
            O => \N__55565\,
            I => \N__55560\
        );

    \I__13115\ : Odrv4
    port map (
            O => \N__55560\,
            I => n5235
        );

    \I__13114\ : InMux
    port map (
            O => \N__55557\,
            I => \N__55554\
        );

    \I__13113\ : LocalMux
    port map (
            O => \N__55554\,
            I => \N__55551\
        );

    \I__13112\ : Odrv12
    port map (
            O => \N__55551\,
            I => \GHB\
        );

    \I__13111\ : IoInMux
    port map (
            O => \N__55548\,
            I => \N__55545\
        );

    \I__13110\ : LocalMux
    port map (
            O => \N__55545\,
            I => \N__55542\
        );

    \I__13109\ : Span4Mux_s1_v
    port map (
            O => \N__55542\,
            I => \N__55539\
        );

    \I__13108\ : Span4Mux_h
    port map (
            O => \N__55539\,
            I => \N__55536\
        );

    \I__13107\ : Odrv4
    port map (
            O => \N__55536\,
            I => \INHB_c_0\
        );

    \I__13106\ : InMux
    port map (
            O => \N__55533\,
            I => \N__55530\
        );

    \I__13105\ : LocalMux
    port map (
            O => \N__55530\,
            I => \GHC\
        );

    \I__13104\ : IoInMux
    port map (
            O => \N__55527\,
            I => \N__55524\
        );

    \I__13103\ : LocalMux
    port map (
            O => \N__55524\,
            I => \N__55521\
        );

    \I__13102\ : Span4Mux_s1_v
    port map (
            O => \N__55521\,
            I => \N__55518\
        );

    \I__13101\ : Span4Mux_h
    port map (
            O => \N__55518\,
            I => \N__55515\
        );

    \I__13100\ : Odrv4
    port map (
            O => \N__55515\,
            I => \INHC_c_0\
        );

    \I__13099\ : InMux
    port map (
            O => \N__55512\,
            I => \N__55509\
        );

    \I__13098\ : LocalMux
    port map (
            O => \N__55509\,
            I => \N__55506\
        );

    \I__13097\ : Span4Mux_s1_v
    port map (
            O => \N__55506\,
            I => \N__55501\
        );

    \I__13096\ : InMux
    port map (
            O => \N__55505\,
            I => \N__55496\
        );

    \I__13095\ : InMux
    port map (
            O => \N__55504\,
            I => \N__55496\
        );

    \I__13094\ : Sp12to4
    port map (
            O => \N__55501\,
            I => \N__55491\
        );

    \I__13093\ : LocalMux
    port map (
            O => \N__55496\,
            I => \N__55491\
        );

    \I__13092\ : Odrv12
    port map (
            O => \N__55491\,
            I => pwm_out
        );

    \I__13091\ : InMux
    port map (
            O => \N__55488\,
            I => \N__55485\
        );

    \I__13090\ : LocalMux
    port map (
            O => \N__55485\,
            I => \N__55482\
        );

    \I__13089\ : Odrv12
    port map (
            O => \N__55482\,
            I => \GHA\
        );

    \I__13088\ : IoInMux
    port map (
            O => \N__55479\,
            I => \N__55476\
        );

    \I__13087\ : LocalMux
    port map (
            O => \N__55476\,
            I => \N__55473\
        );

    \I__13086\ : Span4Mux_s0_v
    port map (
            O => \N__55473\,
            I => \N__55470\
        );

    \I__13085\ : Odrv4
    port map (
            O => \N__55470\,
            I => \INHA_c_0\
        );

    \I__13084\ : InMux
    port map (
            O => \N__55467\,
            I => \N__55463\
        );

    \I__13083\ : InMux
    port map (
            O => \N__55466\,
            I => \N__55460\
        );

    \I__13082\ : LocalMux
    port map (
            O => \N__55463\,
            I => sweep_counter_14
        );

    \I__13081\ : LocalMux
    port map (
            O => \N__55460\,
            I => sweep_counter_14
        );

    \I__13080\ : InMux
    port map (
            O => \N__55455\,
            I => n13012
        );

    \I__13079\ : InMux
    port map (
            O => \N__55452\,
            I => \N__55448\
        );

    \I__13078\ : InMux
    port map (
            O => \N__55451\,
            I => \N__55445\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__55448\,
            I => sweep_counter_15
        );

    \I__13076\ : LocalMux
    port map (
            O => \N__55445\,
            I => sweep_counter_15
        );

    \I__13075\ : InMux
    port map (
            O => \N__55440\,
            I => n13013
        );

    \I__13074\ : InMux
    port map (
            O => \N__55437\,
            I => \N__55433\
        );

    \I__13073\ : InMux
    port map (
            O => \N__55436\,
            I => \N__55430\
        );

    \I__13072\ : LocalMux
    port map (
            O => \N__55433\,
            I => \N__55427\
        );

    \I__13071\ : LocalMux
    port map (
            O => \N__55430\,
            I => sweep_counter_16
        );

    \I__13070\ : Odrv4
    port map (
            O => \N__55427\,
            I => sweep_counter_16
        );

    \I__13069\ : InMux
    port map (
            O => \N__55422\,
            I => \bfn_17_28_0_\
        );

    \I__13068\ : InMux
    port map (
            O => \N__55419\,
            I => n13015
        );

    \I__13067\ : InMux
    port map (
            O => \N__55416\,
            I => \N__55412\
        );

    \I__13066\ : InMux
    port map (
            O => \N__55415\,
            I => \N__55409\
        );

    \I__13065\ : LocalMux
    port map (
            O => \N__55412\,
            I => sweep_counter_17
        );

    \I__13064\ : LocalMux
    port map (
            O => \N__55409\,
            I => sweep_counter_17
        );

    \I__13063\ : CEMux
    port map (
            O => \N__55404\,
            I => \N__55396\
        );

    \I__13062\ : SRMux
    port map (
            O => \N__55403\,
            I => \N__55393\
        );

    \I__13061\ : CEMux
    port map (
            O => \N__55402\,
            I => \N__55390\
        );

    \I__13060\ : SRMux
    port map (
            O => \N__55401\,
            I => \N__55386\
        );

    \I__13059\ : SRMux
    port map (
            O => \N__55400\,
            I => \N__55383\
        );

    \I__13058\ : CEMux
    port map (
            O => \N__55399\,
            I => \N__55380\
        );

    \I__13057\ : LocalMux
    port map (
            O => \N__55396\,
            I => \N__55377\
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__55393\,
            I => \N__55374\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__55390\,
            I => \N__55371\
        );

    \I__13054\ : CEMux
    port map (
            O => \N__55389\,
            I => \N__55368\
        );

    \I__13053\ : LocalMux
    port map (
            O => \N__55386\,
            I => \N__55365\
        );

    \I__13052\ : LocalMux
    port map (
            O => \N__55383\,
            I => \N__55362\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__55380\,
            I => \N__55359\
        );

    \I__13050\ : Span4Mux_h
    port map (
            O => \N__55377\,
            I => \N__55354\
        );

    \I__13049\ : Span4Mux_h
    port map (
            O => \N__55374\,
            I => \N__55354\
        );

    \I__13048\ : Span4Mux_h
    port map (
            O => \N__55371\,
            I => \N__55347\
        );

    \I__13047\ : LocalMux
    port map (
            O => \N__55368\,
            I => \N__55347\
        );

    \I__13046\ : Span4Mux_h
    port map (
            O => \N__55365\,
            I => \N__55347\
        );

    \I__13045\ : Span4Mux_h
    port map (
            O => \N__55362\,
            I => \N__55344\
        );

    \I__13044\ : Odrv4
    port map (
            O => \N__55359\,
            I => n5197
        );

    \I__13043\ : Odrv4
    port map (
            O => \N__55354\,
            I => n5197
        );

    \I__13042\ : Odrv4
    port map (
            O => \N__55347\,
            I => n5197
        );

    \I__13041\ : Odrv4
    port map (
            O => \N__55344\,
            I => n5197
        );

    \I__13040\ : InMux
    port map (
            O => \N__55335\,
            I => \N__55319\
        );

    \I__13039\ : InMux
    port map (
            O => \N__55334\,
            I => \N__55316\
        );

    \I__13038\ : InMux
    port map (
            O => \N__55333\,
            I => \N__55311\
        );

    \I__13037\ : InMux
    port map (
            O => \N__55332\,
            I => \N__55311\
        );

    \I__13036\ : InMux
    port map (
            O => \N__55331\,
            I => \N__55301\
        );

    \I__13035\ : InMux
    port map (
            O => \N__55330\,
            I => \N__55301\
        );

    \I__13034\ : InMux
    port map (
            O => \N__55329\,
            I => \N__55298\
        );

    \I__13033\ : InMux
    port map (
            O => \N__55328\,
            I => \N__55291\
        );

    \I__13032\ : InMux
    port map (
            O => \N__55327\,
            I => \N__55291\
        );

    \I__13031\ : InMux
    port map (
            O => \N__55326\,
            I => \N__55291\
        );

    \I__13030\ : InMux
    port map (
            O => \N__55325\,
            I => \N__55284\
        );

    \I__13029\ : InMux
    port map (
            O => \N__55324\,
            I => \N__55284\
        );

    \I__13028\ : InMux
    port map (
            O => \N__55323\,
            I => \N__55284\
        );

    \I__13027\ : InMux
    port map (
            O => \N__55322\,
            I => \N__55281\
        );

    \I__13026\ : LocalMux
    port map (
            O => \N__55319\,
            I => \N__55278\
        );

    \I__13025\ : LocalMux
    port map (
            O => \N__55316\,
            I => \N__55273\
        );

    \I__13024\ : LocalMux
    port map (
            O => \N__55311\,
            I => \N__55273\
        );

    \I__13023\ : InMux
    port map (
            O => \N__55310\,
            I => \N__55264\
        );

    \I__13022\ : InMux
    port map (
            O => \N__55309\,
            I => \N__55264\
        );

    \I__13021\ : InMux
    port map (
            O => \N__55308\,
            I => \N__55264\
        );

    \I__13020\ : InMux
    port map (
            O => \N__55307\,
            I => \N__55255\
        );

    \I__13019\ : InMux
    port map (
            O => \N__55306\,
            I => \N__55255\
        );

    \I__13018\ : LocalMux
    port map (
            O => \N__55301\,
            I => \N__55252\
        );

    \I__13017\ : LocalMux
    port map (
            O => \N__55298\,
            I => \N__55245\
        );

    \I__13016\ : LocalMux
    port map (
            O => \N__55291\,
            I => \N__55245\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__55284\,
            I => \N__55245\
        );

    \I__13014\ : LocalMux
    port map (
            O => \N__55281\,
            I => \N__55242\
        );

    \I__13013\ : Span4Mux_h
    port map (
            O => \N__55278\,
            I => \N__55237\
        );

    \I__13012\ : Span4Mux_h
    port map (
            O => \N__55273\,
            I => \N__55237\
        );

    \I__13011\ : InMux
    port map (
            O => \N__55272\,
            I => \N__55232\
        );

    \I__13010\ : InMux
    port map (
            O => \N__55271\,
            I => \N__55232\
        );

    \I__13009\ : LocalMux
    port map (
            O => \N__55264\,
            I => \N__55229\
        );

    \I__13008\ : InMux
    port map (
            O => \N__55263\,
            I => \N__55224\
        );

    \I__13007\ : InMux
    port map (
            O => \N__55262\,
            I => \N__55224\
        );

    \I__13006\ : InMux
    port map (
            O => \N__55261\,
            I => \N__55221\
        );

    \I__13005\ : InMux
    port map (
            O => \N__55260\,
            I => \N__55218\
        );

    \I__13004\ : LocalMux
    port map (
            O => \N__55255\,
            I => \N__55207\
        );

    \I__13003\ : Span4Mux_v
    port map (
            O => \N__55252\,
            I => \N__55207\
        );

    \I__13002\ : Span4Mux_v
    port map (
            O => \N__55245\,
            I => \N__55207\
        );

    \I__13001\ : Span4Mux_v
    port map (
            O => \N__55242\,
            I => \N__55207\
        );

    \I__13000\ : Span4Mux_v
    port map (
            O => \N__55237\,
            I => \N__55207\
        );

    \I__12999\ : LocalMux
    port map (
            O => \N__55232\,
            I => \N__55202\
        );

    \I__12998\ : Span4Mux_s1_v
    port map (
            O => \N__55229\,
            I => \N__55202\
        );

    \I__12997\ : LocalMux
    port map (
            O => \N__55224\,
            I => duty_23
        );

    \I__12996\ : LocalMux
    port map (
            O => \N__55221\,
            I => duty_23
        );

    \I__12995\ : LocalMux
    port map (
            O => \N__55218\,
            I => duty_23
        );

    \I__12994\ : Odrv4
    port map (
            O => \N__55207\,
            I => duty_23
        );

    \I__12993\ : Odrv4
    port map (
            O => \N__55202\,
            I => duty_23
        );

    \I__12992\ : IoInMux
    port map (
            O => \N__55191\,
            I => \N__55188\
        );

    \I__12991\ : LocalMux
    port map (
            O => \N__55188\,
            I => \N__55185\
        );

    \I__12990\ : IoSpan4Mux
    port map (
            O => \N__55185\,
            I => \N__55182\
        );

    \I__12989\ : Span4Mux_s1_v
    port map (
            O => \N__55182\,
            I => \N__55179\
        );

    \I__12988\ : Odrv4
    port map (
            O => \N__55179\,
            I => \INLB_c_0\
        );

    \I__12987\ : InMux
    port map (
            O => \N__55176\,
            I => \N__55172\
        );

    \I__12986\ : InMux
    port map (
            O => \N__55175\,
            I => \N__55169\
        );

    \I__12985\ : LocalMux
    port map (
            O => \N__55172\,
            I => sweep_counter_5
        );

    \I__12984\ : LocalMux
    port map (
            O => \N__55169\,
            I => sweep_counter_5
        );

    \I__12983\ : InMux
    port map (
            O => \N__55164\,
            I => n13003
        );

    \I__12982\ : InMux
    port map (
            O => \N__55161\,
            I => \N__55157\
        );

    \I__12981\ : InMux
    port map (
            O => \N__55160\,
            I => \N__55154\
        );

    \I__12980\ : LocalMux
    port map (
            O => \N__55157\,
            I => sweep_counter_6
        );

    \I__12979\ : LocalMux
    port map (
            O => \N__55154\,
            I => sweep_counter_6
        );

    \I__12978\ : InMux
    port map (
            O => \N__55149\,
            I => n13004
        );

    \I__12977\ : InMux
    port map (
            O => \N__55146\,
            I => \N__55142\
        );

    \I__12976\ : InMux
    port map (
            O => \N__55145\,
            I => \N__55139\
        );

    \I__12975\ : LocalMux
    port map (
            O => \N__55142\,
            I => sweep_counter_7
        );

    \I__12974\ : LocalMux
    port map (
            O => \N__55139\,
            I => sweep_counter_7
        );

    \I__12973\ : InMux
    port map (
            O => \N__55134\,
            I => n13005
        );

    \I__12972\ : InMux
    port map (
            O => \N__55131\,
            I => \N__55127\
        );

    \I__12971\ : InMux
    port map (
            O => \N__55130\,
            I => \N__55124\
        );

    \I__12970\ : LocalMux
    port map (
            O => \N__55127\,
            I => sweep_counter_8
        );

    \I__12969\ : LocalMux
    port map (
            O => \N__55124\,
            I => sweep_counter_8
        );

    \I__12968\ : InMux
    port map (
            O => \N__55119\,
            I => \bfn_17_27_0_\
        );

    \I__12967\ : InMux
    port map (
            O => \N__55116\,
            I => \N__55112\
        );

    \I__12966\ : InMux
    port map (
            O => \N__55115\,
            I => \N__55109\
        );

    \I__12965\ : LocalMux
    port map (
            O => \N__55112\,
            I => sweep_counter_9
        );

    \I__12964\ : LocalMux
    port map (
            O => \N__55109\,
            I => sweep_counter_9
        );

    \I__12963\ : InMux
    port map (
            O => \N__55104\,
            I => n13007
        );

    \I__12962\ : InMux
    port map (
            O => \N__55101\,
            I => \N__55097\
        );

    \I__12961\ : InMux
    port map (
            O => \N__55100\,
            I => \N__55094\
        );

    \I__12960\ : LocalMux
    port map (
            O => \N__55097\,
            I => sweep_counter_10
        );

    \I__12959\ : LocalMux
    port map (
            O => \N__55094\,
            I => sweep_counter_10
        );

    \I__12958\ : InMux
    port map (
            O => \N__55089\,
            I => n13008
        );

    \I__12957\ : InMux
    port map (
            O => \N__55086\,
            I => \N__55082\
        );

    \I__12956\ : InMux
    port map (
            O => \N__55085\,
            I => \N__55079\
        );

    \I__12955\ : LocalMux
    port map (
            O => \N__55082\,
            I => \N__55076\
        );

    \I__12954\ : LocalMux
    port map (
            O => \N__55079\,
            I => sweep_counter_11
        );

    \I__12953\ : Odrv4
    port map (
            O => \N__55076\,
            I => sweep_counter_11
        );

    \I__12952\ : InMux
    port map (
            O => \N__55071\,
            I => n13009
        );

    \I__12951\ : InMux
    port map (
            O => \N__55068\,
            I => \N__55064\
        );

    \I__12950\ : InMux
    port map (
            O => \N__55067\,
            I => \N__55061\
        );

    \I__12949\ : LocalMux
    port map (
            O => \N__55064\,
            I => sweep_counter_12
        );

    \I__12948\ : LocalMux
    port map (
            O => \N__55061\,
            I => sweep_counter_12
        );

    \I__12947\ : InMux
    port map (
            O => \N__55056\,
            I => n13010
        );

    \I__12946\ : InMux
    port map (
            O => \N__55053\,
            I => \N__55049\
        );

    \I__12945\ : InMux
    port map (
            O => \N__55052\,
            I => \N__55046\
        );

    \I__12944\ : LocalMux
    port map (
            O => \N__55049\,
            I => sweep_counter_13
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__55046\,
            I => sweep_counter_13
        );

    \I__12942\ : InMux
    port map (
            O => \N__55041\,
            I => n13011
        );

    \I__12941\ : CascadeMux
    port map (
            O => \N__55038\,
            I => \n5183_cascade_\
        );

    \I__12940\ : CascadeMux
    port map (
            O => \N__55035\,
            I => \N__55031\
        );

    \I__12939\ : InMux
    port map (
            O => \N__55034\,
            I => \N__55022\
        );

    \I__12938\ : InMux
    port map (
            O => \N__55031\,
            I => \N__55022\
        );

    \I__12937\ : InMux
    port map (
            O => \N__55030\,
            I => \N__55019\
        );

    \I__12936\ : InMux
    port map (
            O => \N__55029\,
            I => \N__55016\
        );

    \I__12935\ : InMux
    port map (
            O => \N__55028\,
            I => \N__55011\
        );

    \I__12934\ : InMux
    port map (
            O => \N__55027\,
            I => \N__55011\
        );

    \I__12933\ : LocalMux
    port map (
            O => \N__55022\,
            I => \N__55008\
        );

    \I__12932\ : LocalMux
    port map (
            O => \N__55019\,
            I => dti
        );

    \I__12931\ : LocalMux
    port map (
            O => \N__55016\,
            I => dti
        );

    \I__12930\ : LocalMux
    port map (
            O => \N__55011\,
            I => dti
        );

    \I__12929\ : Odrv4
    port map (
            O => \N__55008\,
            I => dti
        );

    \I__12928\ : CascadeMux
    port map (
            O => \N__54999\,
            I => \n20_adj_706_cascade_\
        );

    \I__12927\ : InMux
    port map (
            O => \N__54996\,
            I => \N__54993\
        );

    \I__12926\ : LocalMux
    port map (
            O => \N__54993\,
            I => n24_adj_704
        );

    \I__12925\ : InMux
    port map (
            O => \N__54990\,
            I => \N__54987\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__54987\,
            I => \N__54983\
        );

    \I__12923\ : InMux
    port map (
            O => \N__54986\,
            I => \N__54980\
        );

    \I__12922\ : Odrv4
    port map (
            O => \N__54983\,
            I => n13187
        );

    \I__12921\ : LocalMux
    port map (
            O => \N__54980\,
            I => n13187
        );

    \I__12920\ : InMux
    port map (
            O => \N__54975\,
            I => \N__54971\
        );

    \I__12919\ : InMux
    port map (
            O => \N__54974\,
            I => \N__54968\
        );

    \I__12918\ : LocalMux
    port map (
            O => \N__54971\,
            I => sweep_counter_0
        );

    \I__12917\ : LocalMux
    port map (
            O => \N__54968\,
            I => sweep_counter_0
        );

    \I__12916\ : InMux
    port map (
            O => \N__54963\,
            I => \bfn_17_26_0_\
        );

    \I__12915\ : InMux
    port map (
            O => \N__54960\,
            I => \N__54956\
        );

    \I__12914\ : InMux
    port map (
            O => \N__54959\,
            I => \N__54953\
        );

    \I__12913\ : LocalMux
    port map (
            O => \N__54956\,
            I => sweep_counter_1
        );

    \I__12912\ : LocalMux
    port map (
            O => \N__54953\,
            I => sweep_counter_1
        );

    \I__12911\ : InMux
    port map (
            O => \N__54948\,
            I => n12999
        );

    \I__12910\ : InMux
    port map (
            O => \N__54945\,
            I => \N__54941\
        );

    \I__12909\ : InMux
    port map (
            O => \N__54944\,
            I => \N__54938\
        );

    \I__12908\ : LocalMux
    port map (
            O => \N__54941\,
            I => sweep_counter_2
        );

    \I__12907\ : LocalMux
    port map (
            O => \N__54938\,
            I => sweep_counter_2
        );

    \I__12906\ : InMux
    port map (
            O => \N__54933\,
            I => n13000
        );

    \I__12905\ : CascadeMux
    port map (
            O => \N__54930\,
            I => \N__54926\
        );

    \I__12904\ : InMux
    port map (
            O => \N__54929\,
            I => \N__54923\
        );

    \I__12903\ : InMux
    port map (
            O => \N__54926\,
            I => \N__54920\
        );

    \I__12902\ : LocalMux
    port map (
            O => \N__54923\,
            I => sweep_counter_3
        );

    \I__12901\ : LocalMux
    port map (
            O => \N__54920\,
            I => sweep_counter_3
        );

    \I__12900\ : InMux
    port map (
            O => \N__54915\,
            I => n13001
        );

    \I__12899\ : InMux
    port map (
            O => \N__54912\,
            I => \N__54908\
        );

    \I__12898\ : InMux
    port map (
            O => \N__54911\,
            I => \N__54905\
        );

    \I__12897\ : LocalMux
    port map (
            O => \N__54908\,
            I => sweep_counter_4
        );

    \I__12896\ : LocalMux
    port map (
            O => \N__54905\,
            I => sweep_counter_4
        );

    \I__12895\ : InMux
    port map (
            O => \N__54900\,
            I => n13002
        );

    \I__12894\ : CascadeMux
    port map (
            O => \N__54897\,
            I => \n6_adj_582_cascade_\
        );

    \I__12893\ : InMux
    port map (
            O => \N__54894\,
            I => \N__54888\
        );

    \I__12892\ : InMux
    port map (
            O => \N__54893\,
            I => \N__54888\
        );

    \I__12891\ : LocalMux
    port map (
            O => \N__54888\,
            I => \N__54885\
        );

    \I__12890\ : Odrv4
    port map (
            O => \N__54885\,
            I => n14108
        );

    \I__12889\ : CascadeMux
    port map (
            O => \N__54882\,
            I => \N__54878\
        );

    \I__12888\ : InMux
    port map (
            O => \N__54881\,
            I => \N__54875\
        );

    \I__12887\ : InMux
    port map (
            O => \N__54878\,
            I => \N__54870\
        );

    \I__12886\ : LocalMux
    port map (
            O => \N__54875\,
            I => \N__54867\
        );

    \I__12885\ : InMux
    port map (
            O => \N__54874\,
            I => \N__54864\
        );

    \I__12884\ : InMux
    port map (
            O => \N__54873\,
            I => \N__54861\
        );

    \I__12883\ : LocalMux
    port map (
            O => \N__54870\,
            I => encoder0_position_target_15
        );

    \I__12882\ : Odrv12
    port map (
            O => \N__54867\,
            I => encoder0_position_target_15
        );

    \I__12881\ : LocalMux
    port map (
            O => \N__54864\,
            I => encoder0_position_target_15
        );

    \I__12880\ : LocalMux
    port map (
            O => \N__54861\,
            I => encoder0_position_target_15
        );

    \I__12879\ : CascadeMux
    port map (
            O => \N__54852\,
            I => \N__54849\
        );

    \I__12878\ : InMux
    port map (
            O => \N__54849\,
            I => \N__54844\
        );

    \I__12877\ : InMux
    port map (
            O => \N__54848\,
            I => \N__54841\
        );

    \I__12876\ : CascadeMux
    port map (
            O => \N__54847\,
            I => \N__54838\
        );

    \I__12875\ : LocalMux
    port map (
            O => \N__54844\,
            I => \N__54835\
        );

    \I__12874\ : LocalMux
    port map (
            O => \N__54841\,
            I => \N__54831\
        );

    \I__12873\ : InMux
    port map (
            O => \N__54838\,
            I => \N__54828\
        );

    \I__12872\ : Span4Mux_h
    port map (
            O => \N__54835\,
            I => \N__54825\
        );

    \I__12871\ : InMux
    port map (
            O => \N__54834\,
            I => \N__54822\
        );

    \I__12870\ : Span4Mux_h
    port map (
            O => \N__54831\,
            I => \N__54819\
        );

    \I__12869\ : LocalMux
    port map (
            O => \N__54828\,
            I => encoder0_position_target_21
        );

    \I__12868\ : Odrv4
    port map (
            O => \N__54825\,
            I => encoder0_position_target_21
        );

    \I__12867\ : LocalMux
    port map (
            O => \N__54822\,
            I => encoder0_position_target_21
        );

    \I__12866\ : Odrv4
    port map (
            O => \N__54819\,
            I => encoder0_position_target_21
        );

    \I__12865\ : CascadeMux
    port map (
            O => \N__54810\,
            I => \N__54807\
        );

    \I__12864\ : InMux
    port map (
            O => \N__54807\,
            I => \N__54802\
        );

    \I__12863\ : InMux
    port map (
            O => \N__54806\,
            I => \N__54798\
        );

    \I__12862\ : CascadeMux
    port map (
            O => \N__54805\,
            I => \N__54795\
        );

    \I__12861\ : LocalMux
    port map (
            O => \N__54802\,
            I => \N__54792\
        );

    \I__12860\ : CascadeMux
    port map (
            O => \N__54801\,
            I => \N__54789\
        );

    \I__12859\ : LocalMux
    port map (
            O => \N__54798\,
            I => \N__54786\
        );

    \I__12858\ : InMux
    port map (
            O => \N__54795\,
            I => \N__54783\
        );

    \I__12857\ : Span4Mux_v
    port map (
            O => \N__54792\,
            I => \N__54780\
        );

    \I__12856\ : InMux
    port map (
            O => \N__54789\,
            I => \N__54777\
        );

    \I__12855\ : Span4Mux_h
    port map (
            O => \N__54786\,
            I => \N__54774\
        );

    \I__12854\ : LocalMux
    port map (
            O => \N__54783\,
            I => encoder0_position_target_19
        );

    \I__12853\ : Odrv4
    port map (
            O => \N__54780\,
            I => encoder0_position_target_19
        );

    \I__12852\ : LocalMux
    port map (
            O => \N__54777\,
            I => encoder0_position_target_19
        );

    \I__12851\ : Odrv4
    port map (
            O => \N__54774\,
            I => encoder0_position_target_19
        );

    \I__12850\ : CascadeMux
    port map (
            O => \N__54765\,
            I => \N__54759\
        );

    \I__12849\ : InMux
    port map (
            O => \N__54764\,
            I => \N__54756\
        );

    \I__12848\ : InMux
    port map (
            O => \N__54763\,
            I => \N__54752\
        );

    \I__12847\ : InMux
    port map (
            O => \N__54762\,
            I => \N__54749\
        );

    \I__12846\ : InMux
    port map (
            O => \N__54759\,
            I => \N__54745\
        );

    \I__12845\ : LocalMux
    port map (
            O => \N__54756\,
            I => \N__54742\
        );

    \I__12844\ : InMux
    port map (
            O => \N__54755\,
            I => \N__54739\
        );

    \I__12843\ : LocalMux
    port map (
            O => \N__54752\,
            I => \N__54736\
        );

    \I__12842\ : LocalMux
    port map (
            O => \N__54749\,
            I => \N__54733\
        );

    \I__12841\ : InMux
    port map (
            O => \N__54748\,
            I => \N__54730\
        );

    \I__12840\ : LocalMux
    port map (
            O => \N__54745\,
            I => \N__54725\
        );

    \I__12839\ : Span4Mux_h
    port map (
            O => \N__54742\,
            I => \N__54725\
        );

    \I__12838\ : LocalMux
    port map (
            O => \N__54739\,
            I => encoder0_position_target_23
        );

    \I__12837\ : Odrv12
    port map (
            O => \N__54736\,
            I => encoder0_position_target_23
        );

    \I__12836\ : Odrv4
    port map (
            O => \N__54733\,
            I => encoder0_position_target_23
        );

    \I__12835\ : LocalMux
    port map (
            O => \N__54730\,
            I => encoder0_position_target_23
        );

    \I__12834\ : Odrv4
    port map (
            O => \N__54725\,
            I => encoder0_position_target_23
        );

    \I__12833\ : InMux
    port map (
            O => \N__54714\,
            I => \N__54711\
        );

    \I__12832\ : LocalMux
    port map (
            O => \N__54711\,
            I => \N__54708\
        );

    \I__12831\ : Odrv4
    port map (
            O => \N__54708\,
            I => n24_adj_699
        );

    \I__12830\ : InMux
    port map (
            O => \N__54705\,
            I => \N__54702\
        );

    \I__12829\ : LocalMux
    port map (
            O => \N__54702\,
            I => n16_adj_707
        );

    \I__12828\ : CascadeMux
    port map (
            O => \N__54699\,
            I => \N__54694\
        );

    \I__12827\ : CascadeMux
    port map (
            O => \N__54698\,
            I => \N__54690\
        );

    \I__12826\ : InMux
    port map (
            O => \N__54697\,
            I => \N__54685\
        );

    \I__12825\ : InMux
    port map (
            O => \N__54694\,
            I => \N__54679\
        );

    \I__12824\ : InMux
    port map (
            O => \N__54693\,
            I => \N__54679\
        );

    \I__12823\ : InMux
    port map (
            O => \N__54690\,
            I => \N__54672\
        );

    \I__12822\ : InMux
    port map (
            O => \N__54689\,
            I => \N__54672\
        );

    \I__12821\ : InMux
    port map (
            O => \N__54688\,
            I => \N__54672\
        );

    \I__12820\ : LocalMux
    port map (
            O => \N__54685\,
            I => \N__54667\
        );

    \I__12819\ : InMux
    port map (
            O => \N__54684\,
            I => \N__54664\
        );

    \I__12818\ : LocalMux
    port map (
            O => \N__54679\,
            I => \N__54659\
        );

    \I__12817\ : LocalMux
    port map (
            O => \N__54672\,
            I => \N__54659\
        );

    \I__12816\ : InMux
    port map (
            O => \N__54671\,
            I => \N__54656\
        );

    \I__12815\ : InMux
    port map (
            O => \N__54670\,
            I => \N__54653\
        );

    \I__12814\ : Odrv4
    port map (
            O => \N__54667\,
            I => commutation_state_prev_0
        );

    \I__12813\ : LocalMux
    port map (
            O => \N__54664\,
            I => commutation_state_prev_0
        );

    \I__12812\ : Odrv4
    port map (
            O => \N__54659\,
            I => commutation_state_prev_0
        );

    \I__12811\ : LocalMux
    port map (
            O => \N__54656\,
            I => commutation_state_prev_0
        );

    \I__12810\ : LocalMux
    port map (
            O => \N__54653\,
            I => commutation_state_prev_0
        );

    \I__12809\ : CascadeMux
    port map (
            O => \N__54642\,
            I => \dti_N_333_cascade_\
        );

    \I__12808\ : CascadeMux
    port map (
            O => \N__54639\,
            I => \N__54631\
        );

    \I__12807\ : CascadeMux
    port map (
            O => \N__54638\,
            I => \N__54628\
        );

    \I__12806\ : CascadeMux
    port map (
            O => \N__54637\,
            I => \N__54625\
        );

    \I__12805\ : CascadeMux
    port map (
            O => \N__54636\,
            I => \N__54620\
        );

    \I__12804\ : InMux
    port map (
            O => \N__54635\,
            I => \N__54617\
        );

    \I__12803\ : InMux
    port map (
            O => \N__54634\,
            I => \N__54610\
        );

    \I__12802\ : InMux
    port map (
            O => \N__54631\,
            I => \N__54610\
        );

    \I__12801\ : InMux
    port map (
            O => \N__54628\,
            I => \N__54610\
        );

    \I__12800\ : InMux
    port map (
            O => \N__54625\,
            I => \N__54605\
        );

    \I__12799\ : InMux
    port map (
            O => \N__54624\,
            I => \N__54605\
        );

    \I__12798\ : InMux
    port map (
            O => \N__54623\,
            I => \N__54602\
        );

    \I__12797\ : InMux
    port map (
            O => \N__54620\,
            I => \N__54599\
        );

    \I__12796\ : LocalMux
    port map (
            O => \N__54617\,
            I => \N__54596\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__54610\,
            I => \N__54591\
        );

    \I__12794\ : LocalMux
    port map (
            O => \N__54605\,
            I => \N__54591\
        );

    \I__12793\ : LocalMux
    port map (
            O => \N__54602\,
            I => n4_adj_716
        );

    \I__12792\ : LocalMux
    port map (
            O => \N__54599\,
            I => n4_adj_716
        );

    \I__12791\ : Odrv4
    port map (
            O => \N__54596\,
            I => n4_adj_716
        );

    \I__12790\ : Odrv4
    port map (
            O => \N__54591\,
            I => n4_adj_716
        );

    \I__12789\ : CEMux
    port map (
            O => \N__54582\,
            I => \N__54579\
        );

    \I__12788\ : LocalMux
    port map (
            O => \N__54579\,
            I => n5169
        );

    \I__12787\ : CascadeMux
    port map (
            O => \N__54576\,
            I => \N__54573\
        );

    \I__12786\ : InMux
    port map (
            O => \N__54573\,
            I => \N__54570\
        );

    \I__12785\ : LocalMux
    port map (
            O => \N__54570\,
            I => n1377
        );

    \I__12784\ : InMux
    port map (
            O => \N__54567\,
            I => \N__54561\
        );

    \I__12783\ : InMux
    port map (
            O => \N__54566\,
            I => \N__54558\
        );

    \I__12782\ : InMux
    port map (
            O => \N__54565\,
            I => \N__54553\
        );

    \I__12781\ : InMux
    port map (
            O => \N__54564\,
            I => \N__54553\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__54561\,
            I => n5119
        );

    \I__12779\ : LocalMux
    port map (
            O => \N__54558\,
            I => n5119
        );

    \I__12778\ : LocalMux
    port map (
            O => \N__54553\,
            I => n5119
        );

    \I__12777\ : CascadeMux
    port map (
            O => \N__54546\,
            I => \N__54540\
        );

    \I__12776\ : CascadeMux
    port map (
            O => \N__54545\,
            I => \N__54536\
        );

    \I__12775\ : CascadeMux
    port map (
            O => \N__54544\,
            I => \N__54531\
        );

    \I__12774\ : CascadeMux
    port map (
            O => \N__54543\,
            I => \N__54523\
        );

    \I__12773\ : InMux
    port map (
            O => \N__54540\,
            I => \N__54491\
        );

    \I__12772\ : InMux
    port map (
            O => \N__54539\,
            I => \N__54491\
        );

    \I__12771\ : InMux
    port map (
            O => \N__54536\,
            I => \N__54491\
        );

    \I__12770\ : InMux
    port map (
            O => \N__54535\,
            I => \N__54491\
        );

    \I__12769\ : InMux
    port map (
            O => \N__54534\,
            I => \N__54491\
        );

    \I__12768\ : InMux
    port map (
            O => \N__54531\,
            I => \N__54484\
        );

    \I__12767\ : InMux
    port map (
            O => \N__54530\,
            I => \N__54484\
        );

    \I__12766\ : InMux
    port map (
            O => \N__54529\,
            I => \N__54484\
        );

    \I__12765\ : InMux
    port map (
            O => \N__54528\,
            I => \N__54477\
        );

    \I__12764\ : InMux
    port map (
            O => \N__54527\,
            I => \N__54477\
        );

    \I__12763\ : InMux
    port map (
            O => \N__54526\,
            I => \N__54477\
        );

    \I__12762\ : InMux
    port map (
            O => \N__54523\,
            I => \N__54466\
        );

    \I__12761\ : InMux
    port map (
            O => \N__54522\,
            I => \N__54466\
        );

    \I__12760\ : InMux
    port map (
            O => \N__54521\,
            I => \N__54466\
        );

    \I__12759\ : InMux
    port map (
            O => \N__54520\,
            I => \N__54466\
        );

    \I__12758\ : InMux
    port map (
            O => \N__54519\,
            I => \N__54466\
        );

    \I__12757\ : CascadeMux
    port map (
            O => \N__54518\,
            I => \N__54462\
        );

    \I__12756\ : CascadeMux
    port map (
            O => \N__54517\,
            I => \N__54452\
        );

    \I__12755\ : CascadeMux
    port map (
            O => \N__54516\,
            I => \N__54449\
        );

    \I__12754\ : CascadeMux
    port map (
            O => \N__54515\,
            I => \N__54446\
        );

    \I__12753\ : CascadeMux
    port map (
            O => \N__54514\,
            I => \N__54443\
        );

    \I__12752\ : CascadeMux
    port map (
            O => \N__54513\,
            I => \N__54440\
        );

    \I__12751\ : CascadeMux
    port map (
            O => \N__54512\,
            I => \N__54437\
        );

    \I__12750\ : CascadeMux
    port map (
            O => \N__54511\,
            I => \N__54434\
        );

    \I__12749\ : CascadeMux
    port map (
            O => \N__54510\,
            I => \N__54431\
        );

    \I__12748\ : CascadeMux
    port map (
            O => \N__54509\,
            I => \N__54428\
        );

    \I__12747\ : CascadeMux
    port map (
            O => \N__54508\,
            I => \N__54425\
        );

    \I__12746\ : CascadeMux
    port map (
            O => \N__54507\,
            I => \N__54419\
        );

    \I__12745\ : CascadeMux
    port map (
            O => \N__54506\,
            I => \N__54410\
        );

    \I__12744\ : CascadeMux
    port map (
            O => \N__54505\,
            I => \N__54407\
        );

    \I__12743\ : CascadeMux
    port map (
            O => \N__54504\,
            I => \N__54396\
        );

    \I__12742\ : CascadeMux
    port map (
            O => \N__54503\,
            I => \N__54392\
        );

    \I__12741\ : CascadeMux
    port map (
            O => \N__54502\,
            I => \N__54386\
        );

    \I__12740\ : LocalMux
    port map (
            O => \N__54491\,
            I => \N__54381\
        );

    \I__12739\ : LocalMux
    port map (
            O => \N__54484\,
            I => \N__54381\
        );

    \I__12738\ : LocalMux
    port map (
            O => \N__54477\,
            I => \N__54376\
        );

    \I__12737\ : LocalMux
    port map (
            O => \N__54466\,
            I => \N__54376\
        );

    \I__12736\ : InMux
    port map (
            O => \N__54465\,
            I => \N__54371\
        );

    \I__12735\ : InMux
    port map (
            O => \N__54462\,
            I => \N__54371\
        );

    \I__12734\ : InMux
    port map (
            O => \N__54461\,
            I => \N__54366\
        );

    \I__12733\ : InMux
    port map (
            O => \N__54460\,
            I => \N__54366\
        );

    \I__12732\ : CascadeMux
    port map (
            O => \N__54459\,
            I => \N__54362\
        );

    \I__12731\ : CascadeMux
    port map (
            O => \N__54458\,
            I => \N__54355\
        );

    \I__12730\ : CascadeMux
    port map (
            O => \N__54457\,
            I => \N__54347\
        );

    \I__12729\ : CascadeMux
    port map (
            O => \N__54456\,
            I => \N__54342\
        );

    \I__12728\ : InMux
    port map (
            O => \N__54455\,
            I => \N__54337\
        );

    \I__12727\ : InMux
    port map (
            O => \N__54452\,
            I => \N__54337\
        );

    \I__12726\ : InMux
    port map (
            O => \N__54449\,
            I => \N__54334\
        );

    \I__12725\ : InMux
    port map (
            O => \N__54446\,
            I => \N__54325\
        );

    \I__12724\ : InMux
    port map (
            O => \N__54443\,
            I => \N__54325\
        );

    \I__12723\ : InMux
    port map (
            O => \N__54440\,
            I => \N__54325\
        );

    \I__12722\ : InMux
    port map (
            O => \N__54437\,
            I => \N__54325\
        );

    \I__12721\ : InMux
    port map (
            O => \N__54434\,
            I => \N__54316\
        );

    \I__12720\ : InMux
    port map (
            O => \N__54431\,
            I => \N__54316\
        );

    \I__12719\ : InMux
    port map (
            O => \N__54428\,
            I => \N__54316\
        );

    \I__12718\ : InMux
    port map (
            O => \N__54425\,
            I => \N__54316\
        );

    \I__12717\ : InMux
    port map (
            O => \N__54424\,
            I => \N__54309\
        );

    \I__12716\ : InMux
    port map (
            O => \N__54423\,
            I => \N__54309\
        );

    \I__12715\ : InMux
    port map (
            O => \N__54422\,
            I => \N__54309\
        );

    \I__12714\ : InMux
    port map (
            O => \N__54419\,
            I => \N__54298\
        );

    \I__12713\ : InMux
    port map (
            O => \N__54418\,
            I => \N__54298\
        );

    \I__12712\ : InMux
    port map (
            O => \N__54417\,
            I => \N__54298\
        );

    \I__12711\ : InMux
    port map (
            O => \N__54416\,
            I => \N__54298\
        );

    \I__12710\ : InMux
    port map (
            O => \N__54415\,
            I => \N__54298\
        );

    \I__12709\ : InMux
    port map (
            O => \N__54414\,
            I => \N__54259\
        );

    \I__12708\ : InMux
    port map (
            O => \N__54413\,
            I => \N__54252\
        );

    \I__12707\ : InMux
    port map (
            O => \N__54410\,
            I => \N__54252\
        );

    \I__12706\ : InMux
    port map (
            O => \N__54407\,
            I => \N__54252\
        );

    \I__12705\ : InMux
    port map (
            O => \N__54406\,
            I => \N__54249\
        );

    \I__12704\ : InMux
    port map (
            O => \N__54405\,
            I => \N__54242\
        );

    \I__12703\ : InMux
    port map (
            O => \N__54404\,
            I => \N__54242\
        );

    \I__12702\ : InMux
    port map (
            O => \N__54403\,
            I => \N__54242\
        );

    \I__12701\ : InMux
    port map (
            O => \N__54402\,
            I => \N__54239\
        );

    \I__12700\ : InMux
    port map (
            O => \N__54401\,
            I => \N__54232\
        );

    \I__12699\ : InMux
    port map (
            O => \N__54400\,
            I => \N__54232\
        );

    \I__12698\ : InMux
    port map (
            O => \N__54399\,
            I => \N__54232\
        );

    \I__12697\ : InMux
    port map (
            O => \N__54396\,
            I => \N__54219\
        );

    \I__12696\ : InMux
    port map (
            O => \N__54395\,
            I => \N__54219\
        );

    \I__12695\ : InMux
    port map (
            O => \N__54392\,
            I => \N__54219\
        );

    \I__12694\ : InMux
    port map (
            O => \N__54391\,
            I => \N__54219\
        );

    \I__12693\ : InMux
    port map (
            O => \N__54390\,
            I => \N__54219\
        );

    \I__12692\ : InMux
    port map (
            O => \N__54389\,
            I => \N__54219\
        );

    \I__12691\ : InMux
    port map (
            O => \N__54386\,
            I => \N__54216\
        );

    \I__12690\ : Span4Mux_s3_h
    port map (
            O => \N__54381\,
            I => \N__54207\
        );

    \I__12689\ : Span4Mux_v
    port map (
            O => \N__54376\,
            I => \N__54207\
        );

    \I__12688\ : LocalMux
    port map (
            O => \N__54371\,
            I => \N__54207\
        );

    \I__12687\ : LocalMux
    port map (
            O => \N__54366\,
            I => \N__54207\
        );

    \I__12686\ : InMux
    port map (
            O => \N__54365\,
            I => \N__54202\
        );

    \I__12685\ : InMux
    port map (
            O => \N__54362\,
            I => \N__54202\
        );

    \I__12684\ : CascadeMux
    port map (
            O => \N__54361\,
            I => \N__54198\
        );

    \I__12683\ : CascadeMux
    port map (
            O => \N__54360\,
            I => \N__54194\
        );

    \I__12682\ : CascadeMux
    port map (
            O => \N__54359\,
            I => \N__54191\
        );

    \I__12681\ : InMux
    port map (
            O => \N__54358\,
            I => \N__54169\
        );

    \I__12680\ : InMux
    port map (
            O => \N__54355\,
            I => \N__54169\
        );

    \I__12679\ : InMux
    port map (
            O => \N__54354\,
            I => \N__54169\
        );

    \I__12678\ : InMux
    port map (
            O => \N__54353\,
            I => \N__54164\
        );

    \I__12677\ : InMux
    port map (
            O => \N__54352\,
            I => \N__54164\
        );

    \I__12676\ : InMux
    port map (
            O => \N__54351\,
            I => \N__54151\
        );

    \I__12675\ : InMux
    port map (
            O => \N__54350\,
            I => \N__54151\
        );

    \I__12674\ : InMux
    port map (
            O => \N__54347\,
            I => \N__54151\
        );

    \I__12673\ : InMux
    port map (
            O => \N__54346\,
            I => \N__54151\
        );

    \I__12672\ : InMux
    port map (
            O => \N__54345\,
            I => \N__54151\
        );

    \I__12671\ : InMux
    port map (
            O => \N__54342\,
            I => \N__54151\
        );

    \I__12670\ : LocalMux
    port map (
            O => \N__54337\,
            I => \N__54138\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__54334\,
            I => \N__54138\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__54325\,
            I => \N__54138\
        );

    \I__12667\ : LocalMux
    port map (
            O => \N__54316\,
            I => \N__54138\
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__54309\,
            I => \N__54138\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__54298\,
            I => \N__54138\
        );

    \I__12664\ : InMux
    port map (
            O => \N__54297\,
            I => \N__54135\
        );

    \I__12663\ : CascadeMux
    port map (
            O => \N__54296\,
            I => \N__54131\
        );

    \I__12662\ : CascadeMux
    port map (
            O => \N__54295\,
            I => \N__54128\
        );

    \I__12661\ : CascadeMux
    port map (
            O => \N__54294\,
            I => \N__54125\
        );

    \I__12660\ : CascadeMux
    port map (
            O => \N__54293\,
            I => \N__54122\
        );

    \I__12659\ : CascadeMux
    port map (
            O => \N__54292\,
            I => \N__54118\
        );

    \I__12658\ : CascadeMux
    port map (
            O => \N__54291\,
            I => \N__54115\
        );

    \I__12657\ : CascadeMux
    port map (
            O => \N__54290\,
            I => \N__54112\
        );

    \I__12656\ : CascadeMux
    port map (
            O => \N__54289\,
            I => \N__54109\
        );

    \I__12655\ : CascadeMux
    port map (
            O => \N__54288\,
            I => \N__54106\
        );

    \I__12654\ : CascadeMux
    port map (
            O => \N__54287\,
            I => \N__54103\
        );

    \I__12653\ : CascadeMux
    port map (
            O => \N__54286\,
            I => \N__54099\
        );

    \I__12652\ : CascadeMux
    port map (
            O => \N__54285\,
            I => \N__54088\
        );

    \I__12651\ : CascadeMux
    port map (
            O => \N__54284\,
            I => \N__54085\
        );

    \I__12650\ : CascadeMux
    port map (
            O => \N__54283\,
            I => \N__54082\
        );

    \I__12649\ : CascadeMux
    port map (
            O => \N__54282\,
            I => \N__54075\
        );

    \I__12648\ : CascadeMux
    port map (
            O => \N__54281\,
            I => \N__54072\
        );

    \I__12647\ : CascadeMux
    port map (
            O => \N__54280\,
            I => \N__54069\
        );

    \I__12646\ : CascadeMux
    port map (
            O => \N__54279\,
            I => \N__54066\
        );

    \I__12645\ : CascadeMux
    port map (
            O => \N__54278\,
            I => \N__54063\
        );

    \I__12644\ : CascadeMux
    port map (
            O => \N__54277\,
            I => \N__54059\
        );

    \I__12643\ : CascadeMux
    port map (
            O => \N__54276\,
            I => \N__54056\
        );

    \I__12642\ : CascadeMux
    port map (
            O => \N__54275\,
            I => \N__54053\
        );

    \I__12641\ : CascadeMux
    port map (
            O => \N__54274\,
            I => \N__54049\
        );

    \I__12640\ : CascadeMux
    port map (
            O => \N__54273\,
            I => \N__54046\
        );

    \I__12639\ : CascadeMux
    port map (
            O => \N__54272\,
            I => \N__54043\
        );

    \I__12638\ : CascadeMux
    port map (
            O => \N__54271\,
            I => \N__54040\
        );

    \I__12637\ : CascadeMux
    port map (
            O => \N__54270\,
            I => \N__54037\
        );

    \I__12636\ : CascadeMux
    port map (
            O => \N__54269\,
            I => \N__54034\
        );

    \I__12635\ : CascadeMux
    port map (
            O => \N__54268\,
            I => \N__54031\
        );

    \I__12634\ : CascadeMux
    port map (
            O => \N__54267\,
            I => \N__54028\
        );

    \I__12633\ : CascadeMux
    port map (
            O => \N__54266\,
            I => \N__54025\
        );

    \I__12632\ : CascadeMux
    port map (
            O => \N__54265\,
            I => \N__54022\
        );

    \I__12631\ : CascadeMux
    port map (
            O => \N__54264\,
            I => \N__54019\
        );

    \I__12630\ : CascadeMux
    port map (
            O => \N__54263\,
            I => \N__54015\
        );

    \I__12629\ : CascadeMux
    port map (
            O => \N__54262\,
            I => \N__54012\
        );

    \I__12628\ : LocalMux
    port map (
            O => \N__54259\,
            I => \N__53968\
        );

    \I__12627\ : LocalMux
    port map (
            O => \N__54252\,
            I => \N__53968\
        );

    \I__12626\ : LocalMux
    port map (
            O => \N__54249\,
            I => \N__53968\
        );

    \I__12625\ : LocalMux
    port map (
            O => \N__54242\,
            I => \N__53968\
        );

    \I__12624\ : LocalMux
    port map (
            O => \N__54239\,
            I => \N__53968\
        );

    \I__12623\ : LocalMux
    port map (
            O => \N__54232\,
            I => \N__53968\
        );

    \I__12622\ : LocalMux
    port map (
            O => \N__54219\,
            I => \N__53963\
        );

    \I__12621\ : LocalMux
    port map (
            O => \N__54216\,
            I => \N__53963\
        );

    \I__12620\ : Span4Mux_h
    port map (
            O => \N__54207\,
            I => \N__53958\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__54202\,
            I => \N__53958\
        );

    \I__12618\ : InMux
    port map (
            O => \N__54201\,
            I => \N__53955\
        );

    \I__12617\ : InMux
    port map (
            O => \N__54198\,
            I => \N__53948\
        );

    \I__12616\ : InMux
    port map (
            O => \N__54197\,
            I => \N__53948\
        );

    \I__12615\ : InMux
    port map (
            O => \N__54194\,
            I => \N__53948\
        );

    \I__12614\ : InMux
    port map (
            O => \N__54191\,
            I => \N__53943\
        );

    \I__12613\ : InMux
    port map (
            O => \N__54190\,
            I => \N__53943\
        );

    \I__12612\ : InMux
    port map (
            O => \N__54189\,
            I => \N__53938\
        );

    \I__12611\ : InMux
    port map (
            O => \N__54188\,
            I => \N__53938\
        );

    \I__12610\ : CascadeMux
    port map (
            O => \N__54187\,
            I => \N__53930\
        );

    \I__12609\ : CascadeMux
    port map (
            O => \N__54186\,
            I => \N__53927\
        );

    \I__12608\ : CascadeMux
    port map (
            O => \N__54185\,
            I => \N__53922\
        );

    \I__12607\ : CascadeMux
    port map (
            O => \N__54184\,
            I => \N__53918\
        );

    \I__12606\ : CascadeMux
    port map (
            O => \N__54183\,
            I => \N__53912\
        );

    \I__12605\ : CascadeMux
    port map (
            O => \N__54182\,
            I => \N__53909\
        );

    \I__12604\ : CascadeMux
    port map (
            O => \N__54181\,
            I => \N__53906\
        );

    \I__12603\ : CascadeMux
    port map (
            O => \N__54180\,
            I => \N__53899\
        );

    \I__12602\ : CascadeMux
    port map (
            O => \N__54179\,
            I => \N__53893\
        );

    \I__12601\ : CascadeMux
    port map (
            O => \N__54178\,
            I => \N__53885\
        );

    \I__12600\ : CascadeMux
    port map (
            O => \N__54177\,
            I => \N__53882\
        );

    \I__12599\ : CascadeMux
    port map (
            O => \N__54176\,
            I => \N__53879\
        );

    \I__12598\ : LocalMux
    port map (
            O => \N__54169\,
            I => \N__53872\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__54164\,
            I => \N__53872\
        );

    \I__12596\ : LocalMux
    port map (
            O => \N__54151\,
            I => \N__53872\
        );

    \I__12595\ : Span4Mux_v
    port map (
            O => \N__54138\,
            I => \N__53867\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__54135\,
            I => \N__53867\
        );

    \I__12593\ : InMux
    port map (
            O => \N__54134\,
            I => \N__53860\
        );

    \I__12592\ : InMux
    port map (
            O => \N__54131\,
            I => \N__53860\
        );

    \I__12591\ : InMux
    port map (
            O => \N__54128\,
            I => \N__53860\
        );

    \I__12590\ : InMux
    port map (
            O => \N__54125\,
            I => \N__53853\
        );

    \I__12589\ : InMux
    port map (
            O => \N__54122\,
            I => \N__53853\
        );

    \I__12588\ : InMux
    port map (
            O => \N__54121\,
            I => \N__53853\
        );

    \I__12587\ : InMux
    port map (
            O => \N__54118\,
            I => \N__53846\
        );

    \I__12586\ : InMux
    port map (
            O => \N__54115\,
            I => \N__53846\
        );

    \I__12585\ : InMux
    port map (
            O => \N__54112\,
            I => \N__53846\
        );

    \I__12584\ : InMux
    port map (
            O => \N__54109\,
            I => \N__53835\
        );

    \I__12583\ : InMux
    port map (
            O => \N__54106\,
            I => \N__53835\
        );

    \I__12582\ : InMux
    port map (
            O => \N__54103\,
            I => \N__53835\
        );

    \I__12581\ : InMux
    port map (
            O => \N__54102\,
            I => \N__53835\
        );

    \I__12580\ : InMux
    port map (
            O => \N__54099\,
            I => \N__53835\
        );

    \I__12579\ : InMux
    port map (
            O => \N__54098\,
            I => \N__53828\
        );

    \I__12578\ : InMux
    port map (
            O => \N__54097\,
            I => \N__53828\
        );

    \I__12577\ : InMux
    port map (
            O => \N__54096\,
            I => \N__53828\
        );

    \I__12576\ : CascadeMux
    port map (
            O => \N__54095\,
            I => \N__53825\
        );

    \I__12575\ : CascadeMux
    port map (
            O => \N__54094\,
            I => \N__53822\
        );

    \I__12574\ : CascadeMux
    port map (
            O => \N__54093\,
            I => \N__53819\
        );

    \I__12573\ : CascadeMux
    port map (
            O => \N__54092\,
            I => \N__53815\
        );

    \I__12572\ : InMux
    port map (
            O => \N__54091\,
            I => \N__53802\
        );

    \I__12571\ : InMux
    port map (
            O => \N__54088\,
            I => \N__53802\
        );

    \I__12570\ : InMux
    port map (
            O => \N__54085\,
            I => \N__53797\
        );

    \I__12569\ : InMux
    port map (
            O => \N__54082\,
            I => \N__53797\
        );

    \I__12568\ : CascadeMux
    port map (
            O => \N__54081\,
            I => \N__53794\
        );

    \I__12567\ : CascadeMux
    port map (
            O => \N__54080\,
            I => \N__53789\
        );

    \I__12566\ : CascadeMux
    port map (
            O => \N__54079\,
            I => \N__53786\
        );

    \I__12565\ : InMux
    port map (
            O => \N__54078\,
            I => \N__53776\
        );

    \I__12564\ : InMux
    port map (
            O => \N__54075\,
            I => \N__53776\
        );

    \I__12563\ : InMux
    port map (
            O => \N__54072\,
            I => \N__53776\
        );

    \I__12562\ : InMux
    port map (
            O => \N__54069\,
            I => \N__53769\
        );

    \I__12561\ : InMux
    port map (
            O => \N__54066\,
            I => \N__53769\
        );

    \I__12560\ : InMux
    port map (
            O => \N__54063\,
            I => \N__53769\
        );

    \I__12559\ : InMux
    port map (
            O => \N__54062\,
            I => \N__53766\
        );

    \I__12558\ : InMux
    port map (
            O => \N__54059\,
            I => \N__53758\
        );

    \I__12557\ : InMux
    port map (
            O => \N__54056\,
            I => \N__53758\
        );

    \I__12556\ : InMux
    port map (
            O => \N__54053\,
            I => \N__53747\
        );

    \I__12555\ : InMux
    port map (
            O => \N__54052\,
            I => \N__53747\
        );

    \I__12554\ : InMux
    port map (
            O => \N__54049\,
            I => \N__53747\
        );

    \I__12553\ : InMux
    port map (
            O => \N__54046\,
            I => \N__53747\
        );

    \I__12552\ : InMux
    port map (
            O => \N__54043\,
            I => \N__53747\
        );

    \I__12551\ : InMux
    port map (
            O => \N__54040\,
            I => \N__53738\
        );

    \I__12550\ : InMux
    port map (
            O => \N__54037\,
            I => \N__53738\
        );

    \I__12549\ : InMux
    port map (
            O => \N__54034\,
            I => \N__53738\
        );

    \I__12548\ : InMux
    port map (
            O => \N__54031\,
            I => \N__53738\
        );

    \I__12547\ : InMux
    port map (
            O => \N__54028\,
            I => \N__53729\
        );

    \I__12546\ : InMux
    port map (
            O => \N__54025\,
            I => \N__53729\
        );

    \I__12545\ : InMux
    port map (
            O => \N__54022\,
            I => \N__53729\
        );

    \I__12544\ : InMux
    port map (
            O => \N__54019\,
            I => \N__53729\
        );

    \I__12543\ : InMux
    port map (
            O => \N__54018\,
            I => \N__53718\
        );

    \I__12542\ : InMux
    port map (
            O => \N__54015\,
            I => \N__53718\
        );

    \I__12541\ : InMux
    port map (
            O => \N__54012\,
            I => \N__53718\
        );

    \I__12540\ : InMux
    port map (
            O => \N__54011\,
            I => \N__53718\
        );

    \I__12539\ : InMux
    port map (
            O => \N__54010\,
            I => \N__53718\
        );

    \I__12538\ : CascadeMux
    port map (
            O => \N__54009\,
            I => \N__53710\
        );

    \I__12537\ : CascadeMux
    port map (
            O => \N__54008\,
            I => \N__53704\
        );

    \I__12536\ : CascadeMux
    port map (
            O => \N__54007\,
            I => \N__53701\
        );

    \I__12535\ : CascadeMux
    port map (
            O => \N__54006\,
            I => \N__53698\
        );

    \I__12534\ : CascadeMux
    port map (
            O => \N__54005\,
            I => \N__53695\
        );

    \I__12533\ : CascadeMux
    port map (
            O => \N__54004\,
            I => \N__53691\
        );

    \I__12532\ : CascadeMux
    port map (
            O => \N__54003\,
            I => \N__53688\
        );

    \I__12531\ : CascadeMux
    port map (
            O => \N__54002\,
            I => \N__53685\
        );

    \I__12530\ : CascadeMux
    port map (
            O => \N__54001\,
            I => \N__53682\
        );

    \I__12529\ : CascadeMux
    port map (
            O => \N__54000\,
            I => \N__53679\
        );

    \I__12528\ : CascadeMux
    port map (
            O => \N__53999\,
            I => \N__53676\
        );

    \I__12527\ : CascadeMux
    port map (
            O => \N__53998\,
            I => \N__53673\
        );

    \I__12526\ : CascadeMux
    port map (
            O => \N__53997\,
            I => \N__53670\
        );

    \I__12525\ : CascadeMux
    port map (
            O => \N__53996\,
            I => \N__53667\
        );

    \I__12524\ : CascadeMux
    port map (
            O => \N__53995\,
            I => \N__53664\
        );

    \I__12523\ : CascadeMux
    port map (
            O => \N__53994\,
            I => \N__53661\
        );

    \I__12522\ : CascadeMux
    port map (
            O => \N__53993\,
            I => \N__53658\
        );

    \I__12521\ : CascadeMux
    port map (
            O => \N__53992\,
            I => \N__53655\
        );

    \I__12520\ : CascadeMux
    port map (
            O => \N__53991\,
            I => \N__53652\
        );

    \I__12519\ : CascadeMux
    port map (
            O => \N__53990\,
            I => \N__53649\
        );

    \I__12518\ : CascadeMux
    port map (
            O => \N__53989\,
            I => \N__53646\
        );

    \I__12517\ : CascadeMux
    port map (
            O => \N__53988\,
            I => \N__53643\
        );

    \I__12516\ : CascadeMux
    port map (
            O => \N__53987\,
            I => \N__53640\
        );

    \I__12515\ : CascadeMux
    port map (
            O => \N__53986\,
            I => \N__53633\
        );

    \I__12514\ : CascadeMux
    port map (
            O => \N__53985\,
            I => \N__53630\
        );

    \I__12513\ : CascadeMux
    port map (
            O => \N__53984\,
            I => \N__53627\
        );

    \I__12512\ : CascadeMux
    port map (
            O => \N__53983\,
            I => \N__53624\
        );

    \I__12511\ : CascadeMux
    port map (
            O => \N__53982\,
            I => \N__53621\
        );

    \I__12510\ : CascadeMux
    port map (
            O => \N__53981\,
            I => \N__53617\
        );

    \I__12509\ : Span4Mux_h
    port map (
            O => \N__53968\,
            I => \N__53596\
        );

    \I__12508\ : Span4Mux_v
    port map (
            O => \N__53963\,
            I => \N__53596\
        );

    \I__12507\ : Span4Mux_v
    port map (
            O => \N__53958\,
            I => \N__53596\
        );

    \I__12506\ : LocalMux
    port map (
            O => \N__53955\,
            I => \N__53596\
        );

    \I__12505\ : LocalMux
    port map (
            O => \N__53948\,
            I => \N__53596\
        );

    \I__12504\ : LocalMux
    port map (
            O => \N__53943\,
            I => \N__53593\
        );

    \I__12503\ : LocalMux
    port map (
            O => \N__53938\,
            I => \N__53590\
        );

    \I__12502\ : InMux
    port map (
            O => \N__53937\,
            I => \N__53587\
        );

    \I__12501\ : CascadeMux
    port map (
            O => \N__53936\,
            I => \N__53580\
        );

    \I__12500\ : CascadeMux
    port map (
            O => \N__53935\,
            I => \N__53573\
        );

    \I__12499\ : CascadeMux
    port map (
            O => \N__53934\,
            I => \N__53568\
        );

    \I__12498\ : CascadeMux
    port map (
            O => \N__53933\,
            I => \N__53565\
        );

    \I__12497\ : InMux
    port map (
            O => \N__53930\,
            I => \N__53547\
        );

    \I__12496\ : InMux
    port map (
            O => \N__53927\,
            I => \N__53547\
        );

    \I__12495\ : InMux
    port map (
            O => \N__53926\,
            I => \N__53547\
        );

    \I__12494\ : InMux
    port map (
            O => \N__53925\,
            I => \N__53547\
        );

    \I__12493\ : InMux
    port map (
            O => \N__53922\,
            I => \N__53547\
        );

    \I__12492\ : CascadeMux
    port map (
            O => \N__53921\,
            I => \N__53543\
        );

    \I__12491\ : InMux
    port map (
            O => \N__53918\,
            I => \N__53536\
        );

    \I__12490\ : InMux
    port map (
            O => \N__53917\,
            I => \N__53536\
        );

    \I__12489\ : InMux
    port map (
            O => \N__53916\,
            I => \N__53536\
        );

    \I__12488\ : InMux
    port map (
            O => \N__53915\,
            I => \N__53531\
        );

    \I__12487\ : InMux
    port map (
            O => \N__53912\,
            I => \N__53531\
        );

    \I__12486\ : InMux
    port map (
            O => \N__53909\,
            I => \N__53526\
        );

    \I__12485\ : InMux
    port map (
            O => \N__53906\,
            I => \N__53526\
        );

    \I__12484\ : InMux
    port map (
            O => \N__53905\,
            I => \N__53523\
        );

    \I__12483\ : InMux
    port map (
            O => \N__53904\,
            I => \N__53516\
        );

    \I__12482\ : InMux
    port map (
            O => \N__53903\,
            I => \N__53516\
        );

    \I__12481\ : InMux
    port map (
            O => \N__53902\,
            I => \N__53516\
        );

    \I__12480\ : InMux
    port map (
            O => \N__53899\,
            I => \N__53507\
        );

    \I__12479\ : InMux
    port map (
            O => \N__53898\,
            I => \N__53507\
        );

    \I__12478\ : InMux
    port map (
            O => \N__53897\,
            I => \N__53507\
        );

    \I__12477\ : InMux
    port map (
            O => \N__53896\,
            I => \N__53507\
        );

    \I__12476\ : InMux
    port map (
            O => \N__53893\,
            I => \N__53498\
        );

    \I__12475\ : InMux
    port map (
            O => \N__53892\,
            I => \N__53498\
        );

    \I__12474\ : InMux
    port map (
            O => \N__53891\,
            I => \N__53498\
        );

    \I__12473\ : InMux
    port map (
            O => \N__53890\,
            I => \N__53498\
        );

    \I__12472\ : CascadeMux
    port map (
            O => \N__53889\,
            I => \N__53495\
        );

    \I__12471\ : CascadeMux
    port map (
            O => \N__53888\,
            I => \N__53492\
        );

    \I__12470\ : InMux
    port map (
            O => \N__53885\,
            I => \N__53484\
        );

    \I__12469\ : InMux
    port map (
            O => \N__53882\,
            I => \N__53484\
        );

    \I__12468\ : InMux
    port map (
            O => \N__53879\,
            I => \N__53484\
        );

    \I__12467\ : Span4Mux_h
    port map (
            O => \N__53872\,
            I => \N__53471\
        );

    \I__12466\ : Span4Mux_h
    port map (
            O => \N__53867\,
            I => \N__53471\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__53860\,
            I => \N__53471\
        );

    \I__12464\ : LocalMux
    port map (
            O => \N__53853\,
            I => \N__53471\
        );

    \I__12463\ : LocalMux
    port map (
            O => \N__53846\,
            I => \N__53471\
        );

    \I__12462\ : LocalMux
    port map (
            O => \N__53835\,
            I => \N__53471\
        );

    \I__12461\ : LocalMux
    port map (
            O => \N__53828\,
            I => \N__53468\
        );

    \I__12460\ : InMux
    port map (
            O => \N__53825\,
            I => \N__53457\
        );

    \I__12459\ : InMux
    port map (
            O => \N__53822\,
            I => \N__53457\
        );

    \I__12458\ : InMux
    port map (
            O => \N__53819\,
            I => \N__53457\
        );

    \I__12457\ : InMux
    port map (
            O => \N__53818\,
            I => \N__53457\
        );

    \I__12456\ : InMux
    port map (
            O => \N__53815\,
            I => \N__53457\
        );

    \I__12455\ : InMux
    port map (
            O => \N__53814\,
            I => \N__53454\
        );

    \I__12454\ : CascadeMux
    port map (
            O => \N__53813\,
            I => \N__53446\
        );

    \I__12453\ : CascadeMux
    port map (
            O => \N__53812\,
            I => \N__53442\
        );

    \I__12452\ : CascadeMux
    port map (
            O => \N__53811\,
            I => \N__53429\
        );

    \I__12451\ : CascadeMux
    port map (
            O => \N__53810\,
            I => \N__53426\
        );

    \I__12450\ : CascadeMux
    port map (
            O => \N__53809\,
            I => \N__53422\
        );

    \I__12449\ : CascadeMux
    port map (
            O => \N__53808\,
            I => \N__53419\
        );

    \I__12448\ : CascadeMux
    port map (
            O => \N__53807\,
            I => \N__53414\
        );

    \I__12447\ : LocalMux
    port map (
            O => \N__53802\,
            I => \N__53406\
        );

    \I__12446\ : LocalMux
    port map (
            O => \N__53797\,
            I => \N__53406\
        );

    \I__12445\ : InMux
    port map (
            O => \N__53794\,
            I => \N__53399\
        );

    \I__12444\ : InMux
    port map (
            O => \N__53793\,
            I => \N__53399\
        );

    \I__12443\ : InMux
    port map (
            O => \N__53792\,
            I => \N__53399\
        );

    \I__12442\ : InMux
    port map (
            O => \N__53789\,
            I => \N__53388\
        );

    \I__12441\ : InMux
    port map (
            O => \N__53786\,
            I => \N__53388\
        );

    \I__12440\ : InMux
    port map (
            O => \N__53785\,
            I => \N__53388\
        );

    \I__12439\ : InMux
    port map (
            O => \N__53784\,
            I => \N__53388\
        );

    \I__12438\ : InMux
    port map (
            O => \N__53783\,
            I => \N__53388\
        );

    \I__12437\ : LocalMux
    port map (
            O => \N__53776\,
            I => \N__53380\
        );

    \I__12436\ : LocalMux
    port map (
            O => \N__53769\,
            I => \N__53380\
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__53766\,
            I => \N__53377\
        );

    \I__12434\ : InMux
    port map (
            O => \N__53765\,
            I => \N__53370\
        );

    \I__12433\ : InMux
    port map (
            O => \N__53764\,
            I => \N__53370\
        );

    \I__12432\ : InMux
    port map (
            O => \N__53763\,
            I => \N__53370\
        );

    \I__12431\ : LocalMux
    port map (
            O => \N__53758\,
            I => \N__53359\
        );

    \I__12430\ : LocalMux
    port map (
            O => \N__53747\,
            I => \N__53359\
        );

    \I__12429\ : LocalMux
    port map (
            O => \N__53738\,
            I => \N__53359\
        );

    \I__12428\ : LocalMux
    port map (
            O => \N__53729\,
            I => \N__53359\
        );

    \I__12427\ : LocalMux
    port map (
            O => \N__53718\,
            I => \N__53359\
        );

    \I__12426\ : InMux
    port map (
            O => \N__53717\,
            I => \N__53356\
        );

    \I__12425\ : InMux
    port map (
            O => \N__53716\,
            I => \N__53349\
        );

    \I__12424\ : InMux
    port map (
            O => \N__53715\,
            I => \N__53349\
        );

    \I__12423\ : InMux
    port map (
            O => \N__53714\,
            I => \N__53349\
        );

    \I__12422\ : InMux
    port map (
            O => \N__53713\,
            I => \N__53340\
        );

    \I__12421\ : InMux
    port map (
            O => \N__53710\,
            I => \N__53340\
        );

    \I__12420\ : InMux
    port map (
            O => \N__53709\,
            I => \N__53340\
        );

    \I__12419\ : InMux
    port map (
            O => \N__53708\,
            I => \N__53340\
        );

    \I__12418\ : InMux
    port map (
            O => \N__53707\,
            I => \N__53330\
        );

    \I__12417\ : InMux
    port map (
            O => \N__53704\,
            I => \N__53330\
        );

    \I__12416\ : InMux
    port map (
            O => \N__53701\,
            I => \N__53330\
        );

    \I__12415\ : InMux
    port map (
            O => \N__53698\,
            I => \N__53330\
        );

    \I__12414\ : InMux
    port map (
            O => \N__53695\,
            I => \N__53319\
        );

    \I__12413\ : InMux
    port map (
            O => \N__53694\,
            I => \N__53319\
        );

    \I__12412\ : InMux
    port map (
            O => \N__53691\,
            I => \N__53319\
        );

    \I__12411\ : InMux
    port map (
            O => \N__53688\,
            I => \N__53319\
        );

    \I__12410\ : InMux
    port map (
            O => \N__53685\,
            I => \N__53319\
        );

    \I__12409\ : InMux
    port map (
            O => \N__53682\,
            I => \N__53310\
        );

    \I__12408\ : InMux
    port map (
            O => \N__53679\,
            I => \N__53310\
        );

    \I__12407\ : InMux
    port map (
            O => \N__53676\,
            I => \N__53310\
        );

    \I__12406\ : InMux
    port map (
            O => \N__53673\,
            I => \N__53310\
        );

    \I__12405\ : InMux
    port map (
            O => \N__53670\,
            I => \N__53301\
        );

    \I__12404\ : InMux
    port map (
            O => \N__53667\,
            I => \N__53301\
        );

    \I__12403\ : InMux
    port map (
            O => \N__53664\,
            I => \N__53301\
        );

    \I__12402\ : InMux
    port map (
            O => \N__53661\,
            I => \N__53301\
        );

    \I__12401\ : InMux
    port map (
            O => \N__53658\,
            I => \N__53292\
        );

    \I__12400\ : InMux
    port map (
            O => \N__53655\,
            I => \N__53292\
        );

    \I__12399\ : InMux
    port map (
            O => \N__53652\,
            I => \N__53292\
        );

    \I__12398\ : InMux
    port map (
            O => \N__53649\,
            I => \N__53292\
        );

    \I__12397\ : InMux
    port map (
            O => \N__53646\,
            I => \N__53285\
        );

    \I__12396\ : InMux
    port map (
            O => \N__53643\,
            I => \N__53285\
        );

    \I__12395\ : InMux
    port map (
            O => \N__53640\,
            I => \N__53285\
        );

    \I__12394\ : CascadeMux
    port map (
            O => \N__53639\,
            I => \N__53282\
        );

    \I__12393\ : CascadeMux
    port map (
            O => \N__53638\,
            I => \N__53279\
        );

    \I__12392\ : CascadeMux
    port map (
            O => \N__53637\,
            I => \N__53276\
        );

    \I__12391\ : CascadeMux
    port map (
            O => \N__53636\,
            I => \N__53273\
        );

    \I__12390\ : InMux
    port map (
            O => \N__53633\,
            I => \N__53268\
        );

    \I__12389\ : InMux
    port map (
            O => \N__53630\,
            I => \N__53268\
        );

    \I__12388\ : InMux
    port map (
            O => \N__53627\,
            I => \N__53255\
        );

    \I__12387\ : InMux
    port map (
            O => \N__53624\,
            I => \N__53255\
        );

    \I__12386\ : InMux
    port map (
            O => \N__53621\,
            I => \N__53255\
        );

    \I__12385\ : InMux
    port map (
            O => \N__53620\,
            I => \N__53255\
        );

    \I__12384\ : InMux
    port map (
            O => \N__53617\,
            I => \N__53255\
        );

    \I__12383\ : InMux
    port map (
            O => \N__53616\,
            I => \N__53255\
        );

    \I__12382\ : InMux
    port map (
            O => \N__53615\,
            I => \N__53248\
        );

    \I__12381\ : InMux
    port map (
            O => \N__53614\,
            I => \N__53241\
        );

    \I__12380\ : InMux
    port map (
            O => \N__53613\,
            I => \N__53241\
        );

    \I__12379\ : InMux
    port map (
            O => \N__53612\,
            I => \N__53241\
        );

    \I__12378\ : InMux
    port map (
            O => \N__53611\,
            I => \N__53234\
        );

    \I__12377\ : InMux
    port map (
            O => \N__53610\,
            I => \N__53234\
        );

    \I__12376\ : InMux
    port map (
            O => \N__53609\,
            I => \N__53234\
        );

    \I__12375\ : InMux
    port map (
            O => \N__53608\,
            I => \N__53229\
        );

    \I__12374\ : InMux
    port map (
            O => \N__53607\,
            I => \N__53229\
        );

    \I__12373\ : Span4Mux_h
    port map (
            O => \N__53596\,
            I => \N__53220\
        );

    \I__12372\ : Span4Mux_v
    port map (
            O => \N__53593\,
            I => \N__53220\
        );

    \I__12371\ : Span4Mux_v
    port map (
            O => \N__53590\,
            I => \N__53220\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__53587\,
            I => \N__53220\
        );

    \I__12369\ : InMux
    port map (
            O => \N__53586\,
            I => \N__53213\
        );

    \I__12368\ : InMux
    port map (
            O => \N__53585\,
            I => \N__53213\
        );

    \I__12367\ : InMux
    port map (
            O => \N__53584\,
            I => \N__53213\
        );

    \I__12366\ : InMux
    port map (
            O => \N__53583\,
            I => \N__53202\
        );

    \I__12365\ : InMux
    port map (
            O => \N__53580\,
            I => \N__53202\
        );

    \I__12364\ : InMux
    port map (
            O => \N__53579\,
            I => \N__53202\
        );

    \I__12363\ : InMux
    port map (
            O => \N__53578\,
            I => \N__53202\
        );

    \I__12362\ : InMux
    port map (
            O => \N__53577\,
            I => \N__53202\
        );

    \I__12361\ : CascadeMux
    port map (
            O => \N__53576\,
            I => \N__53199\
        );

    \I__12360\ : InMux
    port map (
            O => \N__53573\,
            I => \N__53180\
        );

    \I__12359\ : InMux
    port map (
            O => \N__53572\,
            I => \N__53180\
        );

    \I__12358\ : InMux
    port map (
            O => \N__53571\,
            I => \N__53180\
        );

    \I__12357\ : InMux
    port map (
            O => \N__53568\,
            I => \N__53169\
        );

    \I__12356\ : InMux
    port map (
            O => \N__53565\,
            I => \N__53169\
        );

    \I__12355\ : InMux
    port map (
            O => \N__53564\,
            I => \N__53169\
        );

    \I__12354\ : InMux
    port map (
            O => \N__53563\,
            I => \N__53169\
        );

    \I__12353\ : InMux
    port map (
            O => \N__53562\,
            I => \N__53169\
        );

    \I__12352\ : InMux
    port map (
            O => \N__53561\,
            I => \N__53164\
        );

    \I__12351\ : InMux
    port map (
            O => \N__53560\,
            I => \N__53164\
        );

    \I__12350\ : CascadeMux
    port map (
            O => \N__53559\,
            I => \N__53161\
        );

    \I__12349\ : CascadeMux
    port map (
            O => \N__53558\,
            I => \N__53155\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__53547\,
            I => \N__53149\
        );

    \I__12347\ : InMux
    port map (
            O => \N__53546\,
            I => \N__53144\
        );

    \I__12346\ : InMux
    port map (
            O => \N__53543\,
            I => \N__53144\
        );

    \I__12345\ : LocalMux
    port map (
            O => \N__53536\,
            I => \N__53141\
        );

    \I__12344\ : LocalMux
    port map (
            O => \N__53531\,
            I => \N__53128\
        );

    \I__12343\ : LocalMux
    port map (
            O => \N__53526\,
            I => \N__53128\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__53523\,
            I => \N__53128\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__53516\,
            I => \N__53128\
        );

    \I__12340\ : LocalMux
    port map (
            O => \N__53507\,
            I => \N__53128\
        );

    \I__12339\ : LocalMux
    port map (
            O => \N__53498\,
            I => \N__53128\
        );

    \I__12338\ : InMux
    port map (
            O => \N__53495\,
            I => \N__53121\
        );

    \I__12337\ : InMux
    port map (
            O => \N__53492\,
            I => \N__53121\
        );

    \I__12336\ : InMux
    port map (
            O => \N__53491\,
            I => \N__53121\
        );

    \I__12335\ : LocalMux
    port map (
            O => \N__53484\,
            I => \N__53116\
        );

    \I__12334\ : Span4Mux_v
    port map (
            O => \N__53471\,
            I => \N__53116\
        );

    \I__12333\ : Span4Mux_v
    port map (
            O => \N__53468\,
            I => \N__53109\
        );

    \I__12332\ : LocalMux
    port map (
            O => \N__53457\,
            I => \N__53109\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__53454\,
            I => \N__53109\
        );

    \I__12330\ : InMux
    port map (
            O => \N__53453\,
            I => \N__53104\
        );

    \I__12329\ : InMux
    port map (
            O => \N__53452\,
            I => \N__53104\
        );

    \I__12328\ : CascadeMux
    port map (
            O => \N__53451\,
            I => \N__53096\
        );

    \I__12327\ : CascadeMux
    port map (
            O => \N__53450\,
            I => \N__53092\
        );

    \I__12326\ : CascadeMux
    port map (
            O => \N__53449\,
            I => \N__53087\
        );

    \I__12325\ : InMux
    port map (
            O => \N__53446\,
            I => \N__53082\
        );

    \I__12324\ : InMux
    port map (
            O => \N__53445\,
            I => \N__53075\
        );

    \I__12323\ : InMux
    port map (
            O => \N__53442\,
            I => \N__53075\
        );

    \I__12322\ : InMux
    port map (
            O => \N__53441\,
            I => \N__53075\
        );

    \I__12321\ : InMux
    port map (
            O => \N__53440\,
            I => \N__53066\
        );

    \I__12320\ : InMux
    port map (
            O => \N__53439\,
            I => \N__53066\
        );

    \I__12319\ : InMux
    port map (
            O => \N__53438\,
            I => \N__53066\
        );

    \I__12318\ : InMux
    port map (
            O => \N__53437\,
            I => \N__53066\
        );

    \I__12317\ : InMux
    port map (
            O => \N__53436\,
            I => \N__53057\
        );

    \I__12316\ : InMux
    port map (
            O => \N__53435\,
            I => \N__53057\
        );

    \I__12315\ : InMux
    port map (
            O => \N__53434\,
            I => \N__53057\
        );

    \I__12314\ : InMux
    port map (
            O => \N__53433\,
            I => \N__53057\
        );

    \I__12313\ : InMux
    port map (
            O => \N__53432\,
            I => \N__53048\
        );

    \I__12312\ : InMux
    port map (
            O => \N__53429\,
            I => \N__53048\
        );

    \I__12311\ : InMux
    port map (
            O => \N__53426\,
            I => \N__53048\
        );

    \I__12310\ : InMux
    port map (
            O => \N__53425\,
            I => \N__53048\
        );

    \I__12309\ : InMux
    port map (
            O => \N__53422\,
            I => \N__53041\
        );

    \I__12308\ : InMux
    port map (
            O => \N__53419\,
            I => \N__53041\
        );

    \I__12307\ : InMux
    port map (
            O => \N__53418\,
            I => \N__53041\
        );

    \I__12306\ : InMux
    port map (
            O => \N__53417\,
            I => \N__53032\
        );

    \I__12305\ : InMux
    port map (
            O => \N__53414\,
            I => \N__53032\
        );

    \I__12304\ : InMux
    port map (
            O => \N__53413\,
            I => \N__53032\
        );

    \I__12303\ : InMux
    port map (
            O => \N__53412\,
            I => \N__53032\
        );

    \I__12302\ : CascadeMux
    port map (
            O => \N__53411\,
            I => \N__53025\
        );

    \I__12301\ : Span4Mux_s2_v
    port map (
            O => \N__53406\,
            I => \N__53022\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__53399\,
            I => \N__53017\
        );

    \I__12299\ : LocalMux
    port map (
            O => \N__53388\,
            I => \N__53017\
        );

    \I__12298\ : CascadeMux
    port map (
            O => \N__53387\,
            I => \N__53013\
        );

    \I__12297\ : CascadeMux
    port map (
            O => \N__53386\,
            I => \N__53009\
        );

    \I__12296\ : CascadeMux
    port map (
            O => \N__53385\,
            I => \N__53005\
        );

    \I__12295\ : Span4Mux_s3_v
    port map (
            O => \N__53380\,
            I => \N__52993\
        );

    \I__12294\ : Span4Mux_s2_h
    port map (
            O => \N__53377\,
            I => \N__52993\
        );

    \I__12293\ : LocalMux
    port map (
            O => \N__53370\,
            I => \N__52993\
        );

    \I__12292\ : Span4Mux_s3_v
    port map (
            O => \N__53359\,
            I => \N__52986\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__53356\,
            I => \N__52986\
        );

    \I__12290\ : LocalMux
    port map (
            O => \N__53349\,
            I => \N__52986\
        );

    \I__12289\ : LocalMux
    port map (
            O => \N__53340\,
            I => \N__52983\
        );

    \I__12288\ : CascadeMux
    port map (
            O => \N__53339\,
            I => \N__52976\
        );

    \I__12287\ : LocalMux
    port map (
            O => \N__53330\,
            I => \N__52966\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__53319\,
            I => \N__52966\
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__53310\,
            I => \N__52957\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__53301\,
            I => \N__52957\
        );

    \I__12283\ : LocalMux
    port map (
            O => \N__53292\,
            I => \N__52957\
        );

    \I__12282\ : LocalMux
    port map (
            O => \N__53285\,
            I => \N__52957\
        );

    \I__12281\ : InMux
    port map (
            O => \N__53282\,
            I => \N__52954\
        );

    \I__12280\ : InMux
    port map (
            O => \N__53279\,
            I => \N__52947\
        );

    \I__12279\ : InMux
    port map (
            O => \N__53276\,
            I => \N__52947\
        );

    \I__12278\ : InMux
    port map (
            O => \N__53273\,
            I => \N__52947\
        );

    \I__12277\ : LocalMux
    port map (
            O => \N__53268\,
            I => \N__52942\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__53255\,
            I => \N__52942\
        );

    \I__12275\ : InMux
    port map (
            O => \N__53254\,
            I => \N__52939\
        );

    \I__12274\ : InMux
    port map (
            O => \N__53253\,
            I => \N__52932\
        );

    \I__12273\ : InMux
    port map (
            O => \N__53252\,
            I => \N__52932\
        );

    \I__12272\ : InMux
    port map (
            O => \N__53251\,
            I => \N__52932\
        );

    \I__12271\ : LocalMux
    port map (
            O => \N__53248\,
            I => \N__52927\
        );

    \I__12270\ : LocalMux
    port map (
            O => \N__53241\,
            I => \N__52927\
        );

    \I__12269\ : LocalMux
    port map (
            O => \N__53234\,
            I => \N__52922\
        );

    \I__12268\ : LocalMux
    port map (
            O => \N__53229\,
            I => \N__52922\
        );

    \I__12267\ : Span4Mux_h
    port map (
            O => \N__53220\,
            I => \N__52915\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__53213\,
            I => \N__52915\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__53202\,
            I => \N__52915\
        );

    \I__12264\ : InMux
    port map (
            O => \N__53199\,
            I => \N__52910\
        );

    \I__12263\ : InMux
    port map (
            O => \N__53198\,
            I => \N__52910\
        );

    \I__12262\ : InMux
    port map (
            O => \N__53197\,
            I => \N__52905\
        );

    \I__12261\ : InMux
    port map (
            O => \N__53196\,
            I => \N__52905\
        );

    \I__12260\ : CascadeMux
    port map (
            O => \N__53195\,
            I => \N__52887\
        );

    \I__12259\ : CascadeMux
    port map (
            O => \N__53194\,
            I => \N__52883\
        );

    \I__12258\ : CascadeMux
    port map (
            O => \N__53193\,
            I => \N__52880\
        );

    \I__12257\ : CascadeMux
    port map (
            O => \N__53192\,
            I => \N__52877\
        );

    \I__12256\ : CascadeMux
    port map (
            O => \N__53191\,
            I => \N__52874\
        );

    \I__12255\ : CascadeMux
    port map (
            O => \N__53190\,
            I => \N__52871\
        );

    \I__12254\ : CascadeMux
    port map (
            O => \N__53189\,
            I => \N__52868\
        );

    \I__12253\ : CascadeMux
    port map (
            O => \N__53188\,
            I => \N__52865\
        );

    \I__12252\ : CascadeMux
    port map (
            O => \N__53187\,
            I => \N__52862\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__53180\,
            I => \N__52855\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__53169\,
            I => \N__52855\
        );

    \I__12249\ : LocalMux
    port map (
            O => \N__53164\,
            I => \N__52855\
        );

    \I__12248\ : InMux
    port map (
            O => \N__53161\,
            I => \N__52846\
        );

    \I__12247\ : InMux
    port map (
            O => \N__53160\,
            I => \N__52846\
        );

    \I__12246\ : InMux
    port map (
            O => \N__53159\,
            I => \N__52846\
        );

    \I__12245\ : InMux
    port map (
            O => \N__53158\,
            I => \N__52846\
        );

    \I__12244\ : InMux
    port map (
            O => \N__53155\,
            I => \N__52837\
        );

    \I__12243\ : InMux
    port map (
            O => \N__53154\,
            I => \N__52837\
        );

    \I__12242\ : InMux
    port map (
            O => \N__53153\,
            I => \N__52837\
        );

    \I__12241\ : InMux
    port map (
            O => \N__53152\,
            I => \N__52837\
        );

    \I__12240\ : Span4Mux_h
    port map (
            O => \N__53149\,
            I => \N__52832\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__53144\,
            I => \N__52832\
        );

    \I__12238\ : Span4Mux_v
    port map (
            O => \N__53141\,
            I => \N__52821\
        );

    \I__12237\ : Span4Mux_v
    port map (
            O => \N__53128\,
            I => \N__52821\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__53121\,
            I => \N__52821\
        );

    \I__12235\ : Span4Mux_v
    port map (
            O => \N__53116\,
            I => \N__52821\
        );

    \I__12234\ : Span4Mux_v
    port map (
            O => \N__53109\,
            I => \N__52821\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__53104\,
            I => \N__52818\
        );

    \I__12232\ : InMux
    port map (
            O => \N__53103\,
            I => \N__52811\
        );

    \I__12231\ : InMux
    port map (
            O => \N__53102\,
            I => \N__52811\
        );

    \I__12230\ : InMux
    port map (
            O => \N__53101\,
            I => \N__52811\
        );

    \I__12229\ : InMux
    port map (
            O => \N__53100\,
            I => \N__52801\
        );

    \I__12228\ : InMux
    port map (
            O => \N__53099\,
            I => \N__52801\
        );

    \I__12227\ : InMux
    port map (
            O => \N__53096\,
            I => \N__52801\
        );

    \I__12226\ : InMux
    port map (
            O => \N__53095\,
            I => \N__52801\
        );

    \I__12225\ : InMux
    port map (
            O => \N__53092\,
            I => \N__52794\
        );

    \I__12224\ : InMux
    port map (
            O => \N__53091\,
            I => \N__52794\
        );

    \I__12223\ : InMux
    port map (
            O => \N__53090\,
            I => \N__52794\
        );

    \I__12222\ : InMux
    port map (
            O => \N__53087\,
            I => \N__52787\
        );

    \I__12221\ : InMux
    port map (
            O => \N__53086\,
            I => \N__52787\
        );

    \I__12220\ : InMux
    port map (
            O => \N__53085\,
            I => \N__52787\
        );

    \I__12219\ : LocalMux
    port map (
            O => \N__53082\,
            I => \N__52771\
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__53075\,
            I => \N__52771\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__53066\,
            I => \N__52771\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__53057\,
            I => \N__52771\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__53048\,
            I => \N__52771\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__53041\,
            I => \N__52771\
        );

    \I__12213\ : LocalMux
    port map (
            O => \N__53032\,
            I => \N__52771\
        );

    \I__12212\ : InMux
    port map (
            O => \N__53031\,
            I => \N__52768\
        );

    \I__12211\ : InMux
    port map (
            O => \N__53030\,
            I => \N__52761\
        );

    \I__12210\ : InMux
    port map (
            O => \N__53029\,
            I => \N__52761\
        );

    \I__12209\ : InMux
    port map (
            O => \N__53028\,
            I => \N__52761\
        );

    \I__12208\ : InMux
    port map (
            O => \N__53025\,
            I => \N__52758\
        );

    \I__12207\ : Span4Mux_v
    port map (
            O => \N__53022\,
            I => \N__52753\
        );

    \I__12206\ : Span4Mux_v
    port map (
            O => \N__53017\,
            I => \N__52753\
        );

    \I__12205\ : InMux
    port map (
            O => \N__53016\,
            I => \N__52742\
        );

    \I__12204\ : InMux
    port map (
            O => \N__53013\,
            I => \N__52742\
        );

    \I__12203\ : InMux
    port map (
            O => \N__53012\,
            I => \N__52742\
        );

    \I__12202\ : InMux
    port map (
            O => \N__53009\,
            I => \N__52742\
        );

    \I__12201\ : InMux
    port map (
            O => \N__53008\,
            I => \N__52742\
        );

    \I__12200\ : InMux
    port map (
            O => \N__53005\,
            I => \N__52735\
        );

    \I__12199\ : InMux
    port map (
            O => \N__53004\,
            I => \N__52735\
        );

    \I__12198\ : InMux
    port map (
            O => \N__53003\,
            I => \N__52735\
        );

    \I__12197\ : CascadeMux
    port map (
            O => \N__53002\,
            I => \N__52727\
        );

    \I__12196\ : CascadeMux
    port map (
            O => \N__53001\,
            I => \N__52718\
        );

    \I__12195\ : CascadeMux
    port map (
            O => \N__53000\,
            I => \N__52714\
        );

    \I__12194\ : Span4Mux_v
    port map (
            O => \N__52993\,
            I => \N__52704\
        );

    \I__12193\ : Span4Mux_v
    port map (
            O => \N__52986\,
            I => \N__52704\
        );

    \I__12192\ : Span4Mux_v
    port map (
            O => \N__52983\,
            I => \N__52704\
        );

    \I__12191\ : InMux
    port map (
            O => \N__52982\,
            I => \N__52697\
        );

    \I__12190\ : InMux
    port map (
            O => \N__52981\,
            I => \N__52697\
        );

    \I__12189\ : InMux
    port map (
            O => \N__52980\,
            I => \N__52697\
        );

    \I__12188\ : InMux
    port map (
            O => \N__52979\,
            I => \N__52694\
        );

    \I__12187\ : InMux
    port map (
            O => \N__52976\,
            I => \N__52689\
        );

    \I__12186\ : InMux
    port map (
            O => \N__52975\,
            I => \N__52689\
        );

    \I__12185\ : InMux
    port map (
            O => \N__52974\,
            I => \N__52684\
        );

    \I__12184\ : InMux
    port map (
            O => \N__52973\,
            I => \N__52684\
        );

    \I__12183\ : InMux
    port map (
            O => \N__52972\,
            I => \N__52679\
        );

    \I__12182\ : InMux
    port map (
            O => \N__52971\,
            I => \N__52679\
        );

    \I__12181\ : Span4Mux_s3_v
    port map (
            O => \N__52966\,
            I => \N__52672\
        );

    \I__12180\ : Span4Mux_s3_v
    port map (
            O => \N__52957\,
            I => \N__52672\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__52954\,
            I => \N__52672\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__52947\,
            I => \N__52669\
        );

    \I__12177\ : Span4Mux_s3_h
    port map (
            O => \N__52942\,
            I => \N__52662\
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__52939\,
            I => \N__52662\
        );

    \I__12175\ : LocalMux
    port map (
            O => \N__52932\,
            I => \N__52662\
        );

    \I__12174\ : Span4Mux_v
    port map (
            O => \N__52927\,
            I => \N__52651\
        );

    \I__12173\ : Span4Mux_v
    port map (
            O => \N__52922\,
            I => \N__52651\
        );

    \I__12172\ : Span4Mux_v
    port map (
            O => \N__52915\,
            I => \N__52651\
        );

    \I__12171\ : LocalMux
    port map (
            O => \N__52910\,
            I => \N__52651\
        );

    \I__12170\ : LocalMux
    port map (
            O => \N__52905\,
            I => \N__52651\
        );

    \I__12169\ : InMux
    port map (
            O => \N__52904\,
            I => \N__52646\
        );

    \I__12168\ : InMux
    port map (
            O => \N__52903\,
            I => \N__52646\
        );

    \I__12167\ : InMux
    port map (
            O => \N__52902\,
            I => \N__52641\
        );

    \I__12166\ : InMux
    port map (
            O => \N__52901\,
            I => \N__52641\
        );

    \I__12165\ : InMux
    port map (
            O => \N__52900\,
            I => \N__52634\
        );

    \I__12164\ : InMux
    port map (
            O => \N__52899\,
            I => \N__52634\
        );

    \I__12163\ : InMux
    port map (
            O => \N__52898\,
            I => \N__52634\
        );

    \I__12162\ : InMux
    port map (
            O => \N__52897\,
            I => \N__52631\
        );

    \I__12161\ : InMux
    port map (
            O => \N__52896\,
            I => \N__52624\
        );

    \I__12160\ : InMux
    port map (
            O => \N__52895\,
            I => \N__52624\
        );

    \I__12159\ : InMux
    port map (
            O => \N__52894\,
            I => \N__52624\
        );

    \I__12158\ : InMux
    port map (
            O => \N__52893\,
            I => \N__52619\
        );

    \I__12157\ : InMux
    port map (
            O => \N__52892\,
            I => \N__52619\
        );

    \I__12156\ : InMux
    port map (
            O => \N__52891\,
            I => \N__52616\
        );

    \I__12155\ : InMux
    port map (
            O => \N__52890\,
            I => \N__52609\
        );

    \I__12154\ : InMux
    port map (
            O => \N__52887\,
            I => \N__52609\
        );

    \I__12153\ : InMux
    port map (
            O => \N__52886\,
            I => \N__52609\
        );

    \I__12152\ : InMux
    port map (
            O => \N__52883\,
            I => \N__52600\
        );

    \I__12151\ : InMux
    port map (
            O => \N__52880\,
            I => \N__52600\
        );

    \I__12150\ : InMux
    port map (
            O => \N__52877\,
            I => \N__52600\
        );

    \I__12149\ : InMux
    port map (
            O => \N__52874\,
            I => \N__52600\
        );

    \I__12148\ : InMux
    port map (
            O => \N__52871\,
            I => \N__52591\
        );

    \I__12147\ : InMux
    port map (
            O => \N__52868\,
            I => \N__52591\
        );

    \I__12146\ : InMux
    port map (
            O => \N__52865\,
            I => \N__52591\
        );

    \I__12145\ : InMux
    port map (
            O => \N__52862\,
            I => \N__52591\
        );

    \I__12144\ : Span4Mux_h
    port map (
            O => \N__52855\,
            I => \N__52583\
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__52846\,
            I => \N__52583\
        );

    \I__12142\ : LocalMux
    port map (
            O => \N__52837\,
            I => \N__52583\
        );

    \I__12141\ : Span4Mux_h
    port map (
            O => \N__52832\,
            I => \N__52576\
        );

    \I__12140\ : Span4Mux_h
    port map (
            O => \N__52821\,
            I => \N__52576\
        );

    \I__12139\ : Span4Mux_v
    port map (
            O => \N__52818\,
            I => \N__52576\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__52811\,
            I => \N__52573\
        );

    \I__12137\ : InMux
    port map (
            O => \N__52810\,
            I => \N__52570\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__52801\,
            I => \N__52563\
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__52794\,
            I => \N__52563\
        );

    \I__12134\ : LocalMux
    port map (
            O => \N__52787\,
            I => \N__52563\
        );

    \I__12133\ : InMux
    port map (
            O => \N__52786\,
            I => \N__52560\
        );

    \I__12132\ : Span12Mux_v
    port map (
            O => \N__52771\,
            I => \N__52542\
        );

    \I__12131\ : LocalMux
    port map (
            O => \N__52768\,
            I => \N__52542\
        );

    \I__12130\ : LocalMux
    port map (
            O => \N__52761\,
            I => \N__52542\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__52758\,
            I => \N__52542\
        );

    \I__12128\ : Sp12to4
    port map (
            O => \N__52753\,
            I => \N__52542\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__52742\,
            I => \N__52542\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__52735\,
            I => \N__52542\
        );

    \I__12125\ : InMux
    port map (
            O => \N__52734\,
            I => \N__52539\
        );

    \I__12124\ : InMux
    port map (
            O => \N__52733\,
            I => \N__52532\
        );

    \I__12123\ : InMux
    port map (
            O => \N__52732\,
            I => \N__52532\
        );

    \I__12122\ : InMux
    port map (
            O => \N__52731\,
            I => \N__52532\
        );

    \I__12121\ : InMux
    port map (
            O => \N__52730\,
            I => \N__52521\
        );

    \I__12120\ : InMux
    port map (
            O => \N__52727\,
            I => \N__52521\
        );

    \I__12119\ : InMux
    port map (
            O => \N__52726\,
            I => \N__52521\
        );

    \I__12118\ : InMux
    port map (
            O => \N__52725\,
            I => \N__52521\
        );

    \I__12117\ : InMux
    port map (
            O => \N__52724\,
            I => \N__52521\
        );

    \I__12116\ : InMux
    port map (
            O => \N__52723\,
            I => \N__52514\
        );

    \I__12115\ : InMux
    port map (
            O => \N__52722\,
            I => \N__52514\
        );

    \I__12114\ : InMux
    port map (
            O => \N__52721\,
            I => \N__52514\
        );

    \I__12113\ : InMux
    port map (
            O => \N__52718\,
            I => \N__52505\
        );

    \I__12112\ : InMux
    port map (
            O => \N__52717\,
            I => \N__52505\
        );

    \I__12111\ : InMux
    port map (
            O => \N__52714\,
            I => \N__52505\
        );

    \I__12110\ : InMux
    port map (
            O => \N__52713\,
            I => \N__52505\
        );

    \I__12109\ : InMux
    port map (
            O => \N__52712\,
            I => \N__52500\
        );

    \I__12108\ : InMux
    port map (
            O => \N__52711\,
            I => \N__52500\
        );

    \I__12107\ : Span4Mux_h
    port map (
            O => \N__52704\,
            I => \N__52497\
        );

    \I__12106\ : LocalMux
    port map (
            O => \N__52697\,
            I => \N__52494\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__52694\,
            I => \N__52485\
        );

    \I__12104\ : LocalMux
    port map (
            O => \N__52689\,
            I => \N__52485\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__52684\,
            I => \N__52485\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__52679\,
            I => \N__52485\
        );

    \I__12101\ : Span4Mux_v
    port map (
            O => \N__52672\,
            I => \N__52478\
        );

    \I__12100\ : Span4Mux_v
    port map (
            O => \N__52669\,
            I => \N__52478\
        );

    \I__12099\ : Span4Mux_h
    port map (
            O => \N__52662\,
            I => \N__52478\
        );

    \I__12098\ : Span4Mux_h
    port map (
            O => \N__52651\,
            I => \N__52471\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__52646\,
            I => \N__52471\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__52641\,
            I => \N__52471\
        );

    \I__12095\ : LocalMux
    port map (
            O => \N__52634\,
            I => \N__52460\
        );

    \I__12094\ : LocalMux
    port map (
            O => \N__52631\,
            I => \N__52460\
        );

    \I__12093\ : LocalMux
    port map (
            O => \N__52624\,
            I => \N__52460\
        );

    \I__12092\ : LocalMux
    port map (
            O => \N__52619\,
            I => \N__52460\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__52616\,
            I => \N__52460\
        );

    \I__12090\ : LocalMux
    port map (
            O => \N__52609\,
            I => \N__52453\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__52600\,
            I => \N__52453\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__52591\,
            I => \N__52453\
        );

    \I__12087\ : InMux
    port map (
            O => \N__52590\,
            I => \N__52450\
        );

    \I__12086\ : Span4Mux_h
    port map (
            O => \N__52583\,
            I => \N__52437\
        );

    \I__12085\ : Span4Mux_h
    port map (
            O => \N__52576\,
            I => \N__52437\
        );

    \I__12084\ : Span4Mux_v
    port map (
            O => \N__52573\,
            I => \N__52437\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__52570\,
            I => \N__52437\
        );

    \I__12082\ : Span4Mux_h
    port map (
            O => \N__52563\,
            I => \N__52437\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__52560\,
            I => \N__52437\
        );

    \I__12080\ : InMux
    port map (
            O => \N__52559\,
            I => \N__52430\
        );

    \I__12079\ : InMux
    port map (
            O => \N__52558\,
            I => \N__52430\
        );

    \I__12078\ : InMux
    port map (
            O => \N__52557\,
            I => \N__52430\
        );

    \I__12077\ : Span12Mux_h
    port map (
            O => \N__52542\,
            I => \N__52412\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__52539\,
            I => \N__52412\
        );

    \I__12075\ : LocalMux
    port map (
            O => \N__52532\,
            I => \N__52412\
        );

    \I__12074\ : LocalMux
    port map (
            O => \N__52521\,
            I => \N__52412\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__52514\,
            I => \N__52412\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__52505\,
            I => \N__52412\
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__52500\,
            I => \N__52412\
        );

    \I__12070\ : Span4Mux_h
    port map (
            O => \N__52497\,
            I => \N__52405\
        );

    \I__12069\ : Span4Mux_v
    port map (
            O => \N__52494\,
            I => \N__52405\
        );

    \I__12068\ : Span4Mux_v
    port map (
            O => \N__52485\,
            I => \N__52405\
        );

    \I__12067\ : Span4Mux_h
    port map (
            O => \N__52478\,
            I => \N__52398\
        );

    \I__12066\ : Span4Mux_v
    port map (
            O => \N__52471\,
            I => \N__52398\
        );

    \I__12065\ : Span4Mux_v
    port map (
            O => \N__52460\,
            I => \N__52398\
        );

    \I__12064\ : Span12Mux_h
    port map (
            O => \N__52453\,
            I => \N__52393\
        );

    \I__12063\ : LocalMux
    port map (
            O => \N__52450\,
            I => \N__52393\
        );

    \I__12062\ : Span4Mux_v
    port map (
            O => \N__52437\,
            I => \N__52388\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__52430\,
            I => \N__52388\
        );

    \I__12060\ : InMux
    port map (
            O => \N__52429\,
            I => \N__52385\
        );

    \I__12059\ : InMux
    port map (
            O => \N__52428\,
            I => \N__52380\
        );

    \I__12058\ : InMux
    port map (
            O => \N__52427\,
            I => \N__52380\
        );

    \I__12057\ : Odrv12
    port map (
            O => \N__52412\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12056\ : Odrv4
    port map (
            O => \N__52405\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12055\ : Odrv4
    port map (
            O => \N__52398\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12054\ : Odrv12
    port map (
            O => \N__52393\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12053\ : Odrv4
    port map (
            O => \N__52388\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12052\ : LocalMux
    port map (
            O => \N__52385\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12051\ : LocalMux
    port map (
            O => \N__52380\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12050\ : InMux
    port map (
            O => \N__52365\,
            I => \N__52362\
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__52362\,
            I => \N__52359\
        );

    \I__12048\ : Span4Mux_v
    port map (
            O => \N__52359\,
            I => \N__52356\
        );

    \I__12047\ : Sp12to4
    port map (
            O => \N__52356\,
            I => \N__52352\
        );

    \I__12046\ : InMux
    port map (
            O => \N__52355\,
            I => \N__52349\
        );

    \I__12045\ : Odrv12
    port map (
            O => \N__52352\,
            I => n15513
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__52349\,
            I => n15513
        );

    \I__12043\ : CascadeMux
    port map (
            O => \N__52344\,
            I => \N__52341\
        );

    \I__12042\ : InMux
    port map (
            O => \N__52341\,
            I => \N__52338\
        );

    \I__12041\ : LocalMux
    port map (
            O => \N__52338\,
            I => \N__52334\
        );

    \I__12040\ : InMux
    port map (
            O => \N__52337\,
            I => \N__52331\
        );

    \I__12039\ : Odrv4
    port map (
            O => \N__52334\,
            I => n1125
        );

    \I__12038\ : LocalMux
    port map (
            O => \N__52331\,
            I => n1125
        );

    \I__12037\ : InMux
    port map (
            O => \N__52326\,
            I => n12516
        );

    \I__12036\ : CascadeMux
    port map (
            O => \N__52323\,
            I => \N__52319\
        );

    \I__12035\ : InMux
    port map (
            O => \N__52322\,
            I => \N__52316\
        );

    \I__12034\ : InMux
    port map (
            O => \N__52319\,
            I => \N__52313\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__52316\,
            I => \N__52310\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__52313\,
            I => n1224
        );

    \I__12031\ : Odrv4
    port map (
            O => \N__52310\,
            I => n1224
        );

    \I__12030\ : CascadeMux
    port map (
            O => \N__52305\,
            I => \N__52301\
        );

    \I__12029\ : InMux
    port map (
            O => \N__52304\,
            I => \N__52296\
        );

    \I__12028\ : InMux
    port map (
            O => \N__52301\,
            I => \N__52296\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__52296\,
            I => \N__52293\
        );

    \I__12026\ : Span4Mux_h
    port map (
            O => \N__52293\,
            I => \N__52290\
        );

    \I__12025\ : Odrv4
    port map (
            O => \N__52290\,
            I => n1126
        );

    \I__12024\ : CascadeMux
    port map (
            O => \N__52287\,
            I => \N__52284\
        );

    \I__12023\ : InMux
    port map (
            O => \N__52284\,
            I => \N__52281\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__52281\,
            I => n1193
        );

    \I__12021\ : CascadeMux
    port map (
            O => \N__52278\,
            I => \N__52271\
        );

    \I__12020\ : CascadeMux
    port map (
            O => \N__52277\,
            I => \N__52268\
        );

    \I__12019\ : CascadeMux
    port map (
            O => \N__52276\,
            I => \N__52265\
        );

    \I__12018\ : InMux
    port map (
            O => \N__52275\,
            I => \N__52261\
        );

    \I__12017\ : InMux
    port map (
            O => \N__52274\,
            I => \N__52258\
        );

    \I__12016\ : InMux
    port map (
            O => \N__52271\,
            I => \N__52249\
        );

    \I__12015\ : InMux
    port map (
            O => \N__52268\,
            I => \N__52249\
        );

    \I__12014\ : InMux
    port map (
            O => \N__52265\,
            I => \N__52249\
        );

    \I__12013\ : InMux
    port map (
            O => \N__52264\,
            I => \N__52249\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__52261\,
            I => \N__52246\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__52258\,
            I => \N__52242\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__52249\,
            I => \N__52236\
        );

    \I__12009\ : Span12Mux_s9_v
    port map (
            O => \N__52246\,
            I => \N__52233\
        );

    \I__12008\ : InMux
    port map (
            O => \N__52245\,
            I => \N__52230\
        );

    \I__12007\ : Span4Mux_h
    port map (
            O => \N__52242\,
            I => \N__52227\
        );

    \I__12006\ : InMux
    port map (
            O => \N__52241\,
            I => \N__52224\
        );

    \I__12005\ : InMux
    port map (
            O => \N__52240\,
            I => \N__52221\
        );

    \I__12004\ : InMux
    port map (
            O => \N__52239\,
            I => \N__52218\
        );

    \I__12003\ : Span4Mux_h
    port map (
            O => \N__52236\,
            I => \N__52215\
        );

    \I__12002\ : Odrv12
    port map (
            O => \N__52233\,
            I => n1158
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__52230\,
            I => n1158
        );

    \I__12000\ : Odrv4
    port map (
            O => \N__52227\,
            I => n1158
        );

    \I__11999\ : LocalMux
    port map (
            O => \N__52224\,
            I => n1158
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__52221\,
            I => n1158
        );

    \I__11997\ : LocalMux
    port map (
            O => \N__52218\,
            I => n1158
        );

    \I__11996\ : Odrv4
    port map (
            O => \N__52215\,
            I => n1158
        );

    \I__11995\ : InMux
    port map (
            O => \N__52200\,
            I => \N__52197\
        );

    \I__11994\ : LocalMux
    port map (
            O => \N__52197\,
            I => \N__52192\
        );

    \I__11993\ : CascadeMux
    port map (
            O => \N__52196\,
            I => \N__52189\
        );

    \I__11992\ : InMux
    port map (
            O => \N__52195\,
            I => \N__52186\
        );

    \I__11991\ : Span4Mux_h
    port map (
            O => \N__52192\,
            I => \N__52183\
        );

    \I__11990\ : InMux
    port map (
            O => \N__52189\,
            I => \N__52180\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__52186\,
            I => \N__52177\
        );

    \I__11988\ : Odrv4
    port map (
            O => \N__52183\,
            I => n1225
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__52180\,
            I => n1225
        );

    \I__11986\ : Odrv12
    port map (
            O => \N__52177\,
            I => n1225
        );

    \I__11985\ : InMux
    port map (
            O => \N__52170\,
            I => \N__52167\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__52167\,
            I => \N__52164\
        );

    \I__11983\ : Odrv12
    port map (
            O => \N__52164\,
            I => n23_adj_700
        );

    \I__11982\ : CascadeMux
    port map (
            O => \N__52161\,
            I => \N__52158\
        );

    \I__11981\ : InMux
    port map (
            O => \N__52158\,
            I => \N__52155\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__52155\,
            I => \N__52152\
        );

    \I__11979\ : Odrv4
    port map (
            O => \N__52152\,
            I => n25_adj_698
        );

    \I__11978\ : CascadeMux
    port map (
            O => \N__52149\,
            I => \direction_N_342_cascade_\
        );

    \I__11977\ : CascadeMux
    port map (
            O => \N__52146\,
            I => \N__52143\
        );

    \I__11976\ : InMux
    port map (
            O => \N__52143\,
            I => \N__52140\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__52140\,
            I => n1693
        );

    \I__11974\ : InMux
    port map (
            O => \N__52137\,
            I => \N__52133\
        );

    \I__11973\ : InMux
    port map (
            O => \N__52136\,
            I => \N__52130\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__52133\,
            I => \N__52125\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__52130\,
            I => \N__52125\
        );

    \I__11970\ : Span4Mux_h
    port map (
            O => \N__52125\,
            I => \N__52122\
        );

    \I__11969\ : Odrv4
    port map (
            O => \N__52122\,
            I => \direction_N_340\
        );

    \I__11968\ : InMux
    port map (
            O => \N__52119\,
            I => \N__52116\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__52116\,
            I => \direction_N_342\
        );

    \I__11966\ : CascadeMux
    port map (
            O => \N__52113\,
            I => \n13661_cascade_\
        );

    \I__11965\ : InMux
    port map (
            O => \N__52110\,
            I => \N__52103\
        );

    \I__11964\ : CascadeMux
    port map (
            O => \N__52109\,
            I => \N__52100\
        );

    \I__11963\ : CascadeMux
    port map (
            O => \N__52108\,
            I => \N__52096\
        );

    \I__11962\ : CascadeMux
    port map (
            O => \N__52107\,
            I => \N__52092\
        );

    \I__11961\ : CascadeMux
    port map (
            O => \N__52106\,
            I => \N__52088\
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__52103\,
            I => \N__52078\
        );

    \I__11959\ : InMux
    port map (
            O => \N__52100\,
            I => \N__52061\
        );

    \I__11958\ : InMux
    port map (
            O => \N__52099\,
            I => \N__52061\
        );

    \I__11957\ : InMux
    port map (
            O => \N__52096\,
            I => \N__52061\
        );

    \I__11956\ : InMux
    port map (
            O => \N__52095\,
            I => \N__52061\
        );

    \I__11955\ : InMux
    port map (
            O => \N__52092\,
            I => \N__52061\
        );

    \I__11954\ : InMux
    port map (
            O => \N__52091\,
            I => \N__52061\
        );

    \I__11953\ : InMux
    port map (
            O => \N__52088\,
            I => \N__52061\
        );

    \I__11952\ : InMux
    port map (
            O => \N__52087\,
            I => \N__52061\
        );

    \I__11951\ : CascadeMux
    port map (
            O => \N__52086\,
            I => \N__52058\
        );

    \I__11950\ : CascadeMux
    port map (
            O => \N__52085\,
            I => \N__52054\
        );

    \I__11949\ : CascadeMux
    port map (
            O => \N__52084\,
            I => \N__52050\
        );

    \I__11948\ : CascadeMux
    port map (
            O => \N__52083\,
            I => \N__52046\
        );

    \I__11947\ : CascadeMux
    port map (
            O => \N__52082\,
            I => \N__52039\
        );

    \I__11946\ : InMux
    port map (
            O => \N__52081\,
            I => \N__52030\
        );

    \I__11945\ : Span4Mux_v
    port map (
            O => \N__52078\,
            I => \N__52025\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__52061\,
            I => \N__52025\
        );

    \I__11943\ : InMux
    port map (
            O => \N__52058\,
            I => \N__52008\
        );

    \I__11942\ : InMux
    port map (
            O => \N__52057\,
            I => \N__52008\
        );

    \I__11941\ : InMux
    port map (
            O => \N__52054\,
            I => \N__52008\
        );

    \I__11940\ : InMux
    port map (
            O => \N__52053\,
            I => \N__52008\
        );

    \I__11939\ : InMux
    port map (
            O => \N__52050\,
            I => \N__52008\
        );

    \I__11938\ : InMux
    port map (
            O => \N__52049\,
            I => \N__52008\
        );

    \I__11937\ : InMux
    port map (
            O => \N__52046\,
            I => \N__52008\
        );

    \I__11936\ : InMux
    port map (
            O => \N__52045\,
            I => \N__52008\
        );

    \I__11935\ : InMux
    port map (
            O => \N__52044\,
            I => \N__51999\
        );

    \I__11934\ : InMux
    port map (
            O => \N__52043\,
            I => \N__51999\
        );

    \I__11933\ : InMux
    port map (
            O => \N__52042\,
            I => \N__51999\
        );

    \I__11932\ : InMux
    port map (
            O => \N__52039\,
            I => \N__51999\
        );

    \I__11931\ : InMux
    port map (
            O => \N__52038\,
            I => \N__51990\
        );

    \I__11930\ : InMux
    port map (
            O => \N__52037\,
            I => \N__51990\
        );

    \I__11929\ : InMux
    port map (
            O => \N__52036\,
            I => \N__51990\
        );

    \I__11928\ : InMux
    port map (
            O => \N__52035\,
            I => \N__51990\
        );

    \I__11927\ : InMux
    port map (
            O => \N__52034\,
            I => \N__51985\
        );

    \I__11926\ : InMux
    port map (
            O => \N__52033\,
            I => \N__51985\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__52030\,
            I => direction_c
        );

    \I__11924\ : Odrv4
    port map (
            O => \N__52025\,
            I => direction_c
        );

    \I__11923\ : LocalMux
    port map (
            O => \N__52008\,
            I => direction_c
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__51999\,
            I => direction_c
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__51990\,
            I => direction_c
        );

    \I__11920\ : LocalMux
    port map (
            O => \N__51985\,
            I => direction_c
        );

    \I__11919\ : CascadeMux
    port map (
            O => \N__51972\,
            I => \n22_adj_705_cascade_\
        );

    \I__11918\ : InMux
    port map (
            O => \N__51969\,
            I => \N__51966\
        );

    \I__11917\ : LocalMux
    port map (
            O => \N__51966\,
            I => \N__51963\
        );

    \I__11916\ : Odrv4
    port map (
            O => \N__51963\,
            I => n1200
        );

    \I__11915\ : InMux
    port map (
            O => \N__51960\,
            I => n12508
        );

    \I__11914\ : InMux
    port map (
            O => \N__51957\,
            I => \N__51954\
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__51954\,
            I => \N__51950\
        );

    \I__11912\ : InMux
    port map (
            O => \N__51953\,
            I => \N__51947\
        );

    \I__11911\ : Span4Mux_v
    port map (
            O => \N__51950\,
            I => \N__51944\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__51947\,
            I => n1132
        );

    \I__11909\ : Odrv4
    port map (
            O => \N__51944\,
            I => n1132
        );

    \I__11908\ : InMux
    port map (
            O => \N__51939\,
            I => \N__51936\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__51936\,
            I => \N__51933\
        );

    \I__11906\ : Span4Mux_h
    port map (
            O => \N__51933\,
            I => \N__51930\
        );

    \I__11905\ : Odrv4
    port map (
            O => \N__51930\,
            I => n1199
        );

    \I__11904\ : InMux
    port map (
            O => \N__51927\,
            I => n12509
        );

    \I__11903\ : CascadeMux
    port map (
            O => \N__51924\,
            I => \N__51921\
        );

    \I__11902\ : InMux
    port map (
            O => \N__51921\,
            I => \N__51917\
        );

    \I__11901\ : InMux
    port map (
            O => \N__51920\,
            I => \N__51914\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__51917\,
            I => \N__51910\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__51914\,
            I => \N__51907\
        );

    \I__11898\ : InMux
    port map (
            O => \N__51913\,
            I => \N__51904\
        );

    \I__11897\ : Span4Mux_h
    port map (
            O => \N__51910\,
            I => \N__51901\
        );

    \I__11896\ : Odrv4
    port map (
            O => \N__51907\,
            I => n1131
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__51904\,
            I => n1131
        );

    \I__11894\ : Odrv4
    port map (
            O => \N__51901\,
            I => n1131
        );

    \I__11893\ : CascadeMux
    port map (
            O => \N__51894\,
            I => \N__51891\
        );

    \I__11892\ : InMux
    port map (
            O => \N__51891\,
            I => \N__51888\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__51888\,
            I => n1198
        );

    \I__11890\ : InMux
    port map (
            O => \N__51885\,
            I => n12510
        );

    \I__11889\ : InMux
    port map (
            O => \N__51882\,
            I => \N__51878\
        );

    \I__11888\ : CascadeMux
    port map (
            O => \N__51881\,
            I => \N__51875\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__51878\,
            I => \N__51871\
        );

    \I__11886\ : InMux
    port map (
            O => \N__51875\,
            I => \N__51868\
        );

    \I__11885\ : CascadeMux
    port map (
            O => \N__51874\,
            I => \N__51865\
        );

    \I__11884\ : Span4Mux_v
    port map (
            O => \N__51871\,
            I => \N__51860\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__51868\,
            I => \N__51860\
        );

    \I__11882\ : InMux
    port map (
            O => \N__51865\,
            I => \N__51857\
        );

    \I__11881\ : Odrv4
    port map (
            O => \N__51860\,
            I => n1130
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__51857\,
            I => n1130
        );

    \I__11879\ : InMux
    port map (
            O => \N__51852\,
            I => \N__51849\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__51849\,
            I => n1197
        );

    \I__11877\ : InMux
    port map (
            O => \N__51846\,
            I => n12511
        );

    \I__11876\ : InMux
    port map (
            O => \N__51843\,
            I => \N__51839\
        );

    \I__11875\ : CascadeMux
    port map (
            O => \N__51842\,
            I => \N__51836\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__51839\,
            I => \N__51833\
        );

    \I__11873\ : InMux
    port map (
            O => \N__51836\,
            I => \N__51830\
        );

    \I__11872\ : Span4Mux_v
    port map (
            O => \N__51833\,
            I => \N__51825\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__51830\,
            I => \N__51825\
        );

    \I__11870\ : Span4Mux_h
    port map (
            O => \N__51825\,
            I => \N__51821\
        );

    \I__11869\ : InMux
    port map (
            O => \N__51824\,
            I => \N__51818\
        );

    \I__11868\ : Odrv4
    port map (
            O => \N__51821\,
            I => n1129
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__51818\,
            I => n1129
        );

    \I__11866\ : InMux
    port map (
            O => \N__51813\,
            I => \N__51810\
        );

    \I__11865\ : LocalMux
    port map (
            O => \N__51810\,
            I => n1196
        );

    \I__11864\ : InMux
    port map (
            O => \N__51807\,
            I => n12512
        );

    \I__11863\ : CascadeMux
    port map (
            O => \N__51804\,
            I => \N__51800\
        );

    \I__11862\ : CascadeMux
    port map (
            O => \N__51803\,
            I => \N__51797\
        );

    \I__11861\ : InMux
    port map (
            O => \N__51800\,
            I => \N__51794\
        );

    \I__11860\ : InMux
    port map (
            O => \N__51797\,
            I => \N__51791\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__51794\,
            I => \N__51788\
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__51791\,
            I => \N__51784\
        );

    \I__11857\ : Span4Mux_h
    port map (
            O => \N__51788\,
            I => \N__51781\
        );

    \I__11856\ : InMux
    port map (
            O => \N__51787\,
            I => \N__51778\
        );

    \I__11855\ : Odrv12
    port map (
            O => \N__51784\,
            I => n1128
        );

    \I__11854\ : Odrv4
    port map (
            O => \N__51781\,
            I => n1128
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__51778\,
            I => n1128
        );

    \I__11852\ : InMux
    port map (
            O => \N__51771\,
            I => \N__51768\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__51768\,
            I => n1195
        );

    \I__11850\ : InMux
    port map (
            O => \N__51765\,
            I => n12513
        );

    \I__11849\ : InMux
    port map (
            O => \N__51762\,
            I => \N__51758\
        );

    \I__11848\ : CascadeMux
    port map (
            O => \N__51761\,
            I => \N__51755\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__51758\,
            I => \N__51752\
        );

    \I__11846\ : InMux
    port map (
            O => \N__51755\,
            I => \N__51749\
        );

    \I__11845\ : Span4Mux_h
    port map (
            O => \N__51752\,
            I => \N__51745\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__51749\,
            I => \N__51742\
        );

    \I__11843\ : InMux
    port map (
            O => \N__51748\,
            I => \N__51739\
        );

    \I__11842\ : Odrv4
    port map (
            O => \N__51745\,
            I => n1127
        );

    \I__11841\ : Odrv12
    port map (
            O => \N__51742\,
            I => n1127
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__51739\,
            I => n1127
        );

    \I__11839\ : InMux
    port map (
            O => \N__51732\,
            I => \N__51729\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__51729\,
            I => n1194
        );

    \I__11837\ : InMux
    port map (
            O => \N__51726\,
            I => n12514
        );

    \I__11836\ : InMux
    port map (
            O => \N__51723\,
            I => \bfn_16_24_0_\
        );

    \I__11835\ : CascadeMux
    port map (
            O => \N__51720\,
            I => \N__51716\
        );

    \I__11834\ : CascadeMux
    port map (
            O => \N__51719\,
            I => \N__51713\
        );

    \I__11833\ : InMux
    port map (
            O => \N__51716\,
            I => \N__51710\
        );

    \I__11832\ : InMux
    port map (
            O => \N__51713\,
            I => \N__51707\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__51710\,
            I => \N__51704\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__51707\,
            I => n1226
        );

    \I__11829\ : Odrv4
    port map (
            O => \N__51704\,
            I => n1226
        );

    \I__11828\ : CascadeMux
    port map (
            O => \N__51699\,
            I => \n1226_cascade_\
        );

    \I__11827\ : InMux
    port map (
            O => \N__51696\,
            I => \N__51693\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__51693\,
            I => \N__51690\
        );

    \I__11825\ : Odrv4
    port map (
            O => \N__51690\,
            I => n1293
        );

    \I__11824\ : CascadeMux
    port map (
            O => \N__51687\,
            I => \N__51684\
        );

    \I__11823\ : InMux
    port map (
            O => \N__51684\,
            I => \N__51679\
        );

    \I__11822\ : InMux
    port map (
            O => \N__51683\,
            I => \N__51674\
        );

    \I__11821\ : InMux
    port map (
            O => \N__51682\,
            I => \N__51674\
        );

    \I__11820\ : LocalMux
    port map (
            O => \N__51679\,
            I => n1325
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__51674\,
            I => n1325
        );

    \I__11818\ : CascadeMux
    port map (
            O => \N__51669\,
            I => \N__51665\
        );

    \I__11817\ : InMux
    port map (
            O => \N__51668\,
            I => \N__51662\
        );

    \I__11816\ : InMux
    port map (
            O => \N__51665\,
            I => \N__51659\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__51662\,
            I => n1229
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__51659\,
            I => n1229
        );

    \I__11813\ : InMux
    port map (
            O => \N__51654\,
            I => \N__51651\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__51651\,
            I => \N__51648\
        );

    \I__11811\ : Span4Mux_h
    port map (
            O => \N__51648\,
            I => \N__51645\
        );

    \I__11810\ : Odrv4
    port map (
            O => \N__51645\,
            I => n11910
        );

    \I__11809\ : CascadeMux
    port map (
            O => \N__51642\,
            I => \n1229_cascade_\
        );

    \I__11808\ : InMux
    port map (
            O => \N__51639\,
            I => \N__51634\
        );

    \I__11807\ : InMux
    port map (
            O => \N__51638\,
            I => \N__51631\
        );

    \I__11806\ : CascadeMux
    port map (
            O => \N__51637\,
            I => \N__51628\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__51634\,
            I => \N__51625\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__51631\,
            I => \N__51622\
        );

    \I__11803\ : InMux
    port map (
            O => \N__51628\,
            I => \N__51619\
        );

    \I__11802\ : Span4Mux_h
    port map (
            O => \N__51625\,
            I => \N__51616\
        );

    \I__11801\ : Odrv4
    port map (
            O => \N__51622\,
            I => n1231
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__51619\,
            I => n1231
        );

    \I__11799\ : Odrv4
    port map (
            O => \N__51616\,
            I => n1231
        );

    \I__11798\ : InMux
    port map (
            O => \N__51609\,
            I => \N__51606\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__51606\,
            I => n13711
        );

    \I__11796\ : InMux
    port map (
            O => \N__51603\,
            I => \N__51598\
        );

    \I__11795\ : CascadeMux
    port map (
            O => \N__51602\,
            I => \N__51594\
        );

    \I__11794\ : CascadeMux
    port map (
            O => \N__51601\,
            I => \N__51591\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__51598\,
            I => \N__51586\
        );

    \I__11792\ : CascadeMux
    port map (
            O => \N__51597\,
            I => \N__51583\
        );

    \I__11791\ : InMux
    port map (
            O => \N__51594\,
            I => \N__51576\
        );

    \I__11790\ : InMux
    port map (
            O => \N__51591\,
            I => \N__51576\
        );

    \I__11789\ : InMux
    port map (
            O => \N__51590\,
            I => \N__51573\
        );

    \I__11788\ : CascadeMux
    port map (
            O => \N__51589\,
            I => \N__51570\
        );

    \I__11787\ : Span12Mux_h
    port map (
            O => \N__51586\,
            I => \N__51564\
        );

    \I__11786\ : InMux
    port map (
            O => \N__51583\,
            I => \N__51557\
        );

    \I__11785\ : InMux
    port map (
            O => \N__51582\,
            I => \N__51557\
        );

    \I__11784\ : InMux
    port map (
            O => \N__51581\,
            I => \N__51557\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__51576\,
            I => \N__51552\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__51573\,
            I => \N__51552\
        );

    \I__11781\ : InMux
    port map (
            O => \N__51570\,
            I => \N__51547\
        );

    \I__11780\ : InMux
    port map (
            O => \N__51569\,
            I => \N__51547\
        );

    \I__11779\ : InMux
    port map (
            O => \N__51568\,
            I => \N__51542\
        );

    \I__11778\ : InMux
    port map (
            O => \N__51567\,
            I => \N__51542\
        );

    \I__11777\ : Odrv12
    port map (
            O => \N__51564\,
            I => n1257
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__51557\,
            I => n1257
        );

    \I__11775\ : Odrv4
    port map (
            O => \N__51552\,
            I => n1257
        );

    \I__11774\ : LocalMux
    port map (
            O => \N__51547\,
            I => n1257
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__51542\,
            I => n1257
        );

    \I__11772\ : InMux
    port map (
            O => \N__51531\,
            I => \N__51528\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__51528\,
            I => \N__51525\
        );

    \I__11770\ : Span4Mux_h
    port map (
            O => \N__51525\,
            I => \N__51522\
        );

    \I__11769\ : Span4Mux_h
    port map (
            O => \N__51522\,
            I => \N__51518\
        );

    \I__11768\ : InMux
    port map (
            O => \N__51521\,
            I => \N__51515\
        );

    \I__11767\ : Span4Mux_h
    port map (
            O => \N__51518\,
            I => \N__51510\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__51515\,
            I => \N__51510\
        );

    \I__11765\ : Odrv4
    port map (
            O => \N__51510\,
            I => n15528
        );

    \I__11764\ : CascadeMux
    port map (
            O => \N__51507\,
            I => \N__51502\
        );

    \I__11763\ : InMux
    port map (
            O => \N__51506\,
            I => \N__51497\
        );

    \I__11762\ : InMux
    port map (
            O => \N__51505\,
            I => \N__51497\
        );

    \I__11761\ : InMux
    port map (
            O => \N__51502\,
            I => \N__51494\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__51497\,
            I => n1228
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__51494\,
            I => n1228
        );

    \I__11758\ : CascadeMux
    port map (
            O => \N__51489\,
            I => \N__51484\
        );

    \I__11757\ : InMux
    port map (
            O => \N__51488\,
            I => \N__51481\
        );

    \I__11756\ : InMux
    port map (
            O => \N__51487\,
            I => \N__51478\
        );

    \I__11755\ : InMux
    port map (
            O => \N__51484\,
            I => \N__51475\
        );

    \I__11754\ : LocalMux
    port map (
            O => \N__51481\,
            I => n1230
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__51478\,
            I => n1230
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__51475\,
            I => n1230
        );

    \I__11751\ : CascadeMux
    port map (
            O => \N__51468\,
            I => \N__51465\
        );

    \I__11750\ : InMux
    port map (
            O => \N__51465\,
            I => \N__51460\
        );

    \I__11749\ : InMux
    port map (
            O => \N__51464\,
            I => \N__51455\
        );

    \I__11748\ : InMux
    port map (
            O => \N__51463\,
            I => \N__51455\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__51460\,
            I => \N__51452\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__51455\,
            I => \N__51449\
        );

    \I__11745\ : Span4Mux_h
    port map (
            O => \N__51452\,
            I => \N__51446\
        );

    \I__11744\ : Odrv4
    port map (
            O => \N__51449\,
            I => n297
        );

    \I__11743\ : Odrv4
    port map (
            O => \N__51446\,
            I => n297
        );

    \I__11742\ : InMux
    port map (
            O => \N__51441\,
            I => \N__51438\
        );

    \I__11741\ : LocalMux
    port map (
            O => \N__51438\,
            I => \N__51435\
        );

    \I__11740\ : Odrv12
    port map (
            O => \N__51435\,
            I => n1201
        );

    \I__11739\ : InMux
    port map (
            O => \N__51432\,
            I => \bfn_16_23_0_\
        );

    \I__11738\ : CascadeMux
    port map (
            O => \N__51429\,
            I => \N__51425\
        );

    \I__11737\ : CascadeMux
    port map (
            O => \N__51428\,
            I => \N__51422\
        );

    \I__11736\ : InMux
    port map (
            O => \N__51425\,
            I => \N__51419\
        );

    \I__11735\ : InMux
    port map (
            O => \N__51422\,
            I => \N__51416\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__51419\,
            I => \N__51413\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__51416\,
            I => \N__51410\
        );

    \I__11732\ : Odrv4
    port map (
            O => \N__51413\,
            I => n1133
        );

    \I__11731\ : Odrv4
    port map (
            O => \N__51410\,
            I => n1133
        );

    \I__11730\ : InMux
    port map (
            O => \N__51405\,
            I => \N__51402\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__51402\,
            I => \N__51394\
        );

    \I__11728\ : CascadeMux
    port map (
            O => \N__51401\,
            I => \N__51388\
        );

    \I__11727\ : CascadeMux
    port map (
            O => \N__51400\,
            I => \N__51383\
        );

    \I__11726\ : CascadeMux
    port map (
            O => \N__51399\,
            I => \N__51380\
        );

    \I__11725\ : CascadeMux
    port map (
            O => \N__51398\,
            I => \N__51376\
        );

    \I__11724\ : InMux
    port map (
            O => \N__51397\,
            I => \N__51372\
        );

    \I__11723\ : Span12Mux_h
    port map (
            O => \N__51394\,
            I => \N__51369\
        );

    \I__11722\ : InMux
    port map (
            O => \N__51393\,
            I => \N__51366\
        );

    \I__11721\ : InMux
    port map (
            O => \N__51392\,
            I => \N__51363\
        );

    \I__11720\ : InMux
    port map (
            O => \N__51391\,
            I => \N__51358\
        );

    \I__11719\ : InMux
    port map (
            O => \N__51388\,
            I => \N__51358\
        );

    \I__11718\ : InMux
    port map (
            O => \N__51387\,
            I => \N__51351\
        );

    \I__11717\ : InMux
    port map (
            O => \N__51386\,
            I => \N__51351\
        );

    \I__11716\ : InMux
    port map (
            O => \N__51383\,
            I => \N__51351\
        );

    \I__11715\ : InMux
    port map (
            O => \N__51380\,
            I => \N__51342\
        );

    \I__11714\ : InMux
    port map (
            O => \N__51379\,
            I => \N__51342\
        );

    \I__11713\ : InMux
    port map (
            O => \N__51376\,
            I => \N__51342\
        );

    \I__11712\ : InMux
    port map (
            O => \N__51375\,
            I => \N__51342\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__51372\,
            I => \N__51339\
        );

    \I__11710\ : Odrv12
    port map (
            O => \N__51369\,
            I => n1455
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__51366\,
            I => n1455
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__51363\,
            I => n1455
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__51358\,
            I => n1455
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__51351\,
            I => n1455
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__51342\,
            I => n1455
        );

    \I__11704\ : Odrv4
    port map (
            O => \N__51339\,
            I => n1455
        );

    \I__11703\ : InMux
    port map (
            O => \N__51324\,
            I => \N__51321\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__51321\,
            I => \N__51318\
        );

    \I__11701\ : Span12Mux_h
    port map (
            O => \N__51318\,
            I => \N__51314\
        );

    \I__11700\ : InMux
    port map (
            O => \N__51317\,
            I => \N__51311\
        );

    \I__11699\ : Odrv12
    port map (
            O => \N__51314\,
            I => n15562
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__51311\,
            I => n15562
        );

    \I__11697\ : InMux
    port map (
            O => \N__51306\,
            I => \N__51303\
        );

    \I__11696\ : LocalMux
    port map (
            O => \N__51303\,
            I => n1392
        );

    \I__11695\ : InMux
    port map (
            O => \N__51300\,
            I => \N__51297\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__51297\,
            I => \N__51291\
        );

    \I__11693\ : InMux
    port map (
            O => \N__51296\,
            I => \N__51288\
        );

    \I__11692\ : CascadeMux
    port map (
            O => \N__51295\,
            I => \N__51284\
        );

    \I__11691\ : InMux
    port map (
            O => \N__51294\,
            I => \N__51278\
        );

    \I__11690\ : Span4Mux_h
    port map (
            O => \N__51291\,
            I => \N__51274\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__51288\,
            I => \N__51271\
        );

    \I__11688\ : CascadeMux
    port map (
            O => \N__51287\,
            I => \N__51267\
        );

    \I__11687\ : InMux
    port map (
            O => \N__51284\,
            I => \N__51261\
        );

    \I__11686\ : InMux
    port map (
            O => \N__51283\,
            I => \N__51261\
        );

    \I__11685\ : InMux
    port map (
            O => \N__51282\,
            I => \N__51258\
        );

    \I__11684\ : InMux
    port map (
            O => \N__51281\,
            I => \N__51255\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__51278\,
            I => \N__51252\
        );

    \I__11682\ : CascadeMux
    port map (
            O => \N__51277\,
            I => \N__51249\
        );

    \I__11681\ : Span4Mux_h
    port map (
            O => \N__51274\,
            I => \N__51243\
        );

    \I__11680\ : Span4Mux_h
    port map (
            O => \N__51271\,
            I => \N__51243\
        );

    \I__11679\ : InMux
    port map (
            O => \N__51270\,
            I => \N__51236\
        );

    \I__11678\ : InMux
    port map (
            O => \N__51267\,
            I => \N__51236\
        );

    \I__11677\ : InMux
    port map (
            O => \N__51266\,
            I => \N__51236\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__51261\,
            I => \N__51227\
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__51258\,
            I => \N__51227\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__51255\,
            I => \N__51227\
        );

    \I__11673\ : Span4Mux_h
    port map (
            O => \N__51252\,
            I => \N__51227\
        );

    \I__11672\ : InMux
    port map (
            O => \N__51249\,
            I => \N__51222\
        );

    \I__11671\ : InMux
    port map (
            O => \N__51248\,
            I => \N__51222\
        );

    \I__11670\ : Odrv4
    port map (
            O => \N__51243\,
            I => n1356
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__51236\,
            I => n1356
        );

    \I__11668\ : Odrv4
    port map (
            O => \N__51227\,
            I => n1356
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__51222\,
            I => n1356
        );

    \I__11666\ : CascadeMux
    port map (
            O => \N__51213\,
            I => \N__51208\
        );

    \I__11665\ : InMux
    port map (
            O => \N__51212\,
            I => \N__51205\
        );

    \I__11664\ : InMux
    port map (
            O => \N__51211\,
            I => \N__51202\
        );

    \I__11663\ : InMux
    port map (
            O => \N__51208\,
            I => \N__51199\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__51205\,
            I => \N__51194\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__51202\,
            I => \N__51194\
        );

    \I__11660\ : LocalMux
    port map (
            O => \N__51199\,
            I => n1424
        );

    \I__11659\ : Odrv4
    port map (
            O => \N__51194\,
            I => n1424
        );

    \I__11658\ : InMux
    port map (
            O => \N__51189\,
            I => \N__51186\
        );

    \I__11657\ : LocalMux
    port map (
            O => \N__51186\,
            I => \N__51183\
        );

    \I__11656\ : Odrv4
    port map (
            O => \N__51183\,
            I => n1294
        );

    \I__11655\ : CascadeMux
    port map (
            O => \N__51180\,
            I => \N__51177\
        );

    \I__11654\ : InMux
    port map (
            O => \N__51177\,
            I => \N__51174\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__51174\,
            I => \N__51171\
        );

    \I__11652\ : Odrv4
    port map (
            O => \N__51171\,
            I => n1295
        );

    \I__11651\ : InMux
    port map (
            O => \N__51168\,
            I => \N__51161\
        );

    \I__11650\ : InMux
    port map (
            O => \N__51167\,
            I => \N__51161\
        );

    \I__11649\ : InMux
    port map (
            O => \N__51166\,
            I => \N__51158\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__51161\,
            I => n1227
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__51158\,
            I => n1227
        );

    \I__11646\ : CascadeMux
    port map (
            O => \N__51153\,
            I => \n14482_cascade_\
        );

    \I__11645\ : InMux
    port map (
            O => \N__51150\,
            I => \N__51147\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__51147\,
            I => \N__51144\
        );

    \I__11643\ : Odrv4
    port map (
            O => \N__51144\,
            I => n1296
        );

    \I__11642\ : CascadeMux
    port map (
            O => \N__51141\,
            I => \n1257_cascade_\
        );

    \I__11641\ : InMux
    port map (
            O => \N__51138\,
            I => \N__51134\
        );

    \I__11640\ : CascadeMux
    port map (
            O => \N__51137\,
            I => \N__51131\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__51134\,
            I => \N__51128\
        );

    \I__11638\ : InMux
    port map (
            O => \N__51131\,
            I => \N__51125\
        );

    \I__11637\ : Odrv4
    port map (
            O => \N__51128\,
            I => n1328
        );

    \I__11636\ : LocalMux
    port map (
            O => \N__51125\,
            I => n1328
        );

    \I__11635\ : InMux
    port map (
            O => \N__51120\,
            I => \N__51115\
        );

    \I__11634\ : InMux
    port map (
            O => \N__51119\,
            I => \N__51112\
        );

    \I__11633\ : InMux
    port map (
            O => \N__51118\,
            I => \N__51109\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__51115\,
            I => n1327
        );

    \I__11631\ : LocalMux
    port map (
            O => \N__51112\,
            I => n1327
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__51109\,
            I => n1327
        );

    \I__11629\ : CascadeMux
    port map (
            O => \N__51102\,
            I => \n1328_cascade_\
        );

    \I__11628\ : CascadeMux
    port map (
            O => \N__51099\,
            I => \N__51095\
        );

    \I__11627\ : CascadeMux
    port map (
            O => \N__51098\,
            I => \N__51092\
        );

    \I__11626\ : InMux
    port map (
            O => \N__51095\,
            I => \N__51088\
        );

    \I__11625\ : InMux
    port map (
            O => \N__51092\,
            I => \N__51085\
        );

    \I__11624\ : InMux
    port map (
            O => \N__51091\,
            I => \N__51082\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__51088\,
            I => n1326
        );

    \I__11622\ : LocalMux
    port map (
            O => \N__51085\,
            I => n1326
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__51082\,
            I => n1326
        );

    \I__11620\ : InMux
    port map (
            O => \N__51075\,
            I => \N__51072\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__51072\,
            I => \N__51069\
        );

    \I__11618\ : Span4Mux_h
    port map (
            O => \N__51069\,
            I => \N__51066\
        );

    \I__11617\ : Odrv4
    port map (
            O => \N__51066\,
            I => n14282
        );

    \I__11616\ : CascadeMux
    port map (
            O => \N__51063\,
            I => \N__51060\
        );

    \I__11615\ : InMux
    port map (
            O => \N__51060\,
            I => \N__51057\
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__51057\,
            I => \N__51052\
        );

    \I__11613\ : InMux
    port map (
            O => \N__51056\,
            I => \N__51049\
        );

    \I__11612\ : InMux
    port map (
            O => \N__51055\,
            I => \N__51046\
        );

    \I__11611\ : Span4Mux_h
    port map (
            O => \N__51052\,
            I => \N__51043\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__51049\,
            I => n1429
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__51046\,
            I => n1429
        );

    \I__11608\ : Odrv4
    port map (
            O => \N__51043\,
            I => n1429
        );

    \I__11607\ : InMux
    port map (
            O => \N__51036\,
            I => \N__51033\
        );

    \I__11606\ : LocalMux
    port map (
            O => \N__51033\,
            I => \N__51030\
        );

    \I__11605\ : Odrv4
    port map (
            O => \N__51030\,
            I => n1496
        );

    \I__11604\ : InMux
    port map (
            O => \N__51027\,
            I => n12542
        );

    \I__11603\ : CascadeMux
    port map (
            O => \N__51024\,
            I => \N__51021\
        );

    \I__11602\ : InMux
    port map (
            O => \N__51021\,
            I => \N__51017\
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__51020\,
            I => \N__51013\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__51017\,
            I => \N__51010\
        );

    \I__11599\ : InMux
    port map (
            O => \N__51016\,
            I => \N__51007\
        );

    \I__11598\ : InMux
    port map (
            O => \N__51013\,
            I => \N__51004\
        );

    \I__11597\ : Span4Mux_v
    port map (
            O => \N__51010\,
            I => \N__51001\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__51007\,
            I => n1428
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__51004\,
            I => n1428
        );

    \I__11594\ : Odrv4
    port map (
            O => \N__51001\,
            I => n1428
        );

    \I__11593\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50991\
        );

    \I__11592\ : LocalMux
    port map (
            O => \N__50991\,
            I => \N__50988\
        );

    \I__11591\ : Span4Mux_h
    port map (
            O => \N__50988\,
            I => \N__50985\
        );

    \I__11590\ : Odrv4
    port map (
            O => \N__50985\,
            I => n1495
        );

    \I__11589\ : InMux
    port map (
            O => \N__50982\,
            I => n12543
        );

    \I__11588\ : CascadeMux
    port map (
            O => \N__50979\,
            I => \N__50975\
        );

    \I__11587\ : InMux
    port map (
            O => \N__50978\,
            I => \N__50972\
        );

    \I__11586\ : InMux
    port map (
            O => \N__50975\,
            I => \N__50969\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__50972\,
            I => \N__50966\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__50969\,
            I => n1427
        );

    \I__11583\ : Odrv4
    port map (
            O => \N__50966\,
            I => n1427
        );

    \I__11582\ : InMux
    port map (
            O => \N__50961\,
            I => \N__50958\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__50958\,
            I => n1494
        );

    \I__11580\ : InMux
    port map (
            O => \N__50955\,
            I => n12544
        );

    \I__11579\ : CascadeMux
    port map (
            O => \N__50952\,
            I => \N__50949\
        );

    \I__11578\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50944\
        );

    \I__11577\ : InMux
    port map (
            O => \N__50948\,
            I => \N__50939\
        );

    \I__11576\ : InMux
    port map (
            O => \N__50947\,
            I => \N__50939\
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__50944\,
            I => n1426
        );

    \I__11574\ : LocalMux
    port map (
            O => \N__50939\,
            I => n1426
        );

    \I__11573\ : InMux
    port map (
            O => \N__50934\,
            I => \N__50931\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__50931\,
            I => n1493
        );

    \I__11571\ : InMux
    port map (
            O => \N__50928\,
            I => \bfn_16_20_0_\
        );

    \I__11570\ : CascadeMux
    port map (
            O => \N__50925\,
            I => \N__50922\
        );

    \I__11569\ : InMux
    port map (
            O => \N__50922\,
            I => \N__50917\
        );

    \I__11568\ : InMux
    port map (
            O => \N__50921\,
            I => \N__50912\
        );

    \I__11567\ : InMux
    port map (
            O => \N__50920\,
            I => \N__50912\
        );

    \I__11566\ : LocalMux
    port map (
            O => \N__50917\,
            I => n1425
        );

    \I__11565\ : LocalMux
    port map (
            O => \N__50912\,
            I => n1425
        );

    \I__11564\ : CascadeMux
    port map (
            O => \N__50907\,
            I => \N__50904\
        );

    \I__11563\ : InMux
    port map (
            O => \N__50904\,
            I => \N__50901\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__50901\,
            I => n1492
        );

    \I__11561\ : InMux
    port map (
            O => \N__50898\,
            I => n12546
        );

    \I__11560\ : InMux
    port map (
            O => \N__50895\,
            I => \N__50892\
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__50892\,
            I => n1491
        );

    \I__11558\ : InMux
    port map (
            O => \N__50889\,
            I => n12547
        );

    \I__11557\ : CascadeMux
    port map (
            O => \N__50886\,
            I => \N__50883\
        );

    \I__11556\ : InMux
    port map (
            O => \N__50883\,
            I => \N__50880\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__50880\,
            I => \N__50876\
        );

    \I__11554\ : InMux
    port map (
            O => \N__50879\,
            I => \N__50872\
        );

    \I__11553\ : Span4Mux_h
    port map (
            O => \N__50876\,
            I => \N__50869\
        );

    \I__11552\ : InMux
    port map (
            O => \N__50875\,
            I => \N__50866\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__50872\,
            I => n1423
        );

    \I__11550\ : Odrv4
    port map (
            O => \N__50869\,
            I => n1423
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__50866\,
            I => n1423
        );

    \I__11548\ : CascadeMux
    port map (
            O => \N__50859\,
            I => \N__50856\
        );

    \I__11547\ : InMux
    port map (
            O => \N__50856\,
            I => \N__50853\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__50853\,
            I => \N__50850\
        );

    \I__11545\ : Odrv4
    port map (
            O => \N__50850\,
            I => n1490
        );

    \I__11544\ : InMux
    port map (
            O => \N__50847\,
            I => n12548
        );

    \I__11543\ : CascadeMux
    port map (
            O => \N__50844\,
            I => \N__50841\
        );

    \I__11542\ : InMux
    port map (
            O => \N__50841\,
            I => \N__50837\
        );

    \I__11541\ : InMux
    port map (
            O => \N__50840\,
            I => \N__50834\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__50837\,
            I => \N__50831\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__50834\,
            I => \N__50828\
        );

    \I__11538\ : Odrv4
    port map (
            O => \N__50831\,
            I => n1422
        );

    \I__11537\ : Odrv4
    port map (
            O => \N__50828\,
            I => n1422
        );

    \I__11536\ : InMux
    port map (
            O => \N__50823\,
            I => n12549
        );

    \I__11535\ : CascadeMux
    port map (
            O => \N__50820\,
            I => \N__50817\
        );

    \I__11534\ : InMux
    port map (
            O => \N__50817\,
            I => \N__50814\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__50814\,
            I => \N__50810\
        );

    \I__11532\ : InMux
    port map (
            O => \N__50813\,
            I => \N__50807\
        );

    \I__11531\ : Odrv4
    port map (
            O => \N__50810\,
            I => n1521
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__50807\,
            I => n1521
        );

    \I__11529\ : InMux
    port map (
            O => \N__50802\,
            I => \N__50799\
        );

    \I__11528\ : LocalMux
    port map (
            O => \N__50799\,
            I => \N__50795\
        );

    \I__11527\ : CascadeMux
    port map (
            O => \N__50798\,
            I => \N__50792\
        );

    \I__11526\ : Span4Mux_h
    port map (
            O => \N__50795\,
            I => \N__50789\
        );

    \I__11525\ : InMux
    port map (
            O => \N__50792\,
            I => \N__50786\
        );

    \I__11524\ : Odrv4
    port map (
            O => \N__50789\,
            I => n1527
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__50786\,
            I => n1527
        );

    \I__11522\ : InMux
    port map (
            O => \N__50781\,
            I => \N__50778\
        );

    \I__11521\ : LocalMux
    port map (
            O => \N__50778\,
            I => \N__50775\
        );

    \I__11520\ : Span4Mux_h
    port map (
            O => \N__50775\,
            I => \N__50772\
        );

    \I__11519\ : Odrv4
    port map (
            O => \N__50772\,
            I => n1594
        );

    \I__11518\ : CascadeMux
    port map (
            O => \N__50769\,
            I => \N__50766\
        );

    \I__11517\ : InMux
    port map (
            O => \N__50766\,
            I => \N__50761\
        );

    \I__11516\ : InMux
    port map (
            O => \N__50765\,
            I => \N__50756\
        );

    \I__11515\ : InMux
    port map (
            O => \N__50764\,
            I => \N__50756\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__50761\,
            I => n1626_adj_613
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__50756\,
            I => n1626_adj_613
        );

    \I__11512\ : CascadeMux
    port map (
            O => \N__50751\,
            I => \N__50748\
        );

    \I__11511\ : InMux
    port map (
            O => \N__50748\,
            I => \N__50743\
        );

    \I__11510\ : InMux
    port map (
            O => \N__50747\,
            I => \N__50740\
        );

    \I__11509\ : InMux
    port map (
            O => \N__50746\,
            I => \N__50737\
        );

    \I__11508\ : LocalMux
    port map (
            O => \N__50743\,
            I => \N__50734\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__50740\,
            I => n1529
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__50737\,
            I => n1529
        );

    \I__11505\ : Odrv4
    port map (
            O => \N__50734\,
            I => n1529
        );

    \I__11504\ : CascadeMux
    port map (
            O => \N__50727\,
            I => \N__50724\
        );

    \I__11503\ : InMux
    port map (
            O => \N__50724\,
            I => \N__50721\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__50721\,
            I => \N__50718\
        );

    \I__11501\ : Span4Mux_h
    port map (
            O => \N__50718\,
            I => \N__50715\
        );

    \I__11500\ : Odrv4
    port map (
            O => \N__50715\,
            I => n1596
        );

    \I__11499\ : CascadeMux
    port map (
            O => \N__50712\,
            I => \N__50708\
        );

    \I__11498\ : CascadeMux
    port map (
            O => \N__50711\,
            I => \N__50705\
        );

    \I__11497\ : InMux
    port map (
            O => \N__50708\,
            I => \N__50701\
        );

    \I__11496\ : InMux
    port map (
            O => \N__50705\,
            I => \N__50698\
        );

    \I__11495\ : InMux
    port map (
            O => \N__50704\,
            I => \N__50695\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__50701\,
            I => n1628_adj_615
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__50698\,
            I => n1628_adj_615
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__50695\,
            I => n1628_adj_615
        );

    \I__11491\ : InMux
    port map (
            O => \N__50688\,
            I => \N__50685\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__50685\,
            I => \N__50682\
        );

    \I__11489\ : Span4Mux_h
    port map (
            O => \N__50682\,
            I => \N__50679\
        );

    \I__11488\ : Odrv4
    port map (
            O => \N__50679\,
            I => n1597
        );

    \I__11487\ : InMux
    port map (
            O => \N__50676\,
            I => \N__50673\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__50673\,
            I => \N__50669\
        );

    \I__11485\ : InMux
    port map (
            O => \N__50672\,
            I => \N__50663\
        );

    \I__11484\ : Sp12to4
    port map (
            O => \N__50669\,
            I => \N__50658\
        );

    \I__11483\ : InMux
    port map (
            O => \N__50668\,
            I => \N__50655\
        );

    \I__11482\ : CascadeMux
    port map (
            O => \N__50667\,
            I => \N__50649\
        );

    \I__11481\ : CascadeMux
    port map (
            O => \N__50666\,
            I => \N__50643\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__50663\,
            I => \N__50640\
        );

    \I__11479\ : CascadeMux
    port map (
            O => \N__50662\,
            I => \N__50637\
        );

    \I__11478\ : CascadeMux
    port map (
            O => \N__50661\,
            I => \N__50634\
        );

    \I__11477\ : Span12Mux_v
    port map (
            O => \N__50658\,
            I => \N__50629\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__50655\,
            I => \N__50626\
        );

    \I__11475\ : InMux
    port map (
            O => \N__50654\,
            I => \N__50623\
        );

    \I__11474\ : InMux
    port map (
            O => \N__50653\,
            I => \N__50618\
        );

    \I__11473\ : InMux
    port map (
            O => \N__50652\,
            I => \N__50618\
        );

    \I__11472\ : InMux
    port map (
            O => \N__50649\,
            I => \N__50607\
        );

    \I__11471\ : InMux
    port map (
            O => \N__50648\,
            I => \N__50607\
        );

    \I__11470\ : InMux
    port map (
            O => \N__50647\,
            I => \N__50607\
        );

    \I__11469\ : InMux
    port map (
            O => \N__50646\,
            I => \N__50607\
        );

    \I__11468\ : InMux
    port map (
            O => \N__50643\,
            I => \N__50607\
        );

    \I__11467\ : Span4Mux_h
    port map (
            O => \N__50640\,
            I => \N__50604\
        );

    \I__11466\ : InMux
    port map (
            O => \N__50637\,
            I => \N__50595\
        );

    \I__11465\ : InMux
    port map (
            O => \N__50634\,
            I => \N__50595\
        );

    \I__11464\ : InMux
    port map (
            O => \N__50633\,
            I => \N__50595\
        );

    \I__11463\ : InMux
    port map (
            O => \N__50632\,
            I => \N__50595\
        );

    \I__11462\ : Odrv12
    port map (
            O => \N__50629\,
            I => n1554
        );

    \I__11461\ : Odrv4
    port map (
            O => \N__50626\,
            I => n1554
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__50623\,
            I => n1554
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__50618\,
            I => n1554
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__50607\,
            I => n1554
        );

    \I__11457\ : Odrv4
    port map (
            O => \N__50604\,
            I => n1554
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__50595\,
            I => n1554
        );

    \I__11455\ : CascadeMux
    port map (
            O => \N__50580\,
            I => \N__50577\
        );

    \I__11454\ : InMux
    port map (
            O => \N__50577\,
            I => \N__50572\
        );

    \I__11453\ : InMux
    port map (
            O => \N__50576\,
            I => \N__50569\
        );

    \I__11452\ : InMux
    port map (
            O => \N__50575\,
            I => \N__50566\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__50572\,
            I => \N__50563\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__50569\,
            I => n1530
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__50566\,
            I => n1530
        );

    \I__11448\ : Odrv4
    port map (
            O => \N__50563\,
            I => n1530
        );

    \I__11447\ : CascadeMux
    port map (
            O => \N__50556\,
            I => \N__50551\
        );

    \I__11446\ : CascadeMux
    port map (
            O => \N__50555\,
            I => \N__50548\
        );

    \I__11445\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50545\
        );

    \I__11444\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50542\
        );

    \I__11443\ : InMux
    port map (
            O => \N__50548\,
            I => \N__50539\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__50545\,
            I => \N__50536\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__50542\,
            I => n1629_adj_616
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__50539\,
            I => n1629_adj_616
        );

    \I__11439\ : Odrv4
    port map (
            O => \N__50536\,
            I => n1629_adj_616
        );

    \I__11438\ : InMux
    port map (
            O => \N__50529\,
            I => \N__50525\
        );

    \I__11437\ : InMux
    port map (
            O => \N__50528\,
            I => \N__50522\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__50525\,
            I => \N__50516\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__50522\,
            I => \N__50516\
        );

    \I__11434\ : InMux
    port map (
            O => \N__50521\,
            I => \N__50513\
        );

    \I__11433\ : Span4Mux_h
    port map (
            O => \N__50516\,
            I => \N__50510\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__50513\,
            I => \N__50507\
        );

    \I__11431\ : Odrv4
    port map (
            O => \N__50510\,
            I => n300
        );

    \I__11430\ : Odrv4
    port map (
            O => \N__50507\,
            I => n300
        );

    \I__11429\ : InMux
    port map (
            O => \N__50502\,
            I => \N__50499\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__50499\,
            I => \N__50496\
        );

    \I__11427\ : Odrv12
    port map (
            O => \N__50496\,
            I => n1501
        );

    \I__11426\ : InMux
    port map (
            O => \N__50493\,
            I => \bfn_16_19_0_\
        );

    \I__11425\ : CascadeMux
    port map (
            O => \N__50490\,
            I => \N__50486\
        );

    \I__11424\ : CascadeMux
    port map (
            O => \N__50489\,
            I => \N__50483\
        );

    \I__11423\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50480\
        );

    \I__11422\ : InMux
    port map (
            O => \N__50483\,
            I => \N__50477\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__50480\,
            I => \N__50472\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__50477\,
            I => \N__50472\
        );

    \I__11419\ : Span4Mux_h
    port map (
            O => \N__50472\,
            I => \N__50469\
        );

    \I__11418\ : Odrv4
    port map (
            O => \N__50469\,
            I => n1433
        );

    \I__11417\ : InMux
    port map (
            O => \N__50466\,
            I => \N__50463\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__50463\,
            I => n1500
        );

    \I__11415\ : InMux
    port map (
            O => \N__50460\,
            I => n12538
        );

    \I__11414\ : CascadeMux
    port map (
            O => \N__50457\,
            I => \N__50454\
        );

    \I__11413\ : InMux
    port map (
            O => \N__50454\,
            I => \N__50450\
        );

    \I__11412\ : InMux
    port map (
            O => \N__50453\,
            I => \N__50447\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__50450\,
            I => \N__50444\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__50447\,
            I => \N__50440\
        );

    \I__11409\ : Span4Mux_v
    port map (
            O => \N__50444\,
            I => \N__50437\
        );

    \I__11408\ : InMux
    port map (
            O => \N__50443\,
            I => \N__50434\
        );

    \I__11407\ : Odrv4
    port map (
            O => \N__50440\,
            I => n1432
        );

    \I__11406\ : Odrv4
    port map (
            O => \N__50437\,
            I => n1432
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__50434\,
            I => n1432
        );

    \I__11404\ : InMux
    port map (
            O => \N__50427\,
            I => \N__50424\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__50424\,
            I => \N__50421\
        );

    \I__11402\ : Odrv4
    port map (
            O => \N__50421\,
            I => n1499
        );

    \I__11401\ : InMux
    port map (
            O => \N__50418\,
            I => n12539
        );

    \I__11400\ : CascadeMux
    port map (
            O => \N__50415\,
            I => \N__50411\
        );

    \I__11399\ : InMux
    port map (
            O => \N__50414\,
            I => \N__50407\
        );

    \I__11398\ : InMux
    port map (
            O => \N__50411\,
            I => \N__50404\
        );

    \I__11397\ : InMux
    port map (
            O => \N__50410\,
            I => \N__50401\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__50407\,
            I => n1431
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__50404\,
            I => n1431
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__50401\,
            I => n1431
        );

    \I__11393\ : InMux
    port map (
            O => \N__50394\,
            I => \N__50391\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__50391\,
            I => n1498
        );

    \I__11391\ : InMux
    port map (
            O => \N__50388\,
            I => n12540
        );

    \I__11390\ : CascadeMux
    port map (
            O => \N__50385\,
            I => \N__50381\
        );

    \I__11389\ : CascadeMux
    port map (
            O => \N__50384\,
            I => \N__50378\
        );

    \I__11388\ : InMux
    port map (
            O => \N__50381\,
            I => \N__50375\
        );

    \I__11387\ : InMux
    port map (
            O => \N__50378\,
            I => \N__50372\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__50375\,
            I => \N__50366\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__50372\,
            I => \N__50366\
        );

    \I__11384\ : InMux
    port map (
            O => \N__50371\,
            I => \N__50363\
        );

    \I__11383\ : Span4Mux_h
    port map (
            O => \N__50366\,
            I => \N__50360\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__50363\,
            I => n1430
        );

    \I__11381\ : Odrv4
    port map (
            O => \N__50360\,
            I => n1430
        );

    \I__11380\ : InMux
    port map (
            O => \N__50355\,
            I => \N__50352\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__50352\,
            I => n1497
        );

    \I__11378\ : InMux
    port map (
            O => \N__50349\,
            I => n12541
        );

    \I__11377\ : CascadeMux
    port map (
            O => \N__50346\,
            I => \n1727_cascade_\
        );

    \I__11376\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50340\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__50340\,
            I => \N__50335\
        );

    \I__11374\ : CascadeMux
    port map (
            O => \N__50339\,
            I => \N__50332\
        );

    \I__11373\ : InMux
    port map (
            O => \N__50338\,
            I => \N__50329\
        );

    \I__11372\ : Span4Mux_h
    port map (
            O => \N__50335\,
            I => \N__50326\
        );

    \I__11371\ : InMux
    port map (
            O => \N__50332\,
            I => \N__50323\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__50329\,
            I => \N__50320\
        );

    \I__11369\ : Odrv4
    port map (
            O => \N__50326\,
            I => n1726
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__50323\,
            I => n1726
        );

    \I__11367\ : Odrv4
    port map (
            O => \N__50320\,
            I => n1726
        );

    \I__11366\ : InMux
    port map (
            O => \N__50313\,
            I => \N__50309\
        );

    \I__11365\ : CascadeMux
    port map (
            O => \N__50312\,
            I => \N__50306\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__50309\,
            I => \N__50303\
        );

    \I__11363\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50300\
        );

    \I__11362\ : Span4Mux_h
    port map (
            O => \N__50303\,
            I => \N__50294\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__50300\,
            I => \N__50294\
        );

    \I__11360\ : InMux
    port map (
            O => \N__50299\,
            I => \N__50291\
        );

    \I__11359\ : Odrv4
    port map (
            O => \N__50294\,
            I => n1724
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__50291\,
            I => n1724
        );

    \I__11357\ : InMux
    port map (
            O => \N__50286\,
            I => \N__50282\
        );

    \I__11356\ : CascadeMux
    port map (
            O => \N__50285\,
            I => \N__50279\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__50282\,
            I => \N__50276\
        );

    \I__11354\ : InMux
    port map (
            O => \N__50279\,
            I => \N__50273\
        );

    \I__11353\ : Span4Mux_h
    port map (
            O => \N__50276\,
            I => \N__50268\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__50273\,
            I => \N__50268\
        );

    \I__11351\ : Span4Mux_h
    port map (
            O => \N__50268\,
            I => \N__50264\
        );

    \I__11350\ : InMux
    port map (
            O => \N__50267\,
            I => \N__50261\
        );

    \I__11349\ : Odrv4
    port map (
            O => \N__50264\,
            I => n1725
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__50261\,
            I => n1725
        );

    \I__11347\ : CascadeMux
    port map (
            O => \N__50256\,
            I => \n14166_cascade_\
        );

    \I__11346\ : InMux
    port map (
            O => \N__50253\,
            I => \N__50250\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__50250\,
            I => \N__50245\
        );

    \I__11344\ : CascadeMux
    port map (
            O => \N__50249\,
            I => \N__50242\
        );

    \I__11343\ : InMux
    port map (
            O => \N__50248\,
            I => \N__50239\
        );

    \I__11342\ : Span4Mux_h
    port map (
            O => \N__50245\,
            I => \N__50236\
        );

    \I__11341\ : InMux
    port map (
            O => \N__50242\,
            I => \N__50233\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__50239\,
            I => \N__50230\
        );

    \I__11339\ : Odrv4
    port map (
            O => \N__50236\,
            I => n1723
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__50233\,
            I => n1723
        );

    \I__11337\ : Odrv4
    port map (
            O => \N__50230\,
            I => n1723
        );

    \I__11336\ : InMux
    port map (
            O => \N__50223\,
            I => \N__50220\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__50220\,
            I => \N__50217\
        );

    \I__11334\ : Span4Mux_v
    port map (
            O => \N__50217\,
            I => \N__50214\
        );

    \I__11333\ : Span4Mux_h
    port map (
            O => \N__50214\,
            I => \N__50211\
        );

    \I__11332\ : Odrv4
    port map (
            O => \N__50211\,
            I => n14172
        );

    \I__11331\ : InMux
    port map (
            O => \N__50208\,
            I => \N__50205\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__50205\,
            I => n1696
        );

    \I__11329\ : InMux
    port map (
            O => \N__50202\,
            I => \N__50199\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__50199\,
            I => \N__50196\
        );

    \I__11327\ : Span4Mux_h
    port map (
            O => \N__50196\,
            I => \N__50192\
        );

    \I__11326\ : CascadeMux
    port map (
            O => \N__50195\,
            I => \N__50189\
        );

    \I__11325\ : Span4Mux_h
    port map (
            O => \N__50192\,
            I => \N__50183\
        );

    \I__11324\ : InMux
    port map (
            O => \N__50189\,
            I => \N__50176\
        );

    \I__11323\ : InMux
    port map (
            O => \N__50188\,
            I => \N__50176\
        );

    \I__11322\ : InMux
    port map (
            O => \N__50187\,
            I => \N__50176\
        );

    \I__11321\ : CascadeMux
    port map (
            O => \N__50186\,
            I => \N__50172\
        );

    \I__11320\ : Span4Mux_v
    port map (
            O => \N__50183\,
            I => \N__50160\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__50176\,
            I => \N__50160\
        );

    \I__11318\ : InMux
    port map (
            O => \N__50175\,
            I => \N__50153\
        );

    \I__11317\ : InMux
    port map (
            O => \N__50172\,
            I => \N__50153\
        );

    \I__11316\ : InMux
    port map (
            O => \N__50171\,
            I => \N__50153\
        );

    \I__11315\ : CascadeMux
    port map (
            O => \N__50170\,
            I => \N__50150\
        );

    \I__11314\ : CascadeMux
    port map (
            O => \N__50169\,
            I => \N__50147\
        );

    \I__11313\ : InMux
    port map (
            O => \N__50168\,
            I => \N__50137\
        );

    \I__11312\ : InMux
    port map (
            O => \N__50167\,
            I => \N__50137\
        );

    \I__11311\ : InMux
    port map (
            O => \N__50166\,
            I => \N__50137\
        );

    \I__11310\ : InMux
    port map (
            O => \N__50165\,
            I => \N__50134\
        );

    \I__11309\ : Span4Mux_v
    port map (
            O => \N__50160\,
            I => \N__50129\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__50153\,
            I => \N__50129\
        );

    \I__11307\ : InMux
    port map (
            O => \N__50150\,
            I => \N__50118\
        );

    \I__11306\ : InMux
    port map (
            O => \N__50147\,
            I => \N__50118\
        );

    \I__11305\ : InMux
    port map (
            O => \N__50146\,
            I => \N__50118\
        );

    \I__11304\ : InMux
    port map (
            O => \N__50145\,
            I => \N__50118\
        );

    \I__11303\ : InMux
    port map (
            O => \N__50144\,
            I => \N__50118\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__50137\,
            I => n1653
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__50134\,
            I => n1653
        );

    \I__11300\ : Odrv4
    port map (
            O => \N__50129\,
            I => n1653
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__50118\,
            I => n1653
        );

    \I__11298\ : CascadeMux
    port map (
            O => \N__50109\,
            I => \N__50106\
        );

    \I__11297\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50102\
        );

    \I__11296\ : CascadeMux
    port map (
            O => \N__50105\,
            I => \N__50099\
        );

    \I__11295\ : LocalMux
    port map (
            O => \N__50102\,
            I => \N__50096\
        );

    \I__11294\ : InMux
    port map (
            O => \N__50099\,
            I => \N__50093\
        );

    \I__11293\ : Span4Mux_v
    port map (
            O => \N__50096\,
            I => \N__50087\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__50093\,
            I => \N__50087\
        );

    \I__11291\ : InMux
    port map (
            O => \N__50092\,
            I => \N__50084\
        );

    \I__11290\ : Odrv4
    port map (
            O => \N__50087\,
            I => n1728
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__50084\,
            I => n1728
        );

    \I__11288\ : InMux
    port map (
            O => \N__50079\,
            I => \N__50076\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__50076\,
            I => \N__50073\
        );

    \I__11286\ : Odrv4
    port map (
            O => \N__50073\,
            I => n14508
        );

    \I__11285\ : CascadeMux
    port map (
            O => \N__50070\,
            I => \N__50067\
        );

    \I__11284\ : InMux
    port map (
            O => \N__50067\,
            I => \N__50064\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__50064\,
            I => \N__50061\
        );

    \I__11282\ : Span4Mux_h
    port map (
            O => \N__50061\,
            I => \N__50058\
        );

    \I__11281\ : Odrv4
    port map (
            O => \N__50058\,
            I => n1395
        );

    \I__11280\ : CascadeMux
    port map (
            O => \N__50055\,
            I => \n1427_cascade_\
        );

    \I__11279\ : CascadeMux
    port map (
            O => \N__50052\,
            I => \N__50048\
        );

    \I__11278\ : CascadeMux
    port map (
            O => \N__50051\,
            I => \N__50045\
        );

    \I__11277\ : InMux
    port map (
            O => \N__50048\,
            I => \N__50042\
        );

    \I__11276\ : InMux
    port map (
            O => \N__50045\,
            I => \N__50039\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__50042\,
            I => \N__50034\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__50039\,
            I => \N__50034\
        );

    \I__11273\ : Span4Mux_h
    port map (
            O => \N__50034\,
            I => \N__50031\
        );

    \I__11272\ : Odrv4
    port map (
            O => \N__50031\,
            I => n1526
        );

    \I__11271\ : CascadeMux
    port map (
            O => \N__50028\,
            I => \n1526_cascade_\
        );

    \I__11270\ : InMux
    port map (
            O => \N__50025\,
            I => \N__50022\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__50022\,
            I => \N__50019\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__50019\,
            I => \N__50016\
        );

    \I__11267\ : Odrv4
    port map (
            O => \N__50016\,
            I => n1593
        );

    \I__11266\ : CascadeMux
    port map (
            O => \N__50013\,
            I => \N__50009\
        );

    \I__11265\ : CascadeMux
    port map (
            O => \N__50012\,
            I => \N__50006\
        );

    \I__11264\ : InMux
    port map (
            O => \N__50009\,
            I => \N__50000\
        );

    \I__11263\ : InMux
    port map (
            O => \N__50006\,
            I => \N__50000\
        );

    \I__11262\ : InMux
    port map (
            O => \N__50005\,
            I => \N__49997\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__50000\,
            I => n1625_adj_612
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__49997\,
            I => n1625_adj_612
        );

    \I__11259\ : InMux
    port map (
            O => \N__49992\,
            I => \N__49988\
        );

    \I__11258\ : InMux
    port map (
            O => \N__49991\,
            I => \N__49984\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__49988\,
            I => \N__49981\
        );

    \I__11256\ : CascadeMux
    port map (
            O => \N__49987\,
            I => \N__49978\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__49984\,
            I => \N__49974\
        );

    \I__11254\ : Span4Mux_v
    port map (
            O => \N__49981\,
            I => \N__49971\
        );

    \I__11253\ : InMux
    port map (
            O => \N__49978\,
            I => \N__49968\
        );

    \I__11252\ : InMux
    port map (
            O => \N__49977\,
            I => \N__49965\
        );

    \I__11251\ : Odrv4
    port map (
            O => \N__49974\,
            I => n1528
        );

    \I__11250\ : Odrv4
    port map (
            O => \N__49971\,
            I => n1528
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__49968\,
            I => n1528
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__49965\,
            I => n1528
        );

    \I__11247\ : CascadeMux
    port map (
            O => \N__49956\,
            I => \N__49952\
        );

    \I__11246\ : CascadeMux
    port map (
            O => \N__49955\,
            I => \N__49949\
        );

    \I__11245\ : InMux
    port map (
            O => \N__49952\,
            I => \N__49946\
        );

    \I__11244\ : InMux
    port map (
            O => \N__49949\,
            I => \N__49943\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__49946\,
            I => \N__49940\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__49943\,
            I => \N__49937\
        );

    \I__11241\ : Span4Mux_h
    port map (
            O => \N__49940\,
            I => \N__49934\
        );

    \I__11240\ : Odrv4
    port map (
            O => \N__49937\,
            I => n1595
        );

    \I__11239\ : Odrv4
    port map (
            O => \N__49934\,
            I => n1595
        );

    \I__11238\ : CascadeMux
    port map (
            O => \N__49929\,
            I => \N__49925\
        );

    \I__11237\ : InMux
    port map (
            O => \N__49928\,
            I => \N__49922\
        );

    \I__11236\ : InMux
    port map (
            O => \N__49925\,
            I => \N__49919\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__49922\,
            I => n1627_adj_614
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__49919\,
            I => n1627_adj_614
        );

    \I__11233\ : InMux
    port map (
            O => \N__49914\,
            I => n12966
        );

    \I__11232\ : CascadeMux
    port map (
            O => \N__49911\,
            I => \N__49904\
        );

    \I__11231\ : CascadeMux
    port map (
            O => \N__49910\,
            I => \N__49900\
        );

    \I__11230\ : CascadeMux
    port map (
            O => \N__49909\,
            I => \N__49896\
        );

    \I__11229\ : InMux
    port map (
            O => \N__49908\,
            I => \N__49881\
        );

    \I__11228\ : InMux
    port map (
            O => \N__49907\,
            I => \N__49881\
        );

    \I__11227\ : InMux
    port map (
            O => \N__49904\,
            I => \N__49881\
        );

    \I__11226\ : InMux
    port map (
            O => \N__49903\,
            I => \N__49881\
        );

    \I__11225\ : InMux
    port map (
            O => \N__49900\,
            I => \N__49881\
        );

    \I__11224\ : InMux
    port map (
            O => \N__49899\,
            I => \N__49881\
        );

    \I__11223\ : InMux
    port map (
            O => \N__49896\,
            I => \N__49881\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__49881\,
            I => n11514
        );

    \I__11221\ : InMux
    port map (
            O => \N__49878\,
            I => \N__49875\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__49875\,
            I => n15089
        );

    \I__11219\ : InMux
    port map (
            O => \N__49872\,
            I => n12967
        );

    \I__11218\ : CascadeMux
    port map (
            O => \N__49869\,
            I => \N__49866\
        );

    \I__11217\ : InMux
    port map (
            O => \N__49866\,
            I => \N__49863\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__49863\,
            I => \N__49858\
        );

    \I__11215\ : InMux
    port map (
            O => \N__49862\,
            I => \N__49853\
        );

    \I__11214\ : InMux
    port map (
            O => \N__49861\,
            I => \N__49853\
        );

    \I__11213\ : Odrv4
    port map (
            O => \N__49858\,
            I => dti_counter_7
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__49853\,
            I => dti_counter_7
        );

    \I__11211\ : CascadeMux
    port map (
            O => \N__49848\,
            I => \n4_adj_716_cascade_\
        );

    \I__11210\ : CascadeMux
    port map (
            O => \N__49845\,
            I => \N__49842\
        );

    \I__11209\ : InMux
    port map (
            O => \N__49842\,
            I => \N__49837\
        );

    \I__11208\ : InMux
    port map (
            O => \N__49841\,
            I => \N__49834\
        );

    \I__11207\ : InMux
    port map (
            O => \N__49840\,
            I => \N__49831\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__49837\,
            I => dti_counter_6
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__49834\,
            I => dti_counter_6
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__49831\,
            I => dti_counter_6
        );

    \I__11203\ : InMux
    port map (
            O => \N__49824\,
            I => \N__49821\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__49821\,
            I => n15090
        );

    \I__11201\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49815\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__49815\,
            I => commutation_state_prev_1
        );

    \I__11199\ : InMux
    port map (
            O => \N__49812\,
            I => \N__49809\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__49809\,
            I => commutation_state_prev_2
        );

    \I__11197\ : InMux
    port map (
            O => \N__49806\,
            I => \N__49803\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__49803\,
            I => n1693_adj_621
        );

    \I__11195\ : InMux
    port map (
            O => \N__49800\,
            I => \N__49797\
        );

    \I__11194\ : LocalMux
    port map (
            O => \N__49797\,
            I => \N__49794\
        );

    \I__11193\ : Odrv4
    port map (
            O => \N__49794\,
            I => n1695
        );

    \I__11192\ : CascadeMux
    port map (
            O => \N__49791\,
            I => \N__49787\
        );

    \I__11191\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49784\
        );

    \I__11190\ : InMux
    port map (
            O => \N__49787\,
            I => \N__49781\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__49784\,
            I => \N__49776\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__49781\,
            I => \N__49776\
        );

    \I__11187\ : Odrv12
    port map (
            O => \N__49776\,
            I => n1727
        );

    \I__11186\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49770\
        );

    \I__11185\ : LocalMux
    port map (
            O => \N__49770\,
            I => \N__49767\
        );

    \I__11184\ : Odrv4
    port map (
            O => \N__49767\,
            I => n15088
        );

    \I__11183\ : InMux
    port map (
            O => \N__49764\,
            I => \N__49759\
        );

    \I__11182\ : InMux
    port map (
            O => \N__49763\,
            I => \N__49756\
        );

    \I__11181\ : InMux
    port map (
            O => \N__49762\,
            I => \N__49753\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__49759\,
            I => dti_counter_0
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__49756\,
            I => dti_counter_0
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__49753\,
            I => dti_counter_0
        );

    \I__11177\ : InMux
    port map (
            O => \N__49746\,
            I => \bfn_15_31_0_\
        );

    \I__11176\ : InMux
    port map (
            O => \N__49743\,
            I => \N__49740\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__49740\,
            I => n15095
        );

    \I__11174\ : InMux
    port map (
            O => \N__49737\,
            I => \N__49732\
        );

    \I__11173\ : InMux
    port map (
            O => \N__49736\,
            I => \N__49729\
        );

    \I__11172\ : InMux
    port map (
            O => \N__49735\,
            I => \N__49726\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__49732\,
            I => \N__49723\
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__49729\,
            I => \N__49720\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__49726\,
            I => dti_counter_1
        );

    \I__11168\ : Odrv4
    port map (
            O => \N__49723\,
            I => dti_counter_1
        );

    \I__11167\ : Odrv4
    port map (
            O => \N__49720\,
            I => dti_counter_1
        );

    \I__11166\ : InMux
    port map (
            O => \N__49713\,
            I => n12961
        );

    \I__11165\ : InMux
    port map (
            O => \N__49710\,
            I => \N__49707\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__49707\,
            I => n15094
        );

    \I__11163\ : CascadeMux
    port map (
            O => \N__49704\,
            I => \N__49700\
        );

    \I__11162\ : CascadeMux
    port map (
            O => \N__49703\,
            I => \N__49696\
        );

    \I__11161\ : InMux
    port map (
            O => \N__49700\,
            I => \N__49693\
        );

    \I__11160\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49690\
        );

    \I__11159\ : InMux
    port map (
            O => \N__49696\,
            I => \N__49687\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__49693\,
            I => \N__49682\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__49690\,
            I => \N__49682\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__49687\,
            I => dti_counter_2
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__49682\,
            I => dti_counter_2
        );

    \I__11154\ : InMux
    port map (
            O => \N__49677\,
            I => n12962
        );

    \I__11153\ : InMux
    port map (
            O => \N__49674\,
            I => \N__49671\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__49671\,
            I => n15093
        );

    \I__11151\ : InMux
    port map (
            O => \N__49668\,
            I => \N__49663\
        );

    \I__11150\ : InMux
    port map (
            O => \N__49667\,
            I => \N__49658\
        );

    \I__11149\ : InMux
    port map (
            O => \N__49666\,
            I => \N__49658\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__49663\,
            I => dti_counter_3
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__49658\,
            I => dti_counter_3
        );

    \I__11146\ : InMux
    port map (
            O => \N__49653\,
            I => n12963
        );

    \I__11145\ : InMux
    port map (
            O => \N__49650\,
            I => \N__49647\
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__49647\,
            I => n15092
        );

    \I__11143\ : CascadeMux
    port map (
            O => \N__49644\,
            I => \N__49640\
        );

    \I__11142\ : CascadeMux
    port map (
            O => \N__49643\,
            I => \N__49636\
        );

    \I__11141\ : InMux
    port map (
            O => \N__49640\,
            I => \N__49633\
        );

    \I__11140\ : InMux
    port map (
            O => \N__49639\,
            I => \N__49630\
        );

    \I__11139\ : InMux
    port map (
            O => \N__49636\,
            I => \N__49627\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__49633\,
            I => dti_counter_4
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__49630\,
            I => dti_counter_4
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__49627\,
            I => dti_counter_4
        );

    \I__11135\ : InMux
    port map (
            O => \N__49620\,
            I => n12964
        );

    \I__11134\ : InMux
    port map (
            O => \N__49617\,
            I => \N__49614\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__49614\,
            I => n15091
        );

    \I__11132\ : InMux
    port map (
            O => \N__49611\,
            I => \N__49606\
        );

    \I__11131\ : InMux
    port map (
            O => \N__49610\,
            I => \N__49603\
        );

    \I__11130\ : InMux
    port map (
            O => \N__49609\,
            I => \N__49600\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__49606\,
            I => dti_counter_5
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__49603\,
            I => dti_counter_5
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__49600\,
            I => dti_counter_5
        );

    \I__11126\ : InMux
    port map (
            O => \N__49593\,
            I => n12965
        );

    \I__11125\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49586\
        );

    \I__11124\ : CascadeMux
    port map (
            O => \N__49589\,
            I => \N__49582\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__49586\,
            I => \N__49578\
        );

    \I__11122\ : InMux
    port map (
            O => \N__49585\,
            I => \N__49575\
        );

    \I__11121\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49572\
        );

    \I__11120\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49569\
        );

    \I__11119\ : Span4Mux_v
    port map (
            O => \N__49578\,
            I => \N__49566\
        );

    \I__11118\ : LocalMux
    port map (
            O => \N__49575\,
            I => \N__49561\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__49572\,
            I => \N__49561\
        );

    \I__11116\ : LocalMux
    port map (
            O => \N__49569\,
            I => encoder0_position_target_20
        );

    \I__11115\ : Odrv4
    port map (
            O => \N__49566\,
            I => encoder0_position_target_20
        );

    \I__11114\ : Odrv4
    port map (
            O => \N__49561\,
            I => encoder0_position_target_20
        );

    \I__11113\ : InMux
    port map (
            O => \N__49554\,
            I => n12455
        );

    \I__11112\ : InMux
    port map (
            O => \N__49551\,
            I => n12456
        );

    \I__11111\ : CascadeMux
    port map (
            O => \N__49548\,
            I => \N__49544\
        );

    \I__11110\ : InMux
    port map (
            O => \N__49547\,
            I => \N__49541\
        );

    \I__11109\ : InMux
    port map (
            O => \N__49544\,
            I => \N__49538\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__49541\,
            I => \N__49534\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__49538\,
            I => \N__49530\
        );

    \I__11106\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49527\
        );

    \I__11105\ : Span4Mux_h
    port map (
            O => \N__49534\,
            I => \N__49524\
        );

    \I__11104\ : InMux
    port map (
            O => \N__49533\,
            I => \N__49521\
        );

    \I__11103\ : Span4Mux_h
    port map (
            O => \N__49530\,
            I => \N__49516\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__49527\,
            I => \N__49516\
        );

    \I__11101\ : Span4Mux_h
    port map (
            O => \N__49524\,
            I => \N__49513\
        );

    \I__11100\ : LocalMux
    port map (
            O => \N__49521\,
            I => encoder0_position_target_22
        );

    \I__11099\ : Odrv4
    port map (
            O => \N__49516\,
            I => encoder0_position_target_22
        );

    \I__11098\ : Odrv4
    port map (
            O => \N__49513\,
            I => encoder0_position_target_22
        );

    \I__11097\ : InMux
    port map (
            O => \N__49506\,
            I => n12457
        );

    \I__11096\ : InMux
    port map (
            O => \N__49503\,
            I => \bfn_15_28_0_\
        );

    \I__11095\ : CascadeMux
    port map (
            O => \N__49500\,
            I => \n14_adj_718_cascade_\
        );

    \I__11094\ : InMux
    port map (
            O => \N__49497\,
            I => \N__49494\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__49494\,
            I => n10_adj_719
        );

    \I__11092\ : CascadeMux
    port map (
            O => \N__49491\,
            I => \n5119_cascade_\
        );

    \I__11091\ : CascadeMux
    port map (
            O => \N__49488\,
            I => \N__49485\
        );

    \I__11090\ : InMux
    port map (
            O => \N__49485\,
            I => \N__49480\
        );

    \I__11089\ : InMux
    port map (
            O => \N__49484\,
            I => \N__49477\
        );

    \I__11088\ : CascadeMux
    port map (
            O => \N__49483\,
            I => \N__49474\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__49480\,
            I => \N__49471\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__49477\,
            I => \N__49467\
        );

    \I__11085\ : InMux
    port map (
            O => \N__49474\,
            I => \N__49464\
        );

    \I__11084\ : Span4Mux_v
    port map (
            O => \N__49471\,
            I => \N__49461\
        );

    \I__11083\ : InMux
    port map (
            O => \N__49470\,
            I => \N__49458\
        );

    \I__11082\ : Span4Mux_v
    port map (
            O => \N__49467\,
            I => \N__49455\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__49464\,
            I => encoder0_position_target_11
        );

    \I__11080\ : Odrv4
    port map (
            O => \N__49461\,
            I => encoder0_position_target_11
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__49458\,
            I => encoder0_position_target_11
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__49455\,
            I => encoder0_position_target_11
        );

    \I__11077\ : InMux
    port map (
            O => \N__49446\,
            I => n12446
        );

    \I__11076\ : CascadeMux
    port map (
            O => \N__49443\,
            I => \N__49439\
        );

    \I__11075\ : CascadeMux
    port map (
            O => \N__49442\,
            I => \N__49436\
        );

    \I__11074\ : InMux
    port map (
            O => \N__49439\,
            I => \N__49432\
        );

    \I__11073\ : InMux
    port map (
            O => \N__49436\,
            I => \N__49429\
        );

    \I__11072\ : InMux
    port map (
            O => \N__49435\,
            I => \N__49426\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__49432\,
            I => \N__49422\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__49429\,
            I => \N__49419\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__49426\,
            I => \N__49416\
        );

    \I__11068\ : InMux
    port map (
            O => \N__49425\,
            I => \N__49413\
        );

    \I__11067\ : Span4Mux_v
    port map (
            O => \N__49422\,
            I => \N__49410\
        );

    \I__11066\ : Span4Mux_h
    port map (
            O => \N__49419\,
            I => \N__49407\
        );

    \I__11065\ : Span4Mux_h
    port map (
            O => \N__49416\,
            I => \N__49404\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__49413\,
            I => encoder0_position_target_12
        );

    \I__11063\ : Odrv4
    port map (
            O => \N__49410\,
            I => encoder0_position_target_12
        );

    \I__11062\ : Odrv4
    port map (
            O => \N__49407\,
            I => encoder0_position_target_12
        );

    \I__11061\ : Odrv4
    port map (
            O => \N__49404\,
            I => encoder0_position_target_12
        );

    \I__11060\ : InMux
    port map (
            O => \N__49395\,
            I => n12447
        );

    \I__11059\ : CascadeMux
    port map (
            O => \N__49392\,
            I => \N__49389\
        );

    \I__11058\ : InMux
    port map (
            O => \N__49389\,
            I => \N__49384\
        );

    \I__11057\ : InMux
    port map (
            O => \N__49388\,
            I => \N__49381\
        );

    \I__11056\ : CascadeMux
    port map (
            O => \N__49387\,
            I => \N__49377\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__49384\,
            I => \N__49374\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__49381\,
            I => \N__49371\
        );

    \I__11053\ : InMux
    port map (
            O => \N__49380\,
            I => \N__49368\
        );

    \I__11052\ : InMux
    port map (
            O => \N__49377\,
            I => \N__49365\
        );

    \I__11051\ : Span4Mux_h
    port map (
            O => \N__49374\,
            I => \N__49362\
        );

    \I__11050\ : Span4Mux_h
    port map (
            O => \N__49371\,
            I => \N__49359\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__49368\,
            I => \N__49356\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__49365\,
            I => encoder0_position_target_13
        );

    \I__11047\ : Odrv4
    port map (
            O => \N__49362\,
            I => encoder0_position_target_13
        );

    \I__11046\ : Odrv4
    port map (
            O => \N__49359\,
            I => encoder0_position_target_13
        );

    \I__11045\ : Odrv12
    port map (
            O => \N__49356\,
            I => encoder0_position_target_13
        );

    \I__11044\ : InMux
    port map (
            O => \N__49347\,
            I => n12448
        );

    \I__11043\ : CascadeMux
    port map (
            O => \N__49344\,
            I => \N__49341\
        );

    \I__11042\ : InMux
    port map (
            O => \N__49341\,
            I => \N__49337\
        );

    \I__11041\ : InMux
    port map (
            O => \N__49340\,
            I => \N__49334\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__49337\,
            I => \N__49329\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__49334\,
            I => \N__49326\
        );

    \I__11038\ : CascadeMux
    port map (
            O => \N__49333\,
            I => \N__49323\
        );

    \I__11037\ : InMux
    port map (
            O => \N__49332\,
            I => \N__49320\
        );

    \I__11036\ : Span4Mux_h
    port map (
            O => \N__49329\,
            I => \N__49317\
        );

    \I__11035\ : Span4Mux_h
    port map (
            O => \N__49326\,
            I => \N__49314\
        );

    \I__11034\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49311\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__49320\,
            I => encoder0_position_target_14
        );

    \I__11032\ : Odrv4
    port map (
            O => \N__49317\,
            I => encoder0_position_target_14
        );

    \I__11031\ : Odrv4
    port map (
            O => \N__49314\,
            I => encoder0_position_target_14
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__49311\,
            I => encoder0_position_target_14
        );

    \I__11029\ : InMux
    port map (
            O => \N__49302\,
            I => n12449
        );

    \I__11028\ : InMux
    port map (
            O => \N__49299\,
            I => \bfn_15_27_0_\
        );

    \I__11027\ : CascadeMux
    port map (
            O => \N__49296\,
            I => \N__49293\
        );

    \I__11026\ : InMux
    port map (
            O => \N__49293\,
            I => \N__49290\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__49290\,
            I => \N__49285\
        );

    \I__11024\ : InMux
    port map (
            O => \N__49289\,
            I => \N__49282\
        );

    \I__11023\ : InMux
    port map (
            O => \N__49288\,
            I => \N__49278\
        );

    \I__11022\ : Span4Mux_h
    port map (
            O => \N__49285\,
            I => \N__49275\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__49282\,
            I => \N__49272\
        );

    \I__11020\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49269\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__49278\,
            I => encoder0_position_target_16
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__49275\,
            I => encoder0_position_target_16
        );

    \I__11017\ : Odrv4
    port map (
            O => \N__49272\,
            I => encoder0_position_target_16
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__49269\,
            I => encoder0_position_target_16
        );

    \I__11015\ : InMux
    port map (
            O => \N__49260\,
            I => n12451
        );

    \I__11014\ : CascadeMux
    port map (
            O => \N__49257\,
            I => \N__49254\
        );

    \I__11013\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49250\
        );

    \I__11012\ : CascadeMux
    port map (
            O => \N__49253\,
            I => \N__49246\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__49250\,
            I => \N__49243\
        );

    \I__11010\ : InMux
    port map (
            O => \N__49249\,
            I => \N__49239\
        );

    \I__11009\ : InMux
    port map (
            O => \N__49246\,
            I => \N__49236\
        );

    \I__11008\ : Span4Mux_h
    port map (
            O => \N__49243\,
            I => \N__49233\
        );

    \I__11007\ : InMux
    port map (
            O => \N__49242\,
            I => \N__49230\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__49239\,
            I => \N__49227\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__49236\,
            I => encoder0_position_target_17
        );

    \I__11004\ : Odrv4
    port map (
            O => \N__49233\,
            I => encoder0_position_target_17
        );

    \I__11003\ : LocalMux
    port map (
            O => \N__49230\,
            I => encoder0_position_target_17
        );

    \I__11002\ : Odrv4
    port map (
            O => \N__49227\,
            I => encoder0_position_target_17
        );

    \I__11001\ : InMux
    port map (
            O => \N__49218\,
            I => n12452
        );

    \I__11000\ : CascadeMux
    port map (
            O => \N__49215\,
            I => \N__49212\
        );

    \I__10999\ : InMux
    port map (
            O => \N__49212\,
            I => \N__49208\
        );

    \I__10998\ : InMux
    port map (
            O => \N__49211\,
            I => \N__49204\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__49208\,
            I => \N__49201\
        );

    \I__10996\ : InMux
    port map (
            O => \N__49207\,
            I => \N__49198\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__49204\,
            I => \N__49195\
        );

    \I__10994\ : Span4Mux_h
    port map (
            O => \N__49201\,
            I => \N__49191\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__49198\,
            I => \N__49186\
        );

    \I__10992\ : Span4Mux_v
    port map (
            O => \N__49195\,
            I => \N__49186\
        );

    \I__10991\ : InMux
    port map (
            O => \N__49194\,
            I => \N__49183\
        );

    \I__10990\ : Odrv4
    port map (
            O => \N__49191\,
            I => encoder0_position_target_18
        );

    \I__10989\ : Odrv4
    port map (
            O => \N__49186\,
            I => encoder0_position_target_18
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__49183\,
            I => encoder0_position_target_18
        );

    \I__10987\ : InMux
    port map (
            O => \N__49176\,
            I => n12453
        );

    \I__10986\ : InMux
    port map (
            O => \N__49173\,
            I => n12454
        );

    \I__10985\ : CascadeMux
    port map (
            O => \N__49170\,
            I => \N__49167\
        );

    \I__10984\ : InMux
    port map (
            O => \N__49167\,
            I => \N__49163\
        );

    \I__10983\ : CascadeMux
    port map (
            O => \N__49166\,
            I => \N__49160\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__49163\,
            I => \N__49157\
        );

    \I__10981\ : InMux
    port map (
            O => \N__49160\,
            I => \N__49153\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__49157\,
            I => \N__49150\
        );

    \I__10979\ : InMux
    port map (
            O => \N__49156\,
            I => \N__49147\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__49153\,
            I => encoder0_position_target_3
        );

    \I__10977\ : Odrv4
    port map (
            O => \N__49150\,
            I => encoder0_position_target_3
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__49147\,
            I => encoder0_position_target_3
        );

    \I__10975\ : InMux
    port map (
            O => \N__49140\,
            I => n12438
        );

    \I__10974\ : InMux
    port map (
            O => \N__49137\,
            I => \N__49133\
        );

    \I__10973\ : CascadeMux
    port map (
            O => \N__49136\,
            I => \N__49130\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__49133\,
            I => \N__49127\
        );

    \I__10971\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49122\
        );

    \I__10970\ : Span4Mux_v
    port map (
            O => \N__49127\,
            I => \N__49119\
        );

    \I__10969\ : InMux
    port map (
            O => \N__49126\,
            I => \N__49114\
        );

    \I__10968\ : InMux
    port map (
            O => \N__49125\,
            I => \N__49114\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__49122\,
            I => encoder0_position_target_4
        );

    \I__10966\ : Odrv4
    port map (
            O => \N__49119\,
            I => encoder0_position_target_4
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__49114\,
            I => encoder0_position_target_4
        );

    \I__10964\ : InMux
    port map (
            O => \N__49107\,
            I => n12439
        );

    \I__10963\ : CascadeMux
    port map (
            O => \N__49104\,
            I => \N__49101\
        );

    \I__10962\ : InMux
    port map (
            O => \N__49101\,
            I => \N__49097\
        );

    \I__10961\ : CascadeMux
    port map (
            O => \N__49100\,
            I => \N__49094\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__49097\,
            I => \N__49091\
        );

    \I__10959\ : InMux
    port map (
            O => \N__49094\,
            I => \N__49086\
        );

    \I__10958\ : Span4Mux_h
    port map (
            O => \N__49091\,
            I => \N__49083\
        );

    \I__10957\ : InMux
    port map (
            O => \N__49090\,
            I => \N__49078\
        );

    \I__10956\ : InMux
    port map (
            O => \N__49089\,
            I => \N__49078\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__49086\,
            I => encoder0_position_target_5
        );

    \I__10954\ : Odrv4
    port map (
            O => \N__49083\,
            I => encoder0_position_target_5
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__49078\,
            I => encoder0_position_target_5
        );

    \I__10952\ : InMux
    port map (
            O => \N__49071\,
            I => n12440
        );

    \I__10951\ : CascadeMux
    port map (
            O => \N__49068\,
            I => \N__49064\
        );

    \I__10950\ : CascadeMux
    port map (
            O => \N__49067\,
            I => \N__49061\
        );

    \I__10949\ : InMux
    port map (
            O => \N__49064\,
            I => \N__49058\
        );

    \I__10948\ : InMux
    port map (
            O => \N__49061\,
            I => \N__49053\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__49058\,
            I => \N__49050\
        );

    \I__10946\ : CascadeMux
    port map (
            O => \N__49057\,
            I => \N__49047\
        );

    \I__10945\ : CascadeMux
    port map (
            O => \N__49056\,
            I => \N__49044\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__49053\,
            I => \N__49039\
        );

    \I__10943\ : Span4Mux_h
    port map (
            O => \N__49050\,
            I => \N__49039\
        );

    \I__10942\ : InMux
    port map (
            O => \N__49047\,
            I => \N__49036\
        );

    \I__10941\ : InMux
    port map (
            O => \N__49044\,
            I => \N__49033\
        );

    \I__10940\ : Span4Mux_h
    port map (
            O => \N__49039\,
            I => \N__49030\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__49036\,
            I => encoder0_position_target_6
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__49033\,
            I => encoder0_position_target_6
        );

    \I__10937\ : Odrv4
    port map (
            O => \N__49030\,
            I => encoder0_position_target_6
        );

    \I__10936\ : InMux
    port map (
            O => \N__49023\,
            I => n12441
        );

    \I__10935\ : InMux
    port map (
            O => \N__49020\,
            I => \N__49015\
        );

    \I__10934\ : InMux
    port map (
            O => \N__49019\,
            I => \N__49012\
        );

    \I__10933\ : CascadeMux
    port map (
            O => \N__49018\,
            I => \N__49009\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__49015\,
            I => \N__49003\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__49012\,
            I => \N__49003\
        );

    \I__10930\ : InMux
    port map (
            O => \N__49009\,
            I => \N__49000\
        );

    \I__10929\ : InMux
    port map (
            O => \N__49008\,
            I => \N__48997\
        );

    \I__10928\ : Span4Mux_h
    port map (
            O => \N__49003\,
            I => \N__48994\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__49000\,
            I => encoder0_position_target_7
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__48997\,
            I => encoder0_position_target_7
        );

    \I__10925\ : Odrv4
    port map (
            O => \N__48994\,
            I => encoder0_position_target_7
        );

    \I__10924\ : InMux
    port map (
            O => \N__48987\,
            I => \bfn_15_26_0_\
        );

    \I__10923\ : CascadeMux
    port map (
            O => \N__48984\,
            I => \N__48981\
        );

    \I__10922\ : InMux
    port map (
            O => \N__48981\,
            I => \N__48978\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__48978\,
            I => \N__48973\
        );

    \I__10920\ : InMux
    port map (
            O => \N__48977\,
            I => \N__48969\
        );

    \I__10919\ : InMux
    port map (
            O => \N__48976\,
            I => \N__48966\
        );

    \I__10918\ : Span4Mux_h
    port map (
            O => \N__48973\,
            I => \N__48963\
        );

    \I__10917\ : InMux
    port map (
            O => \N__48972\,
            I => \N__48960\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__48969\,
            I => \N__48957\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__48966\,
            I => encoder0_position_target_8
        );

    \I__10914\ : Odrv4
    port map (
            O => \N__48963\,
            I => encoder0_position_target_8
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__48960\,
            I => encoder0_position_target_8
        );

    \I__10912\ : Odrv12
    port map (
            O => \N__48957\,
            I => encoder0_position_target_8
        );

    \I__10911\ : InMux
    port map (
            O => \N__48948\,
            I => n12443
        );

    \I__10910\ : CascadeMux
    port map (
            O => \N__48945\,
            I => \N__48942\
        );

    \I__10909\ : InMux
    port map (
            O => \N__48942\,
            I => \N__48937\
        );

    \I__10908\ : CascadeMux
    port map (
            O => \N__48941\,
            I => \N__48934\
        );

    \I__10907\ : InMux
    port map (
            O => \N__48940\,
            I => \N__48931\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48928\
        );

    \I__10905\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48924\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__48931\,
            I => \N__48921\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__48928\,
            I => \N__48918\
        );

    \I__10902\ : InMux
    port map (
            O => \N__48927\,
            I => \N__48915\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__48924\,
            I => \N__48910\
        );

    \I__10900\ : Span4Mux_h
    port map (
            O => \N__48921\,
            I => \N__48910\
        );

    \I__10899\ : Odrv4
    port map (
            O => \N__48918\,
            I => encoder0_position_target_9
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__48915\,
            I => encoder0_position_target_9
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__48910\,
            I => encoder0_position_target_9
        );

    \I__10896\ : InMux
    port map (
            O => \N__48903\,
            I => n12444
        );

    \I__10895\ : CascadeMux
    port map (
            O => \N__48900\,
            I => \N__48897\
        );

    \I__10894\ : InMux
    port map (
            O => \N__48897\,
            I => \N__48893\
        );

    \I__10893\ : InMux
    port map (
            O => \N__48896\,
            I => \N__48890\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__48893\,
            I => \N__48885\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__48890\,
            I => \N__48882\
        );

    \I__10890\ : InMux
    port map (
            O => \N__48889\,
            I => \N__48879\
        );

    \I__10889\ : InMux
    port map (
            O => \N__48888\,
            I => \N__48876\
        );

    \I__10888\ : Span4Mux_v
    port map (
            O => \N__48885\,
            I => \N__48871\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__48882\,
            I => \N__48871\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__48879\,
            I => encoder0_position_target_10
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__48876\,
            I => encoder0_position_target_10
        );

    \I__10884\ : Odrv4
    port map (
            O => \N__48871\,
            I => encoder0_position_target_10
        );

    \I__10883\ : InMux
    port map (
            O => \N__48864\,
            I => n12445
        );

    \I__10882\ : InMux
    port map (
            O => \N__48861\,
            I => n12523
        );

    \I__10881\ : InMux
    port map (
            O => \N__48858\,
            I => \bfn_15_24_0_\
        );

    \I__10880\ : InMux
    port map (
            O => \N__48855\,
            I => \N__48852\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__48852\,
            I => \N__48849\
        );

    \I__10878\ : Odrv4
    port map (
            O => \N__48849\,
            I => n1292
        );

    \I__10877\ : InMux
    port map (
            O => \N__48846\,
            I => n12525
        );

    \I__10876\ : InMux
    port map (
            O => \N__48843\,
            I => n12526
        );

    \I__10875\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48836\
        );

    \I__10874\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48833\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__48836\,
            I => \N__48828\
        );

    \I__10872\ : LocalMux
    port map (
            O => \N__48833\,
            I => \N__48828\
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__48828\,
            I => n1323
        );

    \I__10870\ : CascadeMux
    port map (
            O => \N__48825\,
            I => \N__48822\
        );

    \I__10869\ : InMux
    port map (
            O => \N__48822\,
            I => \N__48819\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__48819\,
            I => \N__48816\
        );

    \I__10867\ : Span4Mux_h
    port map (
            O => \N__48816\,
            I => \N__48812\
        );

    \I__10866\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48808\
        );

    \I__10865\ : Span4Mux_h
    port map (
            O => \N__48812\,
            I => \N__48805\
        );

    \I__10864\ : InMux
    port map (
            O => \N__48811\,
            I => \N__48802\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__48808\,
            I => encoder0_position_target_0
        );

    \I__10862\ : Odrv4
    port map (
            O => \N__48805\,
            I => encoder0_position_target_0
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__48802\,
            I => encoder0_position_target_0
        );

    \I__10860\ : InMux
    port map (
            O => \N__48795\,
            I => n12435
        );

    \I__10859\ : CascadeMux
    port map (
            O => \N__48792\,
            I => \N__48789\
        );

    \I__10858\ : InMux
    port map (
            O => \N__48789\,
            I => \N__48785\
        );

    \I__10857\ : CascadeMux
    port map (
            O => \N__48788\,
            I => \N__48781\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__48785\,
            I => \N__48778\
        );

    \I__10855\ : CascadeMux
    port map (
            O => \N__48784\,
            I => \N__48775\
        );

    \I__10854\ : InMux
    port map (
            O => \N__48781\,
            I => \N__48772\
        );

    \I__10853\ : Span4Mux_h
    port map (
            O => \N__48778\,
            I => \N__48769\
        );

    \I__10852\ : InMux
    port map (
            O => \N__48775\,
            I => \N__48766\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__48772\,
            I => encoder0_position_target_1
        );

    \I__10850\ : Odrv4
    port map (
            O => \N__48769\,
            I => encoder0_position_target_1
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__48766\,
            I => encoder0_position_target_1
        );

    \I__10848\ : InMux
    port map (
            O => \N__48759\,
            I => n12436
        );

    \I__10847\ : InMux
    port map (
            O => \N__48756\,
            I => \N__48752\
        );

    \I__10846\ : CascadeMux
    port map (
            O => \N__48755\,
            I => \N__48749\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__48752\,
            I => \N__48746\
        );

    \I__10844\ : InMux
    port map (
            O => \N__48749\,
            I => \N__48742\
        );

    \I__10843\ : Span4Mux_h
    port map (
            O => \N__48746\,
            I => \N__48739\
        );

    \I__10842\ : InMux
    port map (
            O => \N__48745\,
            I => \N__48736\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__48742\,
            I => encoder0_position_target_2
        );

    \I__10840\ : Odrv4
    port map (
            O => \N__48739\,
            I => encoder0_position_target_2
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__48736\,
            I => encoder0_position_target_2
        );

    \I__10838\ : InMux
    port map (
            O => \N__48729\,
            I => n12437
        );

    \I__10837\ : CascadeMux
    port map (
            O => \N__48726\,
            I => \N__48722\
        );

    \I__10836\ : InMux
    port map (
            O => \N__48725\,
            I => \N__48718\
        );

    \I__10835\ : InMux
    port map (
            O => \N__48722\,
            I => \N__48715\
        );

    \I__10834\ : InMux
    port map (
            O => \N__48721\,
            I => \N__48712\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__48718\,
            I => n1329
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__48715\,
            I => n1329
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__48712\,
            I => n1329
        );

    \I__10830\ : CascadeMux
    port map (
            O => \N__48705\,
            I => \N__48700\
        );

    \I__10829\ : InMux
    port map (
            O => \N__48704\,
            I => \N__48695\
        );

    \I__10828\ : InMux
    port map (
            O => \N__48703\,
            I => \N__48695\
        );

    \I__10827\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48692\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__48695\,
            I => n1333
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__48692\,
            I => n1333
        );

    \I__10824\ : InMux
    port map (
            O => \N__48687\,
            I => \N__48682\
        );

    \I__10823\ : InMux
    port map (
            O => \N__48686\,
            I => \N__48679\
        );

    \I__10822\ : InMux
    port map (
            O => \N__48685\,
            I => \N__48676\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__48682\,
            I => n298
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__48679\,
            I => n298
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__48676\,
            I => n298
        );

    \I__10818\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48666\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__48666\,
            I => n1301
        );

    \I__10816\ : InMux
    port map (
            O => \N__48663\,
            I => \bfn_15_23_0_\
        );

    \I__10815\ : CascadeMux
    port map (
            O => \N__48660\,
            I => \N__48656\
        );

    \I__10814\ : InMux
    port map (
            O => \N__48659\,
            I => \N__48652\
        );

    \I__10813\ : InMux
    port map (
            O => \N__48656\,
            I => \N__48649\
        );

    \I__10812\ : InMux
    port map (
            O => \N__48655\,
            I => \N__48646\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__48652\,
            I => n1233
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__48649\,
            I => n1233
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__48646\,
            I => n1233
        );

    \I__10808\ : CascadeMux
    port map (
            O => \N__48639\,
            I => \N__48636\
        );

    \I__10807\ : InMux
    port map (
            O => \N__48636\,
            I => \N__48633\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__48633\,
            I => n1300
        );

    \I__10805\ : InMux
    port map (
            O => \N__48630\,
            I => n12517
        );

    \I__10804\ : CascadeMux
    port map (
            O => \N__48627\,
            I => \N__48624\
        );

    \I__10803\ : InMux
    port map (
            O => \N__48624\,
            I => \N__48620\
        );

    \I__10802\ : CascadeMux
    port map (
            O => \N__48623\,
            I => \N__48617\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__48620\,
            I => \N__48614\
        );

    \I__10800\ : InMux
    port map (
            O => \N__48617\,
            I => \N__48611\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__48614\,
            I => n1232
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__48611\,
            I => n1232
        );

    \I__10797\ : InMux
    port map (
            O => \N__48606\,
            I => \N__48603\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__48603\,
            I => \N__48600\
        );

    \I__10795\ : Span4Mux_v
    port map (
            O => \N__48600\,
            I => \N__48597\
        );

    \I__10794\ : Odrv4
    port map (
            O => \N__48597\,
            I => n1299
        );

    \I__10793\ : InMux
    port map (
            O => \N__48594\,
            I => n12518
        );

    \I__10792\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48588\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__48588\,
            I => \N__48585\
        );

    \I__10790\ : Odrv4
    port map (
            O => \N__48585\,
            I => n1298
        );

    \I__10789\ : InMux
    port map (
            O => \N__48582\,
            I => n12519
        );

    \I__10788\ : InMux
    port map (
            O => \N__48579\,
            I => \N__48576\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__48576\,
            I => n1297
        );

    \I__10786\ : InMux
    port map (
            O => \N__48573\,
            I => n12520
        );

    \I__10785\ : InMux
    port map (
            O => \N__48570\,
            I => n12521
        );

    \I__10784\ : InMux
    port map (
            O => \N__48567\,
            I => n12522
        );

    \I__10783\ : InMux
    port map (
            O => \N__48564\,
            I => n12532
        );

    \I__10782\ : InMux
    port map (
            O => \N__48561\,
            I => \N__48558\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__48558\,
            I => n1394
        );

    \I__10780\ : InMux
    port map (
            O => \N__48555\,
            I => n12533
        );

    \I__10779\ : InMux
    port map (
            O => \N__48552\,
            I => \N__48549\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__48549\,
            I => \N__48546\
        );

    \I__10777\ : Odrv12
    port map (
            O => \N__48546\,
            I => n1393
        );

    \I__10776\ : InMux
    port map (
            O => \N__48543\,
            I => \bfn_15_22_0_\
        );

    \I__10775\ : InMux
    port map (
            O => \N__48540\,
            I => n12535
        );

    \I__10774\ : CascadeMux
    port map (
            O => \N__48537\,
            I => \N__48534\
        );

    \I__10773\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48530\
        );

    \I__10772\ : InMux
    port map (
            O => \N__48533\,
            I => \N__48527\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__48530\,
            I => n1324
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__48527\,
            I => n1324
        );

    \I__10769\ : InMux
    port map (
            O => \N__48522\,
            I => \N__48519\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__48519\,
            I => n1391
        );

    \I__10767\ : InMux
    port map (
            O => \N__48516\,
            I => n12536
        );

    \I__10766\ : InMux
    port map (
            O => \N__48513\,
            I => \N__48510\
        );

    \I__10765\ : LocalMux
    port map (
            O => \N__48510\,
            I => \N__48507\
        );

    \I__10764\ : Span4Mux_h
    port map (
            O => \N__48507\,
            I => \N__48503\
        );

    \I__10763\ : CascadeMux
    port map (
            O => \N__48506\,
            I => \N__48500\
        );

    \I__10762\ : Span4Mux_h
    port map (
            O => \N__48503\,
            I => \N__48497\
        );

    \I__10761\ : InMux
    port map (
            O => \N__48500\,
            I => \N__48494\
        );

    \I__10760\ : Odrv4
    port map (
            O => \N__48497\,
            I => n15544
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__48494\,
            I => n15544
        );

    \I__10758\ : InMux
    port map (
            O => \N__48489\,
            I => n12537
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__48486\,
            I => \N__48483\
        );

    \I__10756\ : InMux
    port map (
            O => \N__48483\,
            I => \N__48478\
        );

    \I__10755\ : CascadeMux
    port map (
            O => \N__48482\,
            I => \N__48475\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__48481\,
            I => \N__48472\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__48478\,
            I => \N__48469\
        );

    \I__10752\ : InMux
    port map (
            O => \N__48475\,
            I => \N__48466\
        );

    \I__10751\ : InMux
    port map (
            O => \N__48472\,
            I => \N__48463\
        );

    \I__10750\ : Odrv4
    port map (
            O => \N__48469\,
            I => n1332
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__48466\,
            I => n1332
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__48463\,
            I => n1332
        );

    \I__10747\ : InMux
    port map (
            O => \N__48456\,
            I => \N__48453\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__48453\,
            I => n13727
        );

    \I__10745\ : CascadeMux
    port map (
            O => \N__48450\,
            I => \n14496_cascade_\
        );

    \I__10744\ : CascadeMux
    port map (
            O => \N__48447\,
            I => \n1455_cascade_\
        );

    \I__10743\ : CascadeMux
    port map (
            O => \N__48444\,
            I => \N__48441\
        );

    \I__10742\ : InMux
    port map (
            O => \N__48441\,
            I => \N__48437\
        );

    \I__10741\ : InMux
    port map (
            O => \N__48440\,
            I => \N__48433\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__48437\,
            I => \N__48430\
        );

    \I__10739\ : InMux
    port map (
            O => \N__48436\,
            I => \N__48427\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__48433\,
            I => n1525
        );

    \I__10737\ : Odrv4
    port map (
            O => \N__48430\,
            I => n1525
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__48427\,
            I => n1525
        );

    \I__10735\ : CascadeMux
    port map (
            O => \N__48420\,
            I => \N__48417\
        );

    \I__10734\ : InMux
    port map (
            O => \N__48417\,
            I => \N__48413\
        );

    \I__10733\ : InMux
    port map (
            O => \N__48416\,
            I => \N__48410\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__48413\,
            I => \N__48406\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__48410\,
            I => \N__48403\
        );

    \I__10730\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48400\
        );

    \I__10729\ : Odrv4
    port map (
            O => \N__48406\,
            I => n1524
        );

    \I__10728\ : Odrv4
    port map (
            O => \N__48403\,
            I => n1524
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__48400\,
            I => n1524
        );

    \I__10726\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48388\
        );

    \I__10725\ : InMux
    port map (
            O => \N__48392\,
            I => \N__48383\
        );

    \I__10724\ : InMux
    port map (
            O => \N__48391\,
            I => \N__48383\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__48388\,
            I => \N__48380\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__48383\,
            I => n299
        );

    \I__10721\ : Odrv4
    port map (
            O => \N__48380\,
            I => n299
        );

    \I__10720\ : CascadeMux
    port map (
            O => \N__48375\,
            I => \N__48372\
        );

    \I__10719\ : InMux
    port map (
            O => \N__48372\,
            I => \N__48369\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__48369\,
            I => n1401
        );

    \I__10717\ : InMux
    port map (
            O => \N__48366\,
            I => \bfn_15_21_0_\
        );

    \I__10716\ : InMux
    port map (
            O => \N__48363\,
            I => \N__48360\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__48360\,
            I => n1400
        );

    \I__10714\ : InMux
    port map (
            O => \N__48357\,
            I => n12527
        );

    \I__10713\ : InMux
    port map (
            O => \N__48354\,
            I => \N__48351\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__48351\,
            I => \N__48348\
        );

    \I__10711\ : Odrv4
    port map (
            O => \N__48348\,
            I => n1399
        );

    \I__10710\ : InMux
    port map (
            O => \N__48345\,
            I => n12528
        );

    \I__10709\ : CascadeMux
    port map (
            O => \N__48342\,
            I => \N__48338\
        );

    \I__10708\ : CascadeMux
    port map (
            O => \N__48341\,
            I => \N__48335\
        );

    \I__10707\ : InMux
    port map (
            O => \N__48338\,
            I => \N__48331\
        );

    \I__10706\ : InMux
    port map (
            O => \N__48335\,
            I => \N__48328\
        );

    \I__10705\ : InMux
    port map (
            O => \N__48334\,
            I => \N__48325\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__48331\,
            I => \N__48322\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__48328\,
            I => n1331
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__48325\,
            I => n1331
        );

    \I__10701\ : Odrv4
    port map (
            O => \N__48322\,
            I => n1331
        );

    \I__10700\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48312\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__48312\,
            I => n1398
        );

    \I__10698\ : InMux
    port map (
            O => \N__48309\,
            I => n12529
        );

    \I__10697\ : CascadeMux
    port map (
            O => \N__48306\,
            I => \N__48301\
        );

    \I__10696\ : InMux
    port map (
            O => \N__48305\,
            I => \N__48298\
        );

    \I__10695\ : InMux
    port map (
            O => \N__48304\,
            I => \N__48295\
        );

    \I__10694\ : InMux
    port map (
            O => \N__48301\,
            I => \N__48292\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__48298\,
            I => n1330
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__48295\,
            I => n1330
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__48292\,
            I => n1330
        );

    \I__10690\ : CascadeMux
    port map (
            O => \N__48285\,
            I => \N__48282\
        );

    \I__10689\ : InMux
    port map (
            O => \N__48282\,
            I => \N__48279\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__48279\,
            I => n1397
        );

    \I__10687\ : InMux
    port map (
            O => \N__48276\,
            I => n12530
        );

    \I__10686\ : InMux
    port map (
            O => \N__48273\,
            I => \N__48270\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__48270\,
            I => n1396
        );

    \I__10684\ : InMux
    port map (
            O => \N__48267\,
            I => n12531
        );

    \I__10683\ : InMux
    port map (
            O => \N__48264\,
            I => \N__48259\
        );

    \I__10682\ : InMux
    port map (
            O => \N__48263\,
            I => \N__48256\
        );

    \I__10681\ : InMux
    port map (
            O => \N__48262\,
            I => \N__48253\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__48259\,
            I => n1522
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__48256\,
            I => n1522
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__48253\,
            I => n1522
        );

    \I__10677\ : CascadeMux
    port map (
            O => \N__48246\,
            I => \n1523_cascade_\
        );

    \I__10676\ : InMux
    port map (
            O => \N__48243\,
            I => \N__48240\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__48240\,
            I => n14296
        );

    \I__10674\ : InMux
    port map (
            O => \N__48237\,
            I => \N__48234\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__48234\,
            I => \N__48231\
        );

    \I__10672\ : Odrv12
    port map (
            O => \N__48231\,
            I => n1601
        );

    \I__10671\ : CascadeMux
    port map (
            O => \N__48228\,
            I => \n1554_cascade_\
        );

    \I__10670\ : InMux
    port map (
            O => \N__48225\,
            I => \N__48220\
        );

    \I__10669\ : InMux
    port map (
            O => \N__48224\,
            I => \N__48217\
        );

    \I__10668\ : CascadeMux
    port map (
            O => \N__48223\,
            I => \N__48214\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__48220\,
            I => \N__48211\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__48217\,
            I => \N__48208\
        );

    \I__10665\ : InMux
    port map (
            O => \N__48214\,
            I => \N__48205\
        );

    \I__10664\ : Span4Mux_h
    port map (
            O => \N__48211\,
            I => \N__48200\
        );

    \I__10663\ : Span4Mux_h
    port map (
            O => \N__48208\,
            I => \N__48200\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__48205\,
            I => \N__48197\
        );

    \I__10661\ : Odrv4
    port map (
            O => \N__48200\,
            I => n301
        );

    \I__10660\ : Odrv4
    port map (
            O => \N__48197\,
            I => n301
        );

    \I__10659\ : CascadeMux
    port map (
            O => \N__48192\,
            I => \N__48189\
        );

    \I__10658\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48185\
        );

    \I__10657\ : CascadeMux
    port map (
            O => \N__48188\,
            I => \N__48182\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__48185\,
            I => \N__48178\
        );

    \I__10655\ : InMux
    port map (
            O => \N__48182\,
            I => \N__48173\
        );

    \I__10654\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48173\
        );

    \I__10653\ : Odrv4
    port map (
            O => \N__48178\,
            I => n1633_adj_620
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__48173\,
            I => n1633_adj_620
        );

    \I__10651\ : CascadeMux
    port map (
            O => \N__48168\,
            I => \N__48164\
        );

    \I__10650\ : CascadeMux
    port map (
            O => \N__48167\,
            I => \N__48161\
        );

    \I__10649\ : InMux
    port map (
            O => \N__48164\,
            I => \N__48157\
        );

    \I__10648\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48154\
        );

    \I__10647\ : InMux
    port map (
            O => \N__48160\,
            I => \N__48151\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__48157\,
            I => \N__48148\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__48154\,
            I => n1532
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__48151\,
            I => n1532
        );

    \I__10643\ : Odrv4
    port map (
            O => \N__48148\,
            I => n1532
        );

    \I__10642\ : CascadeMux
    port map (
            O => \N__48141\,
            I => \N__48138\
        );

    \I__10641\ : InMux
    port map (
            O => \N__48138\,
            I => \N__48135\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__48135\,
            I => \N__48132\
        );

    \I__10639\ : Odrv4
    port map (
            O => \N__48132\,
            I => n11906
        );

    \I__10638\ : CascadeMux
    port map (
            O => \N__48129\,
            I => \n14490_cascade_\
        );

    \I__10637\ : CascadeMux
    port map (
            O => \N__48126\,
            I => \N__48122\
        );

    \I__10636\ : CascadeMux
    port map (
            O => \N__48125\,
            I => \N__48119\
        );

    \I__10635\ : InMux
    port map (
            O => \N__48122\,
            I => \N__48116\
        );

    \I__10634\ : InMux
    port map (
            O => \N__48119\,
            I => \N__48113\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__48116\,
            I => \N__48109\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__48113\,
            I => \N__48106\
        );

    \I__10631\ : InMux
    port map (
            O => \N__48112\,
            I => \N__48103\
        );

    \I__10630\ : Span4Mux_h
    port map (
            O => \N__48109\,
            I => \N__48100\
        );

    \I__10629\ : Span4Mux_h
    port map (
            O => \N__48106\,
            I => \N__48097\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__48103\,
            I => n1623_adj_610
        );

    \I__10627\ : Odrv4
    port map (
            O => \N__48100\,
            I => n1623_adj_610
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__48097\,
            I => n1623_adj_610
        );

    \I__10625\ : CascadeMux
    port map (
            O => \N__48090\,
            I => \N__48087\
        );

    \I__10624\ : InMux
    port map (
            O => \N__48087\,
            I => \N__48084\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__48084\,
            I => \N__48081\
        );

    \I__10622\ : Span4Mux_v
    port map (
            O => \N__48081\,
            I => \N__48078\
        );

    \I__10621\ : Odrv4
    port map (
            O => \N__48078\,
            I => n1690
        );

    \I__10620\ : InMux
    port map (
            O => \N__48075\,
            I => n12573
        );

    \I__10619\ : InMux
    port map (
            O => \N__48072\,
            I => \N__48067\
        );

    \I__10618\ : CascadeMux
    port map (
            O => \N__48071\,
            I => \N__48064\
        );

    \I__10617\ : InMux
    port map (
            O => \N__48070\,
            I => \N__48061\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__48067\,
            I => \N__48058\
        );

    \I__10615\ : InMux
    port map (
            O => \N__48064\,
            I => \N__48055\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__48061\,
            I => \N__48052\
        );

    \I__10613\ : Odrv4
    port map (
            O => \N__48058\,
            I => n1622_adj_609
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__48055\,
            I => n1622_adj_609
        );

    \I__10611\ : Odrv4
    port map (
            O => \N__48052\,
            I => n1622_adj_609
        );

    \I__10610\ : CascadeMux
    port map (
            O => \N__48045\,
            I => \N__48042\
        );

    \I__10609\ : InMux
    port map (
            O => \N__48042\,
            I => \N__48039\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__48039\,
            I => \N__48036\
        );

    \I__10607\ : Span4Mux_v
    port map (
            O => \N__48036\,
            I => \N__48033\
        );

    \I__10606\ : Odrv4
    port map (
            O => \N__48033\,
            I => n1689
        );

    \I__10605\ : InMux
    port map (
            O => \N__48030\,
            I => n12574
        );

    \I__10604\ : InMux
    port map (
            O => \N__48027\,
            I => \N__48023\
        );

    \I__10603\ : InMux
    port map (
            O => \N__48026\,
            I => \N__48019\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__48023\,
            I => \N__48016\
        );

    \I__10601\ : InMux
    port map (
            O => \N__48022\,
            I => \N__48013\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__48019\,
            I => \N__48010\
        );

    \I__10599\ : Odrv4
    port map (
            O => \N__48016\,
            I => n1621_adj_608
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__48013\,
            I => n1621_adj_608
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__48010\,
            I => n1621_adj_608
        );

    \I__10596\ : InMux
    port map (
            O => \N__48003\,
            I => \N__48000\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__48000\,
            I => \N__47997\
        );

    \I__10594\ : Span4Mux_v
    port map (
            O => \N__47997\,
            I => \N__47994\
        );

    \I__10593\ : Odrv4
    port map (
            O => \N__47994\,
            I => n1688
        );

    \I__10592\ : InMux
    port map (
            O => \N__47991\,
            I => n12575
        );

    \I__10591\ : InMux
    port map (
            O => \N__47988\,
            I => \N__47985\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__47985\,
            I => \N__47982\
        );

    \I__10589\ : Span12Mux_h
    port map (
            O => \N__47982\,
            I => \N__47978\
        );

    \I__10588\ : InMux
    port map (
            O => \N__47981\,
            I => \N__47975\
        );

    \I__10587\ : Odrv12
    port map (
            O => \N__47978\,
            I => n15603
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__47975\,
            I => n15603
        );

    \I__10585\ : CascadeMux
    port map (
            O => \N__47970\,
            I => \N__47967\
        );

    \I__10584\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47964\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__47964\,
            I => \N__47960\
        );

    \I__10582\ : InMux
    port map (
            O => \N__47963\,
            I => \N__47957\
        );

    \I__10581\ : Span4Mux_h
    port map (
            O => \N__47960\,
            I => \N__47954\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__47957\,
            I => \N__47951\
        );

    \I__10579\ : Odrv4
    port map (
            O => \N__47954\,
            I => n1620_adj_607
        );

    \I__10578\ : Odrv4
    port map (
            O => \N__47951\,
            I => n1620_adj_607
        );

    \I__10577\ : InMux
    port map (
            O => \N__47946\,
            I => n12576
        );

    \I__10576\ : CascadeMux
    port map (
            O => \N__47943\,
            I => \N__47939\
        );

    \I__10575\ : InMux
    port map (
            O => \N__47942\,
            I => \N__47936\
        );

    \I__10574\ : InMux
    port map (
            O => \N__47939\,
            I => \N__47933\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__47936\,
            I => \N__47930\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__47933\,
            I => \N__47925\
        );

    \I__10571\ : Span4Mux_v
    port map (
            O => \N__47930\,
            I => \N__47925\
        );

    \I__10570\ : Odrv4
    port map (
            O => \N__47925\,
            I => n1719
        );

    \I__10569\ : InMux
    port map (
            O => \N__47922\,
            I => \N__47919\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__47919\,
            I => n1692
        );

    \I__10567\ : CascadeMux
    port map (
            O => \N__47916\,
            I => \N__47913\
        );

    \I__10566\ : InMux
    port map (
            O => \N__47913\,
            I => \N__47910\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__47910\,
            I => \N__47906\
        );

    \I__10564\ : InMux
    port map (
            O => \N__47909\,
            I => \N__47903\
        );

    \I__10563\ : Span4Mux_h
    port map (
            O => \N__47906\,
            I => \N__47900\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__47903\,
            I => n1523
        );

    \I__10561\ : Odrv4
    port map (
            O => \N__47900\,
            I => n1523
        );

    \I__10560\ : CascadeMux
    port map (
            O => \N__47895\,
            I => \N__47892\
        );

    \I__10559\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47888\
        );

    \I__10558\ : CascadeMux
    port map (
            O => \N__47891\,
            I => \N__47885\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__47888\,
            I => \N__47881\
        );

    \I__10556\ : InMux
    port map (
            O => \N__47885\,
            I => \N__47876\
        );

    \I__10555\ : InMux
    port map (
            O => \N__47884\,
            I => \N__47876\
        );

    \I__10554\ : Odrv4
    port map (
            O => \N__47881\,
            I => n1632_adj_619
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__47876\,
            I => n1632_adj_619
        );

    \I__10552\ : InMux
    port map (
            O => \N__47871\,
            I => \N__47868\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__47868\,
            I => n1699
        );

    \I__10550\ : InMux
    port map (
            O => \N__47865\,
            I => n12564
        );

    \I__10549\ : CascadeMux
    port map (
            O => \N__47862\,
            I => \N__47858\
        );

    \I__10548\ : InMux
    port map (
            O => \N__47861\,
            I => \N__47854\
        );

    \I__10547\ : InMux
    port map (
            O => \N__47858\,
            I => \N__47851\
        );

    \I__10546\ : InMux
    port map (
            O => \N__47857\,
            I => \N__47848\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__47854\,
            I => n1631_adj_618
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__47851\,
            I => n1631_adj_618
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__47848\,
            I => n1631_adj_618
        );

    \I__10542\ : InMux
    port map (
            O => \N__47841\,
            I => \N__47838\
        );

    \I__10541\ : LocalMux
    port map (
            O => \N__47838\,
            I => n1698
        );

    \I__10540\ : InMux
    port map (
            O => \N__47835\,
            I => n12565
        );

    \I__10539\ : CascadeMux
    port map (
            O => \N__47832\,
            I => \N__47829\
        );

    \I__10538\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47825\
        );

    \I__10537\ : InMux
    port map (
            O => \N__47828\,
            I => \N__47822\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__47825\,
            I => n1630_adj_617
        );

    \I__10535\ : LocalMux
    port map (
            O => \N__47822\,
            I => n1630_adj_617
        );

    \I__10534\ : InMux
    port map (
            O => \N__47817\,
            I => \N__47814\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__47814\,
            I => n1697
        );

    \I__10532\ : InMux
    port map (
            O => \N__47811\,
            I => n12566
        );

    \I__10531\ : InMux
    port map (
            O => \N__47808\,
            I => n12567
        );

    \I__10530\ : InMux
    port map (
            O => \N__47805\,
            I => n12568
        );

    \I__10529\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47799\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__47799\,
            I => n1694
        );

    \I__10527\ : InMux
    port map (
            O => \N__47796\,
            I => n12569
        );

    \I__10526\ : InMux
    port map (
            O => \N__47793\,
            I => \bfn_15_18_0_\
        );

    \I__10525\ : InMux
    port map (
            O => \N__47790\,
            I => n12571
        );

    \I__10524\ : InMux
    port map (
            O => \N__47787\,
            I => \N__47780\
        );

    \I__10523\ : InMux
    port map (
            O => \N__47786\,
            I => \N__47780\
        );

    \I__10522\ : InMux
    port map (
            O => \N__47785\,
            I => \N__47777\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__47780\,
            I => \N__47774\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__47777\,
            I => n1624_adj_611
        );

    \I__10519\ : Odrv4
    port map (
            O => \N__47774\,
            I => n1624_adj_611
        );

    \I__10518\ : CascadeMux
    port map (
            O => \N__47769\,
            I => \N__47766\
        );

    \I__10517\ : InMux
    port map (
            O => \N__47766\,
            I => \N__47763\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__47763\,
            I => n1691
        );

    \I__10515\ : InMux
    port map (
            O => \N__47760\,
            I => n12572
        );

    \I__10514\ : InMux
    port map (
            O => \N__47757\,
            I => \N__47753\
        );

    \I__10513\ : InMux
    port map (
            O => \N__47756\,
            I => \N__47750\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__47753\,
            I => n43
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__47750\,
            I => n43
        );

    \I__10510\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47740\
        );

    \I__10509\ : InMux
    port map (
            O => \N__47744\,
            I => \N__47737\
        );

    \I__10508\ : InMux
    port map (
            O => \N__47743\,
            I => \N__47734\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__47740\,
            I => n23_adj_668
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__47737\,
            I => n23_adj_668
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__47734\,
            I => n23_adj_668
        );

    \I__10504\ : CascadeMux
    port map (
            O => \N__47727\,
            I => \n15132_cascade_\
        );

    \I__10503\ : InMux
    port map (
            O => \N__47724\,
            I => \N__47719\
        );

    \I__10502\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47716\
        );

    \I__10501\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47713\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__47719\,
            I => n25_adj_670
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__47716\,
            I => n25_adj_670
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__47713\,
            I => n25_adj_670
        );

    \I__10497\ : InMux
    port map (
            O => \N__47706\,
            I => \N__47703\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__47703\,
            I => \N__47700\
        );

    \I__10495\ : Odrv12
    port map (
            O => \N__47700\,
            I => n15110
        );

    \I__10494\ : SRMux
    port map (
            O => \N__47697\,
            I => \N__47694\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__47694\,
            I => \commutation_state_7__N_261\
        );

    \I__10492\ : InMux
    port map (
            O => \N__47691\,
            I => \N__47686\
        );

    \I__10491\ : InMux
    port map (
            O => \N__47690\,
            I => \N__47682\
        );

    \I__10490\ : InMux
    port map (
            O => \N__47689\,
            I => \N__47679\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__47686\,
            I => \N__47676\
        );

    \I__10488\ : InMux
    port map (
            O => \N__47685\,
            I => \N__47673\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__47682\,
            I => \N__47663\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__47679\,
            I => \N__47663\
        );

    \I__10485\ : Span4Mux_s1_v
    port map (
            O => \N__47676\,
            I => \N__47663\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__47673\,
            I => \N__47663\
        );

    \I__10483\ : InMux
    port map (
            O => \N__47672\,
            I => \N__47659\
        );

    \I__10482\ : Span4Mux_v
    port map (
            O => \N__47663\,
            I => \N__47656\
        );

    \I__10481\ : InMux
    port map (
            O => \N__47662\,
            I => \N__47653\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__47659\,
            I => \N__47650\
        );

    \I__10479\ : Span4Mux_v
    port map (
            O => \N__47656\,
            I => \N__47647\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__47653\,
            I => \N__47640\
        );

    \I__10477\ : Span12Mux_s9_v
    port map (
            O => \N__47650\,
            I => \N__47640\
        );

    \I__10476\ : Sp12to4
    port map (
            O => \N__47647\,
            I => \N__47640\
        );

    \I__10475\ : Odrv12
    port map (
            O => \N__47640\,
            I => h3
        );

    \I__10474\ : InMux
    port map (
            O => \N__47637\,
            I => \N__47630\
        );

    \I__10473\ : InMux
    port map (
            O => \N__47636\,
            I => \N__47627\
        );

    \I__10472\ : InMux
    port map (
            O => \N__47635\,
            I => \N__47622\
        );

    \I__10471\ : InMux
    port map (
            O => \N__47634\,
            I => \N__47622\
        );

    \I__10470\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47618\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__47630\,
            I => \N__47611\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__47627\,
            I => \N__47611\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__47622\,
            I => \N__47611\
        );

    \I__10466\ : InMux
    port map (
            O => \N__47621\,
            I => \N__47608\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__47618\,
            I => \N__47603\
        );

    \I__10464\ : Span4Mux_v
    port map (
            O => \N__47611\,
            I => \N__47603\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__47608\,
            I => h1
        );

    \I__10462\ : Odrv4
    port map (
            O => \N__47603\,
            I => h1
        );

    \I__10461\ : CascadeMux
    port map (
            O => \N__47598\,
            I => \N__47593\
        );

    \I__10460\ : InMux
    port map (
            O => \N__47597\,
            I => \N__47590\
        );

    \I__10459\ : InMux
    port map (
            O => \N__47596\,
            I => \N__47587\
        );

    \I__10458\ : InMux
    port map (
            O => \N__47593\,
            I => \N__47582\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__47590\,
            I => \N__47578\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__47587\,
            I => \N__47575\
        );

    \I__10455\ : InMux
    port map (
            O => \N__47586\,
            I => \N__47570\
        );

    \I__10454\ : InMux
    port map (
            O => \N__47585\,
            I => \N__47570\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__47582\,
            I => \N__47567\
        );

    \I__10452\ : InMux
    port map (
            O => \N__47581\,
            I => \N__47564\
        );

    \I__10451\ : Span4Mux_v
    port map (
            O => \N__47578\,
            I => \N__47559\
        );

    \I__10450\ : Span4Mux_s1_v
    port map (
            O => \N__47575\,
            I => \N__47559\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__47570\,
            I => \N__47556\
        );

    \I__10448\ : Span4Mux_s1_v
    port map (
            O => \N__47567\,
            I => \N__47553\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__47564\,
            I => h2
        );

    \I__10446\ : Odrv4
    port map (
            O => \N__47559\,
            I => h2
        );

    \I__10445\ : Odrv12
    port map (
            O => \N__47556\,
            I => h2
        );

    \I__10444\ : Odrv4
    port map (
            O => \N__47553\,
            I => h2
        );

    \I__10443\ : InMux
    port map (
            O => \N__47544\,
            I => \N__47539\
        );

    \I__10442\ : InMux
    port map (
            O => \N__47543\,
            I => \N__47536\
        );

    \I__10441\ : InMux
    port map (
            O => \N__47542\,
            I => \N__47533\
        );

    \I__10440\ : LocalMux
    port map (
            O => \N__47539\,
            I => \N__47530\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__47536\,
            I => \N__47527\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__47533\,
            I => \N__47524\
        );

    \I__10437\ : Span4Mux_h
    port map (
            O => \N__47530\,
            I => \N__47519\
        );

    \I__10436\ : Span4Mux_h
    port map (
            O => \N__47527\,
            I => \N__47519\
        );

    \I__10435\ : Span4Mux_h
    port map (
            O => \N__47524\,
            I => \N__47516\
        );

    \I__10434\ : Odrv4
    port map (
            O => \N__47519\,
            I => n302
        );

    \I__10433\ : Odrv4
    port map (
            O => \N__47516\,
            I => n302
        );

    \I__10432\ : InMux
    port map (
            O => \N__47511\,
            I => \N__47508\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__47508\,
            I => \N__47505\
        );

    \I__10430\ : Odrv4
    port map (
            O => \N__47505\,
            I => n1701
        );

    \I__10429\ : InMux
    port map (
            O => \N__47502\,
            I => \bfn_15_17_0_\
        );

    \I__10428\ : InMux
    port map (
            O => \N__47499\,
            I => \N__47496\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__47496\,
            I => n1700
        );

    \I__10426\ : InMux
    port map (
            O => \N__47493\,
            I => n12563
        );

    \I__10425\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47486\
        );

    \I__10424\ : InMux
    port map (
            O => \N__47489\,
            I => \N__47483\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__47486\,
            I => \N__47480\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__47483\,
            I => \N__47477\
        );

    \I__10421\ : Span4Mux_h
    port map (
            O => \N__47480\,
            I => \N__47474\
        );

    \I__10420\ : Odrv4
    port map (
            O => \N__47477\,
            I => pwm_setpoint_4
        );

    \I__10419\ : Odrv4
    port map (
            O => \N__47474\,
            I => pwm_setpoint_4
        );

    \I__10418\ : InMux
    port map (
            O => \N__47469\,
            I => \N__47465\
        );

    \I__10417\ : InMux
    port map (
            O => \N__47468\,
            I => \N__47462\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__47465\,
            I => \N__47459\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__47462\,
            I => pwm_counter_4
        );

    \I__10414\ : Odrv4
    port map (
            O => \N__47459\,
            I => pwm_counter_4
        );

    \I__10413\ : InMux
    port map (
            O => \N__47454\,
            I => \N__47451\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__47451\,
            I => \N__47448\
        );

    \I__10411\ : Odrv4
    port map (
            O => \N__47448\,
            I => n15150
        );

    \I__10410\ : InMux
    port map (
            O => \N__47445\,
            I => \N__47442\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__47442\,
            I => \N__47439\
        );

    \I__10408\ : Span4Mux_h
    port map (
            O => \N__47439\,
            I => \N__47436\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__47436\,
            I => \N__47432\
        );

    \I__10406\ : InMux
    port map (
            O => \N__47435\,
            I => \N__47429\
        );

    \I__10405\ : Odrv4
    port map (
            O => \N__47432\,
            I => n11_adj_660
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__47429\,
            I => n11_adj_660
        );

    \I__10403\ : CascadeMux
    port map (
            O => \N__47424\,
            I => \n9_adj_658_cascade_\
        );

    \I__10402\ : InMux
    port map (
            O => \N__47421\,
            I => \N__47418\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__47418\,
            I => \N__47414\
        );

    \I__10400\ : InMux
    port map (
            O => \N__47417\,
            I => \N__47411\
        );

    \I__10399\ : Span4Mux_h
    port map (
            O => \N__47414\,
            I => \N__47408\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__47411\,
            I => n13_adj_662
        );

    \I__10397\ : Odrv4
    port map (
            O => \N__47408\,
            I => n13_adj_662
        );

    \I__10396\ : CascadeMux
    port map (
            O => \N__47403\,
            I => \N__47400\
        );

    \I__10395\ : InMux
    port map (
            O => \N__47400\,
            I => \N__47397\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__47397\,
            I => \N__47394\
        );

    \I__10393\ : Span4Mux_h
    port map (
            O => \N__47394\,
            I => \N__47391\
        );

    \I__10392\ : Odrv4
    port map (
            O => \N__47391\,
            I => n15_adj_663
        );

    \I__10391\ : InMux
    port map (
            O => \N__47388\,
            I => \N__47385\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__47385\,
            I => n15205
        );

    \I__10389\ : CascadeMux
    port map (
            O => \N__47382\,
            I => \n15201_cascade_\
        );

    \I__10388\ : InMux
    port map (
            O => \N__47379\,
            I => \N__47376\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__47376\,
            I => \N__47373\
        );

    \I__10386\ : Span4Mux_v
    port map (
            O => \N__47373\,
            I => \N__47370\
        );

    \I__10385\ : Span4Mux_h
    port map (
            O => \N__47370\,
            I => \N__47367\
        );

    \I__10384\ : Odrv4
    port map (
            O => \N__47367\,
            I => n15261
        );

    \I__10383\ : InMux
    port map (
            O => \N__47364\,
            I => \N__47361\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__47361\,
            I => \N__47358\
        );

    \I__10381\ : Span4Mux_h
    port map (
            O => \N__47358\,
            I => \N__47354\
        );

    \I__10380\ : InMux
    port map (
            O => \N__47357\,
            I => \N__47351\
        );

    \I__10379\ : Odrv4
    port map (
            O => \N__47354\,
            I => pwm_setpoint_8
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__47351\,
            I => pwm_setpoint_8
        );

    \I__10377\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47342\
        );

    \I__10376\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47339\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__47342\,
            I => \N__47334\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__47339\,
            I => \N__47331\
        );

    \I__10373\ : InMux
    port map (
            O => \N__47338\,
            I => \N__47328\
        );

    \I__10372\ : InMux
    port map (
            O => \N__47337\,
            I => \N__47325\
        );

    \I__10371\ : Span4Mux_s3_v
    port map (
            O => \N__47334\,
            I => \N__47322\
        );

    \I__10370\ : Span4Mux_s3_v
    port map (
            O => \N__47331\,
            I => \N__47319\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__47328\,
            I => pwm_counter_8
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__47325\,
            I => pwm_counter_8
        );

    \I__10367\ : Odrv4
    port map (
            O => \N__47322\,
            I => pwm_counter_8
        );

    \I__10366\ : Odrv4
    port map (
            O => \N__47319\,
            I => pwm_counter_8
        );

    \I__10365\ : CascadeMux
    port map (
            O => \N__47310\,
            I => \N__47307\
        );

    \I__10364\ : InMux
    port map (
            O => \N__47307\,
            I => \N__47302\
        );

    \I__10363\ : InMux
    port map (
            O => \N__47306\,
            I => \N__47299\
        );

    \I__10362\ : InMux
    port map (
            O => \N__47305\,
            I => \N__47296\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__47302\,
            I => \N__47291\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__47299\,
            I => \N__47291\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__47296\,
            I => \N__47288\
        );

    \I__10358\ : Span4Mux_s1_v
    port map (
            O => \N__47291\,
            I => \N__47285\
        );

    \I__10357\ : Span4Mux_v
    port map (
            O => \N__47288\,
            I => \N__47282\
        );

    \I__10356\ : Odrv4
    port map (
            O => \N__47285\,
            I => pwm_setpoint_9
        );

    \I__10355\ : Odrv4
    port map (
            O => \N__47282\,
            I => pwm_setpoint_9
        );

    \I__10354\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47273\
        );

    \I__10353\ : InMux
    port map (
            O => \N__47276\,
            I => \N__47270\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__47273\,
            I => \N__47263\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__47270\,
            I => \N__47263\
        );

    \I__10350\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47260\
        );

    \I__10349\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47257\
        );

    \I__10348\ : Span4Mux_s3_v
    port map (
            O => \N__47263\,
            I => \N__47254\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__47260\,
            I => pwm_counter_9
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__47257\,
            I => pwm_counter_9
        );

    \I__10345\ : Odrv4
    port map (
            O => \N__47254\,
            I => pwm_counter_9
        );

    \I__10344\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47242\
        );

    \I__10343\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47239\
        );

    \I__10342\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47236\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__47242\,
            I => n21_adj_667
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__47239\,
            I => n21_adj_667
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__47236\,
            I => n21_adj_667
        );

    \I__10338\ : InMux
    port map (
            O => \N__47229\,
            I => \N__47225\
        );

    \I__10337\ : InMux
    port map (
            O => \N__47228\,
            I => \N__47222\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__47225\,
            I => n19_adj_666
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__47222\,
            I => n19_adj_666
        );

    \I__10334\ : CascadeMux
    port map (
            O => \N__47217\,
            I => \N__47214\
        );

    \I__10333\ : InMux
    port map (
            O => \N__47214\,
            I => \N__47211\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__47211\,
            I => \N__47207\
        );

    \I__10331\ : InMux
    port map (
            O => \N__47210\,
            I => \N__47204\
        );

    \I__10330\ : Odrv12
    port map (
            O => \N__47207\,
            I => n17_adj_665
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__47204\,
            I => n17_adj_665
        );

    \I__10328\ : InMux
    port map (
            O => \N__47199\,
            I => \N__47196\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__47196\,
            I => \N__47193\
        );

    \I__10326\ : Odrv4
    port map (
            O => \N__47193\,
            I => n9_adj_658
        );

    \I__10325\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47183\
        );

    \I__10324\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47183\
        );

    \I__10323\ : InMux
    port map (
            O => \N__47188\,
            I => \N__47180\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__47183\,
            I => \N__47173\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__47180\,
            I => \N__47173\
        );

    \I__10320\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47170\
        );

    \I__10319\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47167\
        );

    \I__10318\ : Span4Mux_s1_v
    port map (
            O => \N__47173\,
            I => \N__47164\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__47170\,
            I => pwm_counter_21
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__47167\,
            I => pwm_counter_21
        );

    \I__10315\ : Odrv4
    port map (
            O => \N__47164\,
            I => pwm_counter_21
        );

    \I__10314\ : InMux
    port map (
            O => \N__47157\,
            I => \N__47152\
        );

    \I__10313\ : InMux
    port map (
            O => \N__47156\,
            I => \N__47149\
        );

    \I__10312\ : InMux
    port map (
            O => \N__47155\,
            I => \N__47146\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__47152\,
            I => \N__47143\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__47149\,
            I => pwm_counter_12
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__47146\,
            I => pwm_counter_12
        );

    \I__10308\ : Odrv4
    port map (
            O => \N__47143\,
            I => pwm_counter_12
        );

    \I__10307\ : CascadeMux
    port map (
            O => \N__47136\,
            I => \PWM.n26_cascade_\
        );

    \I__10306\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47130\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__47130\,
            I => \PWM.n28\
        );

    \I__10304\ : CascadeMux
    port map (
            O => \N__47127\,
            I => \PWM.n29_cascade_\
        );

    \I__10303\ : InMux
    port map (
            O => \N__47124\,
            I => \N__47121\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__47121\,
            I => \PWM.n27\
        );

    \I__10301\ : SRMux
    port map (
            O => \N__47118\,
            I => \N__47115\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__47115\,
            I => \N__47112\
        );

    \I__10299\ : Span4Mux_v
    port map (
            O => \N__47112\,
            I => \N__47106\
        );

    \I__10298\ : SRMux
    port map (
            O => \N__47111\,
            I => \N__47103\
        );

    \I__10297\ : SRMux
    port map (
            O => \N__47110\,
            I => \N__47100\
        );

    \I__10296\ : SRMux
    port map (
            O => \N__47109\,
            I => \N__47097\
        );

    \I__10295\ : Odrv4
    port map (
            O => \N__47106\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__47103\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__47100\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__47097\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10291\ : InMux
    port map (
            O => \N__47088\,
            I => \N__47083\
        );

    \I__10290\ : InMux
    port map (
            O => \N__47087\,
            I => \N__47080\
        );

    \I__10289\ : InMux
    port map (
            O => \N__47086\,
            I => \N__47077\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__47083\,
            I => \N__47074\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__47080\,
            I => pwm_counter_19
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__47077\,
            I => pwm_counter_19
        );

    \I__10285\ : Odrv12
    port map (
            O => \N__47074\,
            I => pwm_counter_19
        );

    \I__10284\ : CascadeMux
    port map (
            O => \N__47067\,
            I => \N__47064\
        );

    \I__10283\ : InMux
    port map (
            O => \N__47064\,
            I => \N__47061\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__47061\,
            I => \PWM.n13995\
        );

    \I__10281\ : InMux
    port map (
            O => \N__47058\,
            I => \N__47055\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__47055\,
            I => \PWM.n17\
        );

    \I__10279\ : InMux
    port map (
            O => \N__47052\,
            I => \N__47048\
        );

    \I__10278\ : InMux
    port map (
            O => \N__47051\,
            I => \N__47045\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__47048\,
            I => pwm_counter_24
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__47045\,
            I => pwm_counter_24
        );

    \I__10275\ : InMux
    port map (
            O => \N__47040\,
            I => \N__47036\
        );

    \I__10274\ : InMux
    port map (
            O => \N__47039\,
            I => \N__47033\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__47036\,
            I => pwm_counter_29
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__47033\,
            I => pwm_counter_29
        );

    \I__10271\ : CascadeMux
    port map (
            O => \N__47028\,
            I => \N__47024\
        );

    \I__10270\ : InMux
    port map (
            O => \N__47027\,
            I => \N__47021\
        );

    \I__10269\ : InMux
    port map (
            O => \N__47024\,
            I => \N__47018\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__47021\,
            I => pwm_counter_27
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__47018\,
            I => pwm_counter_27
        );

    \I__10266\ : InMux
    port map (
            O => \N__47013\,
            I => \N__47009\
        );

    \I__10265\ : InMux
    port map (
            O => \N__47012\,
            I => \N__47006\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__47009\,
            I => pwm_counter_26
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__47006\,
            I => pwm_counter_26
        );

    \I__10262\ : InMux
    port map (
            O => \N__47001\,
            I => \N__46997\
        );

    \I__10261\ : InMux
    port map (
            O => \N__47000\,
            I => \N__46994\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__46997\,
            I => pwm_counter_30
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__46994\,
            I => pwm_counter_30
        );

    \I__10258\ : InMux
    port map (
            O => \N__46989\,
            I => \N__46985\
        );

    \I__10257\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46982\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__46985\,
            I => pwm_counter_25
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__46982\,
            I => pwm_counter_25
        );

    \I__10254\ : CascadeMux
    port map (
            O => \N__46977\,
            I => \n12_adj_566_cascade_\
        );

    \I__10253\ : InMux
    port map (
            O => \N__46974\,
            I => \N__46970\
        );

    \I__10252\ : InMux
    port map (
            O => \N__46973\,
            I => \N__46967\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__46970\,
            I => pwm_counter_28
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__46967\,
            I => pwm_counter_28
        );

    \I__10249\ : InMux
    port map (
            O => \N__46962\,
            I => \N__46959\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__46959\,
            I => n5162
        );

    \I__10247\ : CascadeMux
    port map (
            O => \N__46956\,
            I => \n5162_cascade_\
        );

    \I__10246\ : InMux
    port map (
            O => \N__46953\,
            I => \N__46948\
        );

    \I__10245\ : InMux
    port map (
            O => \N__46952\,
            I => \N__46945\
        );

    \I__10244\ : InMux
    port map (
            O => \N__46951\,
            I => \N__46942\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__46948\,
            I => pwm_counter_31
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__46945\,
            I => pwm_counter_31
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__46942\,
            I => pwm_counter_31
        );

    \I__10240\ : SRMux
    port map (
            O => \N__46935\,
            I => \N__46932\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__46932\,
            I => \N__46929\
        );

    \I__10238\ : Span4Mux_s3_v
    port map (
            O => \N__46929\,
            I => \N__46926\
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__46926\,
            I => n5164
        );

    \I__10236\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46920\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__46920\,
            I => \N__46917\
        );

    \I__10234\ : Span4Mux_h
    port map (
            O => \N__46917\,
            I => \N__46914\
        );

    \I__10233\ : Span4Mux_h
    port map (
            O => \N__46914\,
            I => \N__46911\
        );

    \I__10232\ : Odrv4
    port map (
            O => \N__46911\,
            I => \pwm_setpoint_23_N_171_8\
        );

    \I__10231\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46904\
        );

    \I__10230\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46901\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__46904\,
            I => \N__46898\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__46901\,
            I => \N__46895\
        );

    \I__10227\ : Span4Mux_v
    port map (
            O => \N__46898\,
            I => \N__46892\
        );

    \I__10226\ : Span4Mux_v
    port map (
            O => \N__46895\,
            I => \N__46889\
        );

    \I__10225\ : Span4Mux_h
    port map (
            O => \N__46892\,
            I => \N__46886\
        );

    \I__10224\ : Odrv4
    port map (
            O => \N__46889\,
            I => duty_8
        );

    \I__10223\ : Odrv4
    port map (
            O => \N__46886\,
            I => duty_8
        );

    \I__10222\ : CascadeMux
    port map (
            O => \N__46881\,
            I => \n14110_cascade_\
        );

    \I__10221\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46875\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__46875\,
            I => n10_adj_567
        );

    \I__10219\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46869\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__46869\,
            I => n15_adj_702
        );

    \I__10217\ : InMux
    port map (
            O => \N__46866\,
            I => \N__46863\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__46863\,
            I => \N__46860\
        );

    \I__10215\ : Odrv4
    port map (
            O => \N__46860\,
            I => n11853
        );

    \I__10214\ : InMux
    port map (
            O => \N__46857\,
            I => \N__46854\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__46854\,
            I => \N__46851\
        );

    \I__10212\ : Odrv4
    port map (
            O => \N__46851\,
            I => n23_adj_562
        );

    \I__10211\ : InMux
    port map (
            O => \N__46848\,
            I => \N__46845\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46842\
        );

    \I__10209\ : Span4Mux_h
    port map (
            O => \N__46842\,
            I => \N__46838\
        );

    \I__10208\ : InMux
    port map (
            O => \N__46841\,
            I => \N__46835\
        );

    \I__10207\ : Span4Mux_h
    port map (
            O => \N__46838\,
            I => \N__46832\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__46835\,
            I => pwm_setpoint_2
        );

    \I__10205\ : Odrv4
    port map (
            O => \N__46832\,
            I => pwm_setpoint_2
        );

    \I__10204\ : InMux
    port map (
            O => \N__46827\,
            I => \N__46823\
        );

    \I__10203\ : InMux
    port map (
            O => \N__46826\,
            I => \N__46820\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__46823\,
            I => \N__46817\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__46820\,
            I => pwm_setpoint_3
        );

    \I__10200\ : Odrv4
    port map (
            O => \N__46817\,
            I => pwm_setpoint_3
        );

    \I__10199\ : CascadeMux
    port map (
            O => \N__46812\,
            I => \N__46808\
        );

    \I__10198\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46805\
        );

    \I__10197\ : InMux
    port map (
            O => \N__46808\,
            I => \N__46802\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__46805\,
            I => pwm_counter_2
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__46802\,
            I => pwm_counter_2
        );

    \I__10194\ : InMux
    port map (
            O => \N__46797\,
            I => \N__46794\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__46794\,
            I => \N__46790\
        );

    \I__10192\ : InMux
    port map (
            O => \N__46793\,
            I => \N__46786\
        );

    \I__10191\ : Span4Mux_v
    port map (
            O => \N__46790\,
            I => \N__46783\
        );

    \I__10190\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46780\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__46786\,
            I => pwm_counter_3
        );

    \I__10188\ : Odrv4
    port map (
            O => \N__46783\,
            I => pwm_counter_3
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__46780\,
            I => pwm_counter_3
        );

    \I__10186\ : InMux
    port map (
            O => \N__46773\,
            I => \N__46768\
        );

    \I__10185\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46765\
        );

    \I__10184\ : InMux
    port map (
            O => \N__46771\,
            I => \N__46762\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__46768\,
            I => \N__46759\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__46765\,
            I => pwm_counter_5
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__46762\,
            I => pwm_counter_5
        );

    \I__10180\ : Odrv12
    port map (
            O => \N__46759\,
            I => pwm_counter_5
        );

    \I__10179\ : CascadeMux
    port map (
            O => \N__46752\,
            I => \N__46749\
        );

    \I__10178\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46745\
        );

    \I__10177\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46742\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__46745\,
            I => \N__46737\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46734\
        );

    \I__10174\ : InMux
    port map (
            O => \N__46741\,
            I => \N__46731\
        );

    \I__10173\ : InMux
    port map (
            O => \N__46740\,
            I => \N__46728\
        );

    \I__10172\ : Span4Mux_h
    port map (
            O => \N__46737\,
            I => \N__46725\
        );

    \I__10171\ : Span4Mux_h
    port map (
            O => \N__46734\,
            I => \N__46722\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__46731\,
            I => pwm_counter_7
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__46728\,
            I => pwm_counter_7
        );

    \I__10168\ : Odrv4
    port map (
            O => \N__46725\,
            I => pwm_counter_7
        );

    \I__10167\ : Odrv4
    port map (
            O => \N__46722\,
            I => pwm_counter_7
        );

    \I__10166\ : InMux
    port map (
            O => \N__46713\,
            I => \N__46710\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__46710\,
            I => \N__46704\
        );

    \I__10164\ : InMux
    port map (
            O => \N__46709\,
            I => \N__46701\
        );

    \I__10163\ : InMux
    port map (
            O => \N__46708\,
            I => \N__46698\
        );

    \I__10162\ : InMux
    port map (
            O => \N__46707\,
            I => \N__46695\
        );

    \I__10161\ : Span4Mux_h
    port map (
            O => \N__46704\,
            I => \N__46692\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__46701\,
            I => \N__46689\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__46698\,
            I => pwm_counter_6
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__46695\,
            I => pwm_counter_6
        );

    \I__10157\ : Odrv4
    port map (
            O => \N__46692\,
            I => pwm_counter_6
        );

    \I__10156\ : Odrv12
    port map (
            O => \N__46689\,
            I => pwm_counter_6
        );

    \I__10155\ : InMux
    port map (
            O => \N__46680\,
            I => \N__46675\
        );

    \I__10154\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46672\
        );

    \I__10153\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46669\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__46675\,
            I => \N__46666\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__46672\,
            I => pwm_counter_11
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__46669\,
            I => pwm_counter_11
        );

    \I__10149\ : Odrv4
    port map (
            O => \N__46666\,
            I => pwm_counter_11
        );

    \I__10148\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46654\
        );

    \I__10147\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46651\
        );

    \I__10146\ : InMux
    port map (
            O => \N__46657\,
            I => \N__46648\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__46654\,
            I => \N__46645\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__46651\,
            I => pwm_counter_10
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__46648\,
            I => pwm_counter_10
        );

    \I__10142\ : Odrv4
    port map (
            O => \N__46645\,
            I => pwm_counter_10
        );

    \I__10141\ : CascadeMux
    port map (
            O => \N__46638\,
            I => \N__46634\
        );

    \I__10140\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46630\
        );

    \I__10139\ : InMux
    port map (
            O => \N__46634\,
            I => \N__46627\
        );

    \I__10138\ : InMux
    port map (
            O => \N__46633\,
            I => \N__46624\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__46630\,
            I => \N__46621\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__46627\,
            I => pwm_counter_14
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__46624\,
            I => pwm_counter_14
        );

    \I__10134\ : Odrv4
    port map (
            O => \N__46621\,
            I => pwm_counter_14
        );

    \I__10133\ : InMux
    port map (
            O => \N__46614\,
            I => \N__46609\
        );

    \I__10132\ : InMux
    port map (
            O => \N__46613\,
            I => \N__46606\
        );

    \I__10131\ : InMux
    port map (
            O => \N__46612\,
            I => \N__46603\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__46609\,
            I => \N__46600\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__46606\,
            I => pwm_counter_20
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__46603\,
            I => pwm_counter_20
        );

    \I__10127\ : Odrv4
    port map (
            O => \N__46600\,
            I => pwm_counter_20
        );

    \I__10126\ : InMux
    port map (
            O => \N__46593\,
            I => \N__46586\
        );

    \I__10125\ : InMux
    port map (
            O => \N__46592\,
            I => \N__46581\
        );

    \I__10124\ : InMux
    port map (
            O => \N__46591\,
            I => \N__46581\
        );

    \I__10123\ : InMux
    port map (
            O => \N__46590\,
            I => \N__46578\
        );

    \I__10122\ : InMux
    port map (
            O => \N__46589\,
            I => \N__46575\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__46586\,
            I => \N__46572\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__46581\,
            I => \N__46569\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__46578\,
            I => pwm_counter_16
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__46575\,
            I => pwm_counter_16
        );

    \I__10117\ : Odrv12
    port map (
            O => \N__46572\,
            I => pwm_counter_16
        );

    \I__10116\ : Odrv4
    port map (
            O => \N__46569\,
            I => pwm_counter_16
        );

    \I__10115\ : InMux
    port map (
            O => \N__46560\,
            I => \N__46555\
        );

    \I__10114\ : InMux
    port map (
            O => \N__46559\,
            I => \N__46552\
        );

    \I__10113\ : InMux
    port map (
            O => \N__46558\,
            I => \N__46549\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__46555\,
            I => pwm_counter_17
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__46552\,
            I => pwm_counter_17
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__46549\,
            I => pwm_counter_17
        );

    \I__10109\ : CascadeMux
    port map (
            O => \N__46542\,
            I => \N__46538\
        );

    \I__10108\ : InMux
    port map (
            O => \N__46541\,
            I => \N__46534\
        );

    \I__10107\ : InMux
    port map (
            O => \N__46538\,
            I => \N__46531\
        );

    \I__10106\ : InMux
    port map (
            O => \N__46537\,
            I => \N__46528\
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__46534\,
            I => \N__46525\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__46531\,
            I => pwm_counter_13
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__46528\,
            I => pwm_counter_13
        );

    \I__10102\ : Odrv4
    port map (
            O => \N__46525\,
            I => pwm_counter_13
        );

    \I__10101\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46515\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__46515\,
            I => \N__46510\
        );

    \I__10099\ : InMux
    port map (
            O => \N__46514\,
            I => \N__46507\
        );

    \I__10098\ : InMux
    port map (
            O => \N__46513\,
            I => \N__46504\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__46510\,
            I => pwm_counter_23
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__46507\,
            I => pwm_counter_23
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__46504\,
            I => pwm_counter_23
        );

    \I__10094\ : InMux
    port map (
            O => \N__46497\,
            I => \N__46492\
        );

    \I__10093\ : InMux
    port map (
            O => \N__46496\,
            I => \N__46489\
        );

    \I__10092\ : InMux
    port map (
            O => \N__46495\,
            I => \N__46486\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__46492\,
            I => \N__46483\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__46489\,
            I => pwm_counter_22
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__46486\,
            I => pwm_counter_22
        );

    \I__10088\ : Odrv4
    port map (
            O => \N__46483\,
            I => pwm_counter_22
        );

    \I__10087\ : InMux
    port map (
            O => \N__46476\,
            I => \N__46471\
        );

    \I__10086\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46468\
        );

    \I__10085\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46465\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__46471\,
            I => \N__46462\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__46468\,
            I => pwm_counter_18
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__46465\,
            I => pwm_counter_18
        );

    \I__10081\ : Odrv4
    port map (
            O => \N__46462\,
            I => pwm_counter_18
        );

    \I__10080\ : CascadeMux
    port map (
            O => \N__46455\,
            I => \N__46451\
        );

    \I__10079\ : InMux
    port map (
            O => \N__46454\,
            I => \N__46448\
        );

    \I__10078\ : InMux
    port map (
            O => \N__46451\,
            I => \N__46445\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__46448\,
            I => \N__46441\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__46445\,
            I => \N__46438\
        );

    \I__10075\ : InMux
    port map (
            O => \N__46444\,
            I => \N__46435\
        );

    \I__10074\ : Span4Mux_v
    port map (
            O => \N__46441\,
            I => \N__46432\
        );

    \I__10073\ : Odrv4
    port map (
            O => \N__46438\,
            I => pwm_counter_15
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__46435\,
            I => pwm_counter_15
        );

    \I__10071\ : Odrv4
    port map (
            O => \N__46432\,
            I => pwm_counter_15
        );

    \I__10070\ : InMux
    port map (
            O => \N__46425\,
            I => \N__46421\
        );

    \I__10069\ : CascadeMux
    port map (
            O => \N__46424\,
            I => \N__46415\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__46421\,
            I => \N__46411\
        );

    \I__10067\ : CascadeMux
    port map (
            O => \N__46420\,
            I => \N__46405\
        );

    \I__10066\ : InMux
    port map (
            O => \N__46419\,
            I => \N__46399\
        );

    \I__10065\ : InMux
    port map (
            O => \N__46418\,
            I => \N__46399\
        );

    \I__10064\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46394\
        );

    \I__10063\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46394\
        );

    \I__10062\ : Span12Mux_h
    port map (
            O => \N__46411\,
            I => \N__46391\
        );

    \I__10061\ : InMux
    port map (
            O => \N__46410\,
            I => \N__46388\
        );

    \I__10060\ : InMux
    port map (
            O => \N__46409\,
            I => \N__46385\
        );

    \I__10059\ : InMux
    port map (
            O => \N__46408\,
            I => \N__46382\
        );

    \I__10058\ : InMux
    port map (
            O => \N__46405\,
            I => \N__46377\
        );

    \I__10057\ : InMux
    port map (
            O => \N__46404\,
            I => \N__46377\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__46399\,
            I => \N__46374\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__46394\,
            I => \N__46371\
        );

    \I__10054\ : Odrv12
    port map (
            O => \N__46391\,
            I => n1059
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__46388\,
            I => n1059
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__46385\,
            I => n1059
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__46382\,
            I => n1059
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__46377\,
            I => n1059
        );

    \I__10049\ : Odrv4
    port map (
            O => \N__46374\,
            I => n1059
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__46371\,
            I => n1059
        );

    \I__10047\ : InMux
    port map (
            O => \N__46356\,
            I => \N__46353\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__46353\,
            I => \N__46350\
        );

    \I__10045\ : Span4Mux_h
    port map (
            O => \N__46350\,
            I => \N__46347\
        );

    \I__10044\ : Span4Mux_h
    port map (
            O => \N__46347\,
            I => \N__46344\
        );

    \I__10043\ : Odrv4
    port map (
            O => \N__46344\,
            I => n15499
        );

    \I__10042\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46338\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__46338\,
            I => n14470
        );

    \I__10040\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46332\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__46332\,
            I => \N__46328\
        );

    \I__10038\ : CascadeMux
    port map (
            O => \N__46331\,
            I => \N__46324\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__46328\,
            I => \N__46321\
        );

    \I__10036\ : InMux
    port map (
            O => \N__46327\,
            I => \N__46318\
        );

    \I__10035\ : InMux
    port map (
            O => \N__46324\,
            I => \N__46315\
        );

    \I__10034\ : Sp12to4
    port map (
            O => \N__46321\,
            I => \N__46310\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__46318\,
            I => \N__46310\
        );

    \I__10032\ : LocalMux
    port map (
            O => \N__46315\,
            I => encoder0_position_21
        );

    \I__10031\ : Odrv12
    port map (
            O => \N__46310\,
            I => encoder0_position_21
        );

    \I__10030\ : CascadeMux
    port map (
            O => \N__46305\,
            I => \N__46302\
        );

    \I__10029\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46299\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__46299\,
            I => \N__46296\
        );

    \I__10027\ : Span4Mux_h
    port map (
            O => \N__46296\,
            I => \N__46293\
        );

    \I__10026\ : Odrv4
    port map (
            O => \N__46293\,
            I => n12_adj_633
        );

    \I__10025\ : CascadeMux
    port map (
            O => \N__46290\,
            I => \n16_adj_701_cascade_\
        );

    \I__10024\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46284\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__46284\,
            I => \N__46281\
        );

    \I__10022\ : Odrv12
    port map (
            O => \N__46281\,
            I => n24_adj_561
        );

    \I__10021\ : InMux
    port map (
            O => \N__46278\,
            I => \N__46275\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__46275\,
            I => \N__46272\
        );

    \I__10019\ : Odrv4
    port map (
            O => \N__46272\,
            I => n25
        );

    \I__10018\ : CascadeMux
    port map (
            O => \N__46269\,
            I => \n13932_cascade_\
        );

    \I__10017\ : InMux
    port map (
            O => \N__46266\,
            I => \N__46261\
        );

    \I__10016\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46258\
        );

    \I__10015\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46255\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__46261\,
            I => \N__46252\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__46258\,
            I => \N__46247\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__46255\,
            I => \N__46247\
        );

    \I__10011\ : Span4Mux_h
    port map (
            O => \N__46252\,
            I => \N__46244\
        );

    \I__10010\ : Odrv4
    port map (
            O => \N__46247\,
            I => n296
        );

    \I__10009\ : Odrv4
    port map (
            O => \N__46244\,
            I => n296
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__46239\,
            I => \N__46236\
        );

    \I__10007\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46233\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__46233\,
            I => \N__46230\
        );

    \I__10005\ : Odrv4
    port map (
            O => \N__46230\,
            I => n1101
        );

    \I__10004\ : CascadeMux
    port map (
            O => \N__46227\,
            I => \n1133_cascade_\
        );

    \I__10003\ : InMux
    port map (
            O => \N__46224\,
            I => \N__46221\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__46221\,
            I => n14428
        );

    \I__10001\ : CascadeMux
    port map (
            O => \N__46218\,
            I => \n12000_cascade_\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__46215\,
            I => \n1158_cascade_\
        );

    \I__9999\ : CascadeMux
    port map (
            O => \N__46212\,
            I => \n1232_cascade_\
        );

    \I__9998\ : InMux
    port map (
            O => \N__46209\,
            I => \N__46206\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__46206\,
            I => \N__46203\
        );

    \I__9996\ : Odrv12
    port map (
            O => \N__46203\,
            I => n12
        );

    \I__9995\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46177\
        );

    \I__9994\ : CascadeMux
    port map (
            O => \N__46199\,
            I => \N__46174\
        );

    \I__9993\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46166\
        );

    \I__9992\ : InMux
    port map (
            O => \N__46197\,
            I => \N__46166\
        );

    \I__9991\ : InMux
    port map (
            O => \N__46196\,
            I => \N__46166\
        );

    \I__9990\ : CascadeMux
    port map (
            O => \N__46195\,
            I => \N__46161\
        );

    \I__9989\ : InMux
    port map (
            O => \N__46194\,
            I => \N__46155\
        );

    \I__9988\ : InMux
    port map (
            O => \N__46193\,
            I => \N__46145\
        );

    \I__9987\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46145\
        );

    \I__9986\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46142\
        );

    \I__9985\ : InMux
    port map (
            O => \N__46190\,
            I => \N__46133\
        );

    \I__9984\ : InMux
    port map (
            O => \N__46189\,
            I => \N__46133\
        );

    \I__9983\ : InMux
    port map (
            O => \N__46188\,
            I => \N__46133\
        );

    \I__9982\ : InMux
    port map (
            O => \N__46187\,
            I => \N__46133\
        );

    \I__9981\ : InMux
    port map (
            O => \N__46186\,
            I => \N__46124\
        );

    \I__9980\ : InMux
    port map (
            O => \N__46185\,
            I => \N__46124\
        );

    \I__9979\ : InMux
    port map (
            O => \N__46184\,
            I => \N__46124\
        );

    \I__9978\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46124\
        );

    \I__9977\ : InMux
    port map (
            O => \N__46182\,
            I => \N__46121\
        );

    \I__9976\ : InMux
    port map (
            O => \N__46181\,
            I => \N__46118\
        );

    \I__9975\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46115\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__46177\,
            I => \N__46112\
        );

    \I__9973\ : InMux
    port map (
            O => \N__46174\,
            I => \N__46107\
        );

    \I__9972\ : InMux
    port map (
            O => \N__46173\,
            I => \N__46107\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__46166\,
            I => \N__46104\
        );

    \I__9970\ : CascadeMux
    port map (
            O => \N__46165\,
            I => \N__46099\
        );

    \I__9969\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46091\
        );

    \I__9968\ : InMux
    port map (
            O => \N__46161\,
            I => \N__46091\
        );

    \I__9967\ : InMux
    port map (
            O => \N__46160\,
            I => \N__46091\
        );

    \I__9966\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46086\
        );

    \I__9965\ : InMux
    port map (
            O => \N__46158\,
            I => \N__46086\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__46155\,
            I => \N__46083\
        );

    \I__9963\ : InMux
    port map (
            O => \N__46154\,
            I => \N__46076\
        );

    \I__9962\ : InMux
    port map (
            O => \N__46153\,
            I => \N__46076\
        );

    \I__9961\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46076\
        );

    \I__9960\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46071\
        );

    \I__9959\ : InMux
    port map (
            O => \N__46150\,
            I => \N__46071\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__46145\,
            I => \N__46062\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__46142\,
            I => \N__46062\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__46133\,
            I => \N__46062\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__46124\,
            I => \N__46062\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__46121\,
            I => \N__46057\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__46118\,
            I => \N__46054\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__46115\,
            I => \N__46050\
        );

    \I__9951\ : Span4Mux_v
    port map (
            O => \N__46112\,
            I => \N__46047\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__46107\,
            I => \N__46044\
        );

    \I__9949\ : Span4Mux_v
    port map (
            O => \N__46104\,
            I => \N__46041\
        );

    \I__9948\ : InMux
    port map (
            O => \N__46103\,
            I => \N__46032\
        );

    \I__9947\ : InMux
    port map (
            O => \N__46102\,
            I => \N__46032\
        );

    \I__9946\ : InMux
    port map (
            O => \N__46099\,
            I => \N__46032\
        );

    \I__9945\ : InMux
    port map (
            O => \N__46098\,
            I => \N__46032\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__46091\,
            I => \N__46024\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__46086\,
            I => \N__46024\
        );

    \I__9942\ : Span4Mux_v
    port map (
            O => \N__46083\,
            I => \N__46021\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__46076\,
            I => \N__46018\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__46071\,
            I => \N__46013\
        );

    \I__9939\ : Span4Mux_h
    port map (
            O => \N__46062\,
            I => \N__46013\
        );

    \I__9938\ : InMux
    port map (
            O => \N__46061\,
            I => \N__46010\
        );

    \I__9937\ : InMux
    port map (
            O => \N__46060\,
            I => \N__46007\
        );

    \I__9936\ : Span4Mux_h
    port map (
            O => \N__46057\,
            I => \N__46004\
        );

    \I__9935\ : Span12Mux_v
    port map (
            O => \N__46054\,
            I => \N__46001\
        );

    \I__9934\ : InMux
    port map (
            O => \N__46053\,
            I => \N__45998\
        );

    \I__9933\ : Span4Mux_v
    port map (
            O => \N__46050\,
            I => \N__45987\
        );

    \I__9932\ : Span4Mux_h
    port map (
            O => \N__46047\,
            I => \N__45987\
        );

    \I__9931\ : Span4Mux_v
    port map (
            O => \N__46044\,
            I => \N__45987\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__46041\,
            I => \N__45987\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__46032\,
            I => \N__45987\
        );

    \I__9928\ : InMux
    port map (
            O => \N__46031\,
            I => \N__45980\
        );

    \I__9927\ : InMux
    port map (
            O => \N__46030\,
            I => \N__45980\
        );

    \I__9926\ : InMux
    port map (
            O => \N__46029\,
            I => \N__45980\
        );

    \I__9925\ : Span4Mux_v
    port map (
            O => \N__46024\,
            I => \N__45971\
        );

    \I__9924\ : Span4Mux_h
    port map (
            O => \N__46021\,
            I => \N__45971\
        );

    \I__9923\ : Span4Mux_v
    port map (
            O => \N__46018\,
            I => \N__45971\
        );

    \I__9922\ : Span4Mux_v
    port map (
            O => \N__46013\,
            I => \N__45971\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__46010\,
            I => encoder0_position_31
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__46007\,
            I => encoder0_position_31
        );

    \I__9919\ : Odrv4
    port map (
            O => \N__46004\,
            I => encoder0_position_31
        );

    \I__9918\ : Odrv12
    port map (
            O => \N__46001\,
            I => encoder0_position_31
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__45998\,
            I => encoder0_position_31
        );

    \I__9916\ : Odrv4
    port map (
            O => \N__45987\,
            I => encoder0_position_31
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__45980\,
            I => encoder0_position_31
        );

    \I__9914\ : Odrv4
    port map (
            O => \N__45971\,
            I => encoder0_position_31
        );

    \I__9913\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45951\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__45951\,
            I => n1100
        );

    \I__9911\ : CascadeMux
    port map (
            O => \N__45948\,
            I => \N__45945\
        );

    \I__9910\ : InMux
    port map (
            O => \N__45945\,
            I => \N__45942\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__45942\,
            I => \N__45938\
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__45941\,
            I => \N__45935\
        );

    \I__9907\ : Span4Mux_h
    port map (
            O => \N__45938\,
            I => \N__45931\
        );

    \I__9906\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45928\
        );

    \I__9905\ : InMux
    port map (
            O => \N__45934\,
            I => \N__45925\
        );

    \I__9904\ : Odrv4
    port map (
            O => \N__45931\,
            I => n1033
        );

    \I__9903\ : LocalMux
    port map (
            O => \N__45928\,
            I => n1033
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__45925\,
            I => n1033
        );

    \I__9901\ : CascadeMux
    port map (
            O => \N__45918\,
            I => \n1132_cascade_\
        );

    \I__9900\ : CascadeMux
    port map (
            O => \N__45915\,
            I => \N__45911\
        );

    \I__9899\ : InMux
    port map (
            O => \N__45914\,
            I => \N__45908\
        );

    \I__9898\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45905\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__45908\,
            I => n1032
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__45905\,
            I => n1032
        );

    \I__9895\ : CascadeMux
    port map (
            O => \N__45900\,
            I => \N__45897\
        );

    \I__9894\ : InMux
    port map (
            O => \N__45897\,
            I => \N__45894\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__45894\,
            I => n1099
        );

    \I__9892\ : CascadeMux
    port map (
            O => \N__45891\,
            I => \n11908_cascade_\
        );

    \I__9891\ : CascadeMux
    port map (
            O => \N__45888\,
            I => \n13708_cascade_\
        );

    \I__9890\ : CascadeMux
    port map (
            O => \N__45885\,
            I => \n1356_cascade_\
        );

    \I__9889\ : CascadeMux
    port map (
            O => \N__45882\,
            I => \n1433_cascade_\
        );

    \I__9888\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45876\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__45876\,
            I => \N__45871\
        );

    \I__9886\ : CascadeMux
    port map (
            O => \N__45875\,
            I => \N__45868\
        );

    \I__9885\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45865\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__45871\,
            I => \N__45862\
        );

    \I__9883\ : InMux
    port map (
            O => \N__45868\,
            I => \N__45859\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__45865\,
            I => \N__45856\
        );

    \I__9881\ : Odrv4
    port map (
            O => \N__45862\,
            I => n1031
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__45859\,
            I => n1031
        );

    \I__9879\ : Odrv4
    port map (
            O => \N__45856\,
            I => n1031
        );

    \I__9878\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45846\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__45846\,
            I => n1098
        );

    \I__9876\ : CascadeMux
    port map (
            O => \N__45843\,
            I => \n1527_cascade_\
        );

    \I__9875\ : InMux
    port map (
            O => \N__45840\,
            I => \N__45837\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__45837\,
            I => n14288
        );

    \I__9873\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45831\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__45831\,
            I => \N__45828\
        );

    \I__9871\ : Span4Mux_v
    port map (
            O => \N__45828\,
            I => \N__45825\
        );

    \I__9870\ : Span4Mux_h
    port map (
            O => \N__45825\,
            I => \N__45822\
        );

    \I__9869\ : Odrv4
    port map (
            O => \N__45822\,
            I => n14
        );

    \I__9868\ : CascadeMux
    port map (
            O => \N__45819\,
            I => \n1324_cascade_\
        );

    \I__9867\ : InMux
    port map (
            O => \N__45816\,
            I => \N__45810\
        );

    \I__9866\ : InMux
    port map (
            O => \N__45815\,
            I => \N__45810\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__45810\,
            I => \N__45806\
        );

    \I__9864\ : CascadeMux
    port map (
            O => \N__45809\,
            I => \N__45803\
        );

    \I__9863\ : Span4Mux_h
    port map (
            O => \N__45806\,
            I => \N__45800\
        );

    \I__9862\ : InMux
    port map (
            O => \N__45803\,
            I => \N__45797\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__45800\,
            I => \N__45794\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__45797\,
            I => encoder0_position_19
        );

    \I__9859\ : Odrv4
    port map (
            O => \N__45794\,
            I => encoder0_position_19
        );

    \I__9858\ : CascadeMux
    port map (
            O => \N__45789\,
            I => \N__45786\
        );

    \I__9857\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45783\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__45783\,
            I => \N__45780\
        );

    \I__9855\ : Span4Mux_h
    port map (
            O => \N__45780\,
            I => \N__45777\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__45777\,
            I => n14_adj_635
        );

    \I__9853\ : CascadeMux
    port map (
            O => \N__45774\,
            I => \n1531_cascade_\
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__45771\,
            I => \N__45768\
        );

    \I__9851\ : InMux
    port map (
            O => \N__45768\,
            I => \N__45765\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__45765\,
            I => n1592
        );

    \I__9849\ : CascadeMux
    port map (
            O => \N__45762\,
            I => \N__45758\
        );

    \I__9848\ : InMux
    port map (
            O => \N__45761\,
            I => \N__45755\
        );

    \I__9847\ : InMux
    port map (
            O => \N__45758\,
            I => \N__45752\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__45755\,
            I => n1533
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__45752\,
            I => n1533
        );

    \I__9844\ : InMux
    port map (
            O => \N__45747\,
            I => \N__45744\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__45744\,
            I => n1600
        );

    \I__9842\ : CascadeMux
    port map (
            O => \N__45741\,
            I => \n1533_cascade_\
        );

    \I__9841\ : InMux
    port map (
            O => \N__45738\,
            I => \N__45735\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__45735\,
            I => \N__45732\
        );

    \I__9839\ : Span4Mux_h
    port map (
            O => \N__45732\,
            I => \N__45729\
        );

    \I__9838\ : Span4Mux_h
    port map (
            O => \N__45729\,
            I => \N__45726\
        );

    \I__9837\ : Span4Mux_v
    port map (
            O => \N__45726\,
            I => \N__45722\
        );

    \I__9836\ : InMux
    port map (
            O => \N__45725\,
            I => \N__45719\
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__45722\,
            I => n15582
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__45719\,
            I => n15582
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__45714\,
            I => \n14294_cascade_\
        );

    \I__9832\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45708\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__45708\,
            I => n11974
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__45705\,
            I => \n11902_cascade_\
        );

    \I__9829\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45699\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__45699\,
            I => n13736
        );

    \I__9827\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__45693\,
            I => n1599
        );

    \I__9825\ : InMux
    port map (
            O => \N__45690\,
            I => \N__45687\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__45687\,
            I => \N__45683\
        );

    \I__9823\ : CascadeMux
    port map (
            O => \N__45686\,
            I => \N__45680\
        );

    \I__9822\ : Span4Mux_v
    port map (
            O => \N__45683\,
            I => \N__45677\
        );

    \I__9821\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45674\
        );

    \I__9820\ : Odrv4
    port map (
            O => \N__45677\,
            I => n1731
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__45674\,
            I => n1731
        );

    \I__9818\ : InMux
    port map (
            O => \N__45669\,
            I => \N__45666\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__45666\,
            I => \N__45662\
        );

    \I__9816\ : CascadeMux
    port map (
            O => \N__45665\,
            I => \N__45659\
        );

    \I__9815\ : Span4Mux_h
    port map (
            O => \N__45662\,
            I => \N__45655\
        );

    \I__9814\ : InMux
    port map (
            O => \N__45659\,
            I => \N__45652\
        );

    \I__9813\ : InMux
    port map (
            O => \N__45658\,
            I => \N__45649\
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__45655\,
            I => n1733
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__45652\,
            I => n1733
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__45649\,
            I => n1733
        );

    \I__9809\ : InMux
    port map (
            O => \N__45642\,
            I => \N__45638\
        );

    \I__9808\ : InMux
    port map (
            O => \N__45641\,
            I => \N__45635\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__45638\,
            I => \N__45631\
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__45635\,
            I => \N__45628\
        );

    \I__9805\ : InMux
    port map (
            O => \N__45634\,
            I => \N__45625\
        );

    \I__9804\ : Span4Mux_h
    port map (
            O => \N__45631\,
            I => \N__45622\
        );

    \I__9803\ : Span4Mux_v
    port map (
            O => \N__45628\,
            I => \N__45619\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__45625\,
            I => n303
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__45622\,
            I => n303
        );

    \I__9800\ : Odrv4
    port map (
            O => \N__45619\,
            I => n303
        );

    \I__9799\ : CascadeMux
    port map (
            O => \N__45612\,
            I => \n1731_cascade_\
        );

    \I__9798\ : InMux
    port map (
            O => \N__45609\,
            I => \N__45606\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__45606\,
            I => \N__45603\
        );

    \I__9796\ : Span4Mux_h
    port map (
            O => \N__45603\,
            I => \N__45600\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__45600\,
            I => n11970
        );

    \I__9794\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45594\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__45594\,
            I => \N__45590\
        );

    \I__9792\ : CascadeMux
    port map (
            O => \N__45593\,
            I => \N__45587\
        );

    \I__9791\ : Span4Mux_h
    port map (
            O => \N__45590\,
            I => \N__45583\
        );

    \I__9790\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45580\
        );

    \I__9789\ : InMux
    port map (
            O => \N__45586\,
            I => \N__45577\
        );

    \I__9788\ : Odrv4
    port map (
            O => \N__45583\,
            I => n1732
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__45580\,
            I => n1732
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__45577\,
            I => n1732
        );

    \I__9785\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45567\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__45567\,
            I => n1590
        );

    \I__9783\ : InMux
    port map (
            O => \N__45564\,
            I => \N__45561\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__45561\,
            I => n1589
        );

    \I__9781\ : CascadeMux
    port map (
            O => \N__45558\,
            I => \N__45554\
        );

    \I__9780\ : CascadeMux
    port map (
            O => \N__45557\,
            I => \N__45551\
        );

    \I__9779\ : InMux
    port map (
            O => \N__45554\,
            I => \N__45548\
        );

    \I__9778\ : InMux
    port map (
            O => \N__45551\,
            I => \N__45545\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__45548\,
            I => n1531
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__45545\,
            I => n1531
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__45540\,
            I => \n14910_cascade_\
        );

    \I__9774\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45532\
        );

    \I__9773\ : CascadeMux
    port map (
            O => \N__45536\,
            I => \N__45529\
        );

    \I__9772\ : InMux
    port map (
            O => \N__45535\,
            I => \N__45526\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__45532\,
            I => \N__45523\
        );

    \I__9770\ : InMux
    port map (
            O => \N__45529\,
            I => \N__45520\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__45526\,
            I => \N__45515\
        );

    \I__9768\ : Span4Mux_v
    port map (
            O => \N__45523\,
            I => \N__45515\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__45520\,
            I => n1730
        );

    \I__9766\ : Odrv4
    port map (
            O => \N__45515\,
            I => n1730
        );

    \I__9765\ : CascadeMux
    port map (
            O => \N__45510\,
            I => \n14514_cascade_\
        );

    \I__9764\ : CascadeMux
    port map (
            O => \N__45507\,
            I => \n1653_cascade_\
        );

    \I__9763\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45501\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__45501\,
            I => n1598
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__45498\,
            I => \n1630_adj_617_cascade_\
        );

    \I__9760\ : CascadeMux
    port map (
            O => \N__45495\,
            I => \N__45490\
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__45494\,
            I => \N__45487\
        );

    \I__9758\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45482\
        );

    \I__9757\ : InMux
    port map (
            O => \N__45490\,
            I => \N__45482\
        );

    \I__9756\ : InMux
    port map (
            O => \N__45487\,
            I => \N__45479\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__45482\,
            I => \N__45476\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__45479\,
            I => n1729
        );

    \I__9753\ : Odrv12
    port map (
            O => \N__45476\,
            I => n1729
        );

    \I__9752\ : InMux
    port map (
            O => \N__45471\,
            I => \N__45467\
        );

    \I__9751\ : InMux
    port map (
            O => \N__45470\,
            I => \N__45464\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__45467\,
            I => pwm_setpoint_11
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__45464\,
            I => pwm_setpoint_11
        );

    \I__9748\ : InMux
    port map (
            O => \N__45459\,
            I => \N__45455\
        );

    \I__9747\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45452\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__45455\,
            I => \N__45449\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__45452\,
            I => pwm_setpoint_12
        );

    \I__9744\ : Odrv4
    port map (
            O => \N__45449\,
            I => pwm_setpoint_12
        );

    \I__9743\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45440\
        );

    \I__9742\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45437\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__45440\,
            I => pwm_setpoint_20
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__45437\,
            I => pwm_setpoint_20
        );

    \I__9739\ : InMux
    port map (
            O => \N__45432\,
            I => \N__45429\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__45429\,
            I => n41
        );

    \I__9737\ : CascadeMux
    port map (
            O => \N__45426\,
            I => \n41_cascade_\
        );

    \I__9736\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45420\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__45420\,
            I => \N__45417\
        );

    \I__9734\ : Odrv4
    port map (
            O => \N__45417\,
            I => n15265
        );

    \I__9733\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45411\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__45411\,
            I => n15112
        );

    \I__9731\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45405\
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__45405\,
            I => \N__45402\
        );

    \I__9729\ : Span4Mux_h
    port map (
            O => \N__45402\,
            I => \N__45399\
        );

    \I__9728\ : Odrv4
    port map (
            O => \N__45399\,
            I => pwm_setpoint_23
        );

    \I__9727\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45393\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__45393\,
            I => n15257
        );

    \I__9725\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45387\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__45387\,
            I => \N__45384\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__45384\,
            I => n15108
        );

    \I__9722\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45374\
        );

    \I__9721\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45374\
        );

    \I__9720\ : InMux
    port map (
            O => \N__45379\,
            I => \N__45371\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__45374\,
            I => pwm_setpoint_21
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__45371\,
            I => pwm_setpoint_21
        );

    \I__9717\ : InMux
    port map (
            O => \N__45366\,
            I => \N__45362\
        );

    \I__9716\ : InMux
    port map (
            O => \N__45365\,
            I => \N__45359\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__45362\,
            I => \N__45356\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__45359\,
            I => \N__45353\
        );

    \I__9713\ : Odrv4
    port map (
            O => \N__45356\,
            I => pwm_setpoint_19
        );

    \I__9712\ : Odrv4
    port map (
            O => \N__45353\,
            I => pwm_setpoint_19
        );

    \I__9711\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45344\
        );

    \I__9710\ : InMux
    port map (
            O => \N__45347\,
            I => \N__45341\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__45344\,
            I => \N__45338\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__45341\,
            I => n39
        );

    \I__9707\ : Odrv4
    port map (
            O => \N__45338\,
            I => n39
        );

    \I__9706\ : InMux
    port map (
            O => \N__45333\,
            I => \PWM.n13082\
        );

    \I__9705\ : InMux
    port map (
            O => \N__45330\,
            I => \PWM.n13083\
        );

    \I__9704\ : InMux
    port map (
            O => \N__45327\,
            I => \PWM.n13084\
        );

    \I__9703\ : InMux
    port map (
            O => \N__45324\,
            I => \PWM.n13085\
        );

    \I__9702\ : InMux
    port map (
            O => \N__45321\,
            I => \PWM.n13086\
        );

    \I__9701\ : CEMux
    port map (
            O => \N__45318\,
            I => \N__45315\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__45315\,
            I => \N__45312\
        );

    \I__9699\ : Span4Mux_h
    port map (
            O => \N__45312\,
            I => \N__45309\
        );

    \I__9698\ : Odrv4
    port map (
            O => \N__45309\,
            I => n6_adj_717
        );

    \I__9697\ : InMux
    port map (
            O => \N__45306\,
            I => \N__45303\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__45303\,
            I => \N__45299\
        );

    \I__9695\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45296\
        );

    \I__9694\ : Span4Mux_h
    port map (
            O => \N__45299\,
            I => \N__45293\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__45296\,
            I => \N__45290\
        );

    \I__9692\ : Odrv4
    port map (
            O => \N__45293\,
            I => pwm_setpoint_5
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__45290\,
            I => pwm_setpoint_5
        );

    \I__9690\ : InMux
    port map (
            O => \N__45285\,
            I => \N__45281\
        );

    \I__9689\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45278\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__45281\,
            I => \N__45275\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__45278\,
            I => pwm_setpoint_6
        );

    \I__9686\ : Odrv12
    port map (
            O => \N__45275\,
            I => pwm_setpoint_6
        );

    \I__9685\ : InMux
    port map (
            O => \N__45270\,
            I => \N__45266\
        );

    \I__9684\ : InMux
    port map (
            O => \N__45269\,
            I => \N__45263\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__45266\,
            I => \N__45258\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__45263\,
            I => \N__45258\
        );

    \I__9681\ : Odrv12
    port map (
            O => \N__45258\,
            I => pwm_setpoint_10
        );

    \I__9680\ : InMux
    port map (
            O => \N__45255\,
            I => \PWM.n13073\
        );

    \I__9679\ : InMux
    port map (
            O => \N__45252\,
            I => \PWM.n13074\
        );

    \I__9678\ : InMux
    port map (
            O => \N__45249\,
            I => \PWM.n13075\
        );

    \I__9677\ : InMux
    port map (
            O => \N__45246\,
            I => \PWM.n13076\
        );

    \I__9676\ : InMux
    port map (
            O => \N__45243\,
            I => \PWM.n13077\
        );

    \I__9675\ : InMux
    port map (
            O => \N__45240\,
            I => \PWM.n13078\
        );

    \I__9674\ : InMux
    port map (
            O => \N__45237\,
            I => \bfn_13_29_0_\
        );

    \I__9673\ : InMux
    port map (
            O => \N__45234\,
            I => \PWM.n13080\
        );

    \I__9672\ : InMux
    port map (
            O => \N__45231\,
            I => \PWM.n13081\
        );

    \I__9671\ : InMux
    port map (
            O => \N__45228\,
            I => \PWM.n13064\
        );

    \I__9670\ : InMux
    port map (
            O => \N__45225\,
            I => \PWM.n13065\
        );

    \I__9669\ : InMux
    port map (
            O => \N__45222\,
            I => \PWM.n13066\
        );

    \I__9668\ : InMux
    port map (
            O => \N__45219\,
            I => \PWM.n13067\
        );

    \I__9667\ : InMux
    port map (
            O => \N__45216\,
            I => \PWM.n13068\
        );

    \I__9666\ : InMux
    port map (
            O => \N__45213\,
            I => \PWM.n13069\
        );

    \I__9665\ : InMux
    port map (
            O => \N__45210\,
            I => \PWM.n13070\
        );

    \I__9664\ : InMux
    port map (
            O => \N__45207\,
            I => \bfn_13_28_0_\
        );

    \I__9663\ : InMux
    port map (
            O => \N__45204\,
            I => \PWM.n13072\
        );

    \I__9662\ : CascadeMux
    port map (
            O => \N__45201\,
            I => \N__45198\
        );

    \I__9661\ : InMux
    port map (
            O => \N__45198\,
            I => \N__45194\
        );

    \I__9660\ : InMux
    port map (
            O => \N__45197\,
            I => \N__45191\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__45194\,
            I => \N__45188\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__45191\,
            I => pwm_counter_0
        );

    \I__9657\ : Odrv12
    port map (
            O => \N__45188\,
            I => pwm_counter_0
        );

    \I__9656\ : InMux
    port map (
            O => \N__45183\,
            I => \bfn_13_26_0_\
        );

    \I__9655\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45176\
        );

    \I__9654\ : InMux
    port map (
            O => \N__45179\,
            I => \N__45173\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__45176\,
            I => \N__45170\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__45173\,
            I => pwm_counter_1
        );

    \I__9651\ : Odrv12
    port map (
            O => \N__45170\,
            I => pwm_counter_1
        );

    \I__9650\ : InMux
    port map (
            O => \N__45165\,
            I => \PWM.n13056\
        );

    \I__9649\ : InMux
    port map (
            O => \N__45162\,
            I => \PWM.n13057\
        );

    \I__9648\ : InMux
    port map (
            O => \N__45159\,
            I => \PWM.n13058\
        );

    \I__9647\ : InMux
    port map (
            O => \N__45156\,
            I => \PWM.n13059\
        );

    \I__9646\ : InMux
    port map (
            O => \N__45153\,
            I => \PWM.n13060\
        );

    \I__9645\ : InMux
    port map (
            O => \N__45150\,
            I => \PWM.n13061\
        );

    \I__9644\ : InMux
    port map (
            O => \N__45147\,
            I => \PWM.n13062\
        );

    \I__9643\ : InMux
    port map (
            O => \N__45144\,
            I => \bfn_13_27_0_\
        );

    \I__9642\ : CascadeMux
    port map (
            O => \N__45141\,
            I => \N__45137\
        );

    \I__9641\ : CascadeMux
    port map (
            O => \N__45140\,
            I => \N__45134\
        );

    \I__9640\ : InMux
    port map (
            O => \N__45137\,
            I => \N__45130\
        );

    \I__9639\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45125\
        );

    \I__9638\ : InMux
    port map (
            O => \N__45133\,
            I => \N__45125\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__45130\,
            I => n1029
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__45125\,
            I => n1029
        );

    \I__9635\ : InMux
    port map (
            O => \N__45120\,
            I => \N__45117\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__45117\,
            I => n1096
        );

    \I__9633\ : InMux
    port map (
            O => \N__45114\,
            I => n12504
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__45111\,
            I => \N__45108\
        );

    \I__9631\ : InMux
    port map (
            O => \N__45108\,
            I => \N__45104\
        );

    \I__9630\ : InMux
    port map (
            O => \N__45107\,
            I => \N__45101\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__45104\,
            I => n1028
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__45101\,
            I => n1028
        );

    \I__9627\ : InMux
    port map (
            O => \N__45096\,
            I => \N__45093\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__45093\,
            I => n1095
        );

    \I__9625\ : InMux
    port map (
            O => \N__45090\,
            I => n12505
        );

    \I__9624\ : CascadeMux
    port map (
            O => \N__45087\,
            I => \N__45084\
        );

    \I__9623\ : InMux
    port map (
            O => \N__45084\,
            I => \N__45079\
        );

    \I__9622\ : InMux
    port map (
            O => \N__45083\,
            I => \N__45074\
        );

    \I__9621\ : InMux
    port map (
            O => \N__45082\,
            I => \N__45074\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__45079\,
            I => n1027
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__45074\,
            I => n1027
        );

    \I__9618\ : InMux
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__45066\,
            I => n1094
        );

    \I__9616\ : InMux
    port map (
            O => \N__45063\,
            I => n12506
        );

    \I__9615\ : InMux
    port map (
            O => \N__45060\,
            I => \bfn_13_24_0_\
        );

    \I__9614\ : CascadeMux
    port map (
            O => \N__45057\,
            I => \N__45053\
        );

    \I__9613\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45048\
        );

    \I__9612\ : InMux
    port map (
            O => \N__45053\,
            I => \N__45048\
        );

    \I__9611\ : LocalMux
    port map (
            O => \N__45048\,
            I => \N__45044\
        );

    \I__9610\ : InMux
    port map (
            O => \N__45047\,
            I => \N__45041\
        );

    \I__9609\ : Odrv4
    port map (
            O => \N__45044\,
            I => n1026
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__45041\,
            I => n1026
        );

    \I__9607\ : InMux
    port map (
            O => \N__45036\,
            I => \N__45033\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__45033\,
            I => n1093
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__45030\,
            I => \N__45026\
        );

    \I__9604\ : InMux
    port map (
            O => \N__45029\,
            I => \N__45022\
        );

    \I__9603\ : InMux
    port map (
            O => \N__45026\,
            I => \N__45019\
        );

    \I__9602\ : InMux
    port map (
            O => \N__45025\,
            I => \N__45016\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__45022\,
            I => n1030
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__45019\,
            I => n1030
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__45016\,
            I => n1030
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__45009\,
            I => \N__45006\
        );

    \I__9597\ : InMux
    port map (
            O => \N__45006\,
            I => \N__45003\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__45003\,
            I => n1097
        );

    \I__9595\ : CascadeMux
    port map (
            O => \N__45000\,
            I => \n13716_cascade_\
        );

    \I__9594\ : CascadeMux
    port map (
            O => \N__44997\,
            I => \n1059_cascade_\
        );

    \I__9593\ : CascadeMux
    port map (
            O => \N__44994\,
            I => \n1126_cascade_\
        );

    \I__9592\ : InMux
    port map (
            O => \N__44991\,
            I => \N__44988\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__44988\,
            I => \N__44984\
        );

    \I__9590\ : CascadeMux
    port map (
            O => \N__44987\,
            I => \N__44981\
        );

    \I__9589\ : Span4Mux_v
    port map (
            O => \N__44984\,
            I => \N__44977\
        );

    \I__9588\ : InMux
    port map (
            O => \N__44981\,
            I => \N__44974\
        );

    \I__9587\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44971\
        );

    \I__9586\ : Odrv4
    port map (
            O => \N__44977\,
            I => n928
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__44974\,
            I => n928
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__44971\,
            I => n928
        );

    \I__9583\ : CascadeMux
    port map (
            O => \N__44964\,
            I => \N__44960\
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__44963\,
            I => \N__44957\
        );

    \I__9581\ : InMux
    port map (
            O => \N__44960\,
            I => \N__44949\
        );

    \I__9580\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44944\
        );

    \I__9579\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44944\
        );

    \I__9578\ : InMux
    port map (
            O => \N__44955\,
            I => \N__44941\
        );

    \I__9577\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44934\
        );

    \I__9576\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44934\
        );

    \I__9575\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44934\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__44949\,
            I => n960
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__44944\,
            I => n960
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__44941\,
            I => n960
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__44934\,
            I => n960
        );

    \I__9570\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44922\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__44922\,
            I => n995
        );

    \I__9568\ : InMux
    port map (
            O => \N__44919\,
            I => \bfn_13_23_0_\
        );

    \I__9567\ : InMux
    port map (
            O => \N__44916\,
            I => n12500
        );

    \I__9566\ : InMux
    port map (
            O => \N__44913\,
            I => n12501
        );

    \I__9565\ : InMux
    port map (
            O => \N__44910\,
            I => n12502
        );

    \I__9564\ : InMux
    port map (
            O => \N__44907\,
            I => n12503
        );

    \I__9563\ : InMux
    port map (
            O => \N__44904\,
            I => \N__44901\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__44901\,
            I => \N__44898\
        );

    \I__9561\ : Odrv12
    port map (
            O => \N__44898\,
            I => n27
        );

    \I__9560\ : InMux
    port map (
            O => \N__44895\,
            I => \N__44892\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__44892\,
            I => \N__44888\
        );

    \I__9558\ : InMux
    port map (
            O => \N__44891\,
            I => \N__44884\
        );

    \I__9557\ : Span4Mux_h
    port map (
            O => \N__44888\,
            I => \N__44881\
        );

    \I__9556\ : InMux
    port map (
            O => \N__44887\,
            I => \N__44878\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__44884\,
            I => encoder0_position_6
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__44881\,
            I => encoder0_position_6
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__44878\,
            I => encoder0_position_6
        );

    \I__9552\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44867\
        );

    \I__9551\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44863\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__44867\,
            I => \N__44860\
        );

    \I__9549\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44857\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__44863\,
            I => \N__44854\
        );

    \I__9547\ : Span4Mux_v
    port map (
            O => \N__44860\,
            I => \N__44851\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__44857\,
            I => \N__44848\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__44854\,
            I => \N__44845\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__44851\,
            I => \N__44842\
        );

    \I__9543\ : Span12Mux_s8_v
    port map (
            O => \N__44848\,
            I => \N__44839\
        );

    \I__9542\ : Span4Mux_h
    port map (
            O => \N__44845\,
            I => \N__44836\
        );

    \I__9541\ : Span4Mux_h
    port map (
            O => \N__44842\,
            I => \N__44833\
        );

    \I__9540\ : Span12Mux_h
    port map (
            O => \N__44839\,
            I => \N__44830\
        );

    \I__9539\ : Span4Mux_h
    port map (
            O => \N__44836\,
            I => \N__44827\
        );

    \I__9538\ : Span4Mux_h
    port map (
            O => \N__44833\,
            I => \N__44824\
        );

    \I__9537\ : Odrv12
    port map (
            O => \N__44830\,
            I => n313
        );

    \I__9536\ : Odrv4
    port map (
            O => \N__44827\,
            I => n313
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__44824\,
            I => n313
        );

    \I__9534\ : InMux
    port map (
            O => \N__44817\,
            I => \N__44814\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__44814\,
            I => \N__44811\
        );

    \I__9532\ : Span4Mux_h
    port map (
            O => \N__44811\,
            I => \N__44808\
        );

    \I__9531\ : Odrv4
    port map (
            O => \N__44808\,
            I => n11
        );

    \I__9530\ : InMux
    port map (
            O => \N__44805\,
            I => \N__44799\
        );

    \I__9529\ : InMux
    port map (
            O => \N__44804\,
            I => \N__44799\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__44799\,
            I => \N__44795\
        );

    \I__9527\ : InMux
    port map (
            O => \N__44798\,
            I => \N__44792\
        );

    \I__9526\ : Span4Mux_h
    port map (
            O => \N__44795\,
            I => \N__44789\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__44792\,
            I => encoder0_position_22
        );

    \I__9524\ : Odrv4
    port map (
            O => \N__44789\,
            I => encoder0_position_22
        );

    \I__9523\ : CascadeMux
    port map (
            O => \N__44784\,
            I => \N__44781\
        );

    \I__9522\ : InMux
    port map (
            O => \N__44781\,
            I => \N__44778\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__44778\,
            I => \N__44775\
        );

    \I__9520\ : Span4Mux_h
    port map (
            O => \N__44775\,
            I => \N__44772\
        );

    \I__9519\ : Odrv4
    port map (
            O => \N__44772\,
            I => n11_adj_632
        );

    \I__9518\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44766\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__44766\,
            I => \N__44763\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__44763\,
            I => \N__44760\
        );

    \I__9515\ : Odrv4
    port map (
            O => \N__44760\,
            I => n9
        );

    \I__9514\ : InMux
    port map (
            O => \N__44757\,
            I => \N__44753\
        );

    \I__9513\ : InMux
    port map (
            O => \N__44756\,
            I => \N__44750\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__44753\,
            I => \N__44745\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__44750\,
            I => \N__44745\
        );

    \I__9510\ : Span4Mux_v
    port map (
            O => \N__44745\,
            I => \N__44741\
        );

    \I__9509\ : InMux
    port map (
            O => \N__44744\,
            I => \N__44738\
        );

    \I__9508\ : Sp12to4
    port map (
            O => \N__44741\,
            I => \N__44735\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__44738\,
            I => n295
        );

    \I__9506\ : Odrv12
    port map (
            O => \N__44735\,
            I => n295
        );

    \I__9505\ : InMux
    port map (
            O => \N__44730\,
            I => \N__44723\
        );

    \I__9504\ : InMux
    port map (
            O => \N__44729\,
            I => \N__44723\
        );

    \I__9503\ : CascadeMux
    port map (
            O => \N__44728\,
            I => \N__44720\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__44723\,
            I => \N__44717\
        );

    \I__9501\ : InMux
    port map (
            O => \N__44720\,
            I => \N__44714\
        );

    \I__9500\ : Span4Mux_h
    port map (
            O => \N__44717\,
            I => \N__44711\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__44714\,
            I => encoder0_position_24
        );

    \I__9498\ : Odrv4
    port map (
            O => \N__44711\,
            I => encoder0_position_24
        );

    \I__9497\ : CascadeMux
    port map (
            O => \N__44706\,
            I => \N__44703\
        );

    \I__9496\ : InMux
    port map (
            O => \N__44703\,
            I => \N__44700\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__44700\,
            I => \N__44697\
        );

    \I__9494\ : Span4Mux_h
    port map (
            O => \N__44697\,
            I => \N__44694\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__44694\,
            I => n9_adj_630
        );

    \I__9492\ : InMux
    port map (
            O => \N__44691\,
            I => \N__44688\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__44688\,
            I => \N__44684\
        );

    \I__9490\ : CascadeMux
    port map (
            O => \N__44687\,
            I => \N__44681\
        );

    \I__9489\ : Span4Mux_v
    port map (
            O => \N__44684\,
            I => \N__44677\
        );

    \I__9488\ : InMux
    port map (
            O => \N__44681\,
            I => \N__44674\
        );

    \I__9487\ : InMux
    port map (
            O => \N__44680\,
            I => \N__44671\
        );

    \I__9486\ : Odrv4
    port map (
            O => \N__44677\,
            I => n933
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__44674\,
            I => n933
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__44671\,
            I => n933
        );

    \I__9483\ : CascadeMux
    port map (
            O => \N__44664\,
            I => \N__44661\
        );

    \I__9482\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44658\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__44658\,
            I => n1000
        );

    \I__9480\ : CascadeMux
    port map (
            O => \N__44655\,
            I => \n1032_cascade_\
        );

    \I__9479\ : CascadeMux
    port map (
            O => \N__44652\,
            I => \n11914_cascade_\
        );

    \I__9478\ : InMux
    port map (
            O => \N__44649\,
            I => n12556
        );

    \I__9477\ : InMux
    port map (
            O => \N__44646\,
            I => \bfn_13_20_0_\
        );

    \I__9476\ : InMux
    port map (
            O => \N__44643\,
            I => n12558
        );

    \I__9475\ : InMux
    port map (
            O => \N__44640\,
            I => \N__44637\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__44637\,
            I => n1591
        );

    \I__9473\ : InMux
    port map (
            O => \N__44634\,
            I => n12559
        );

    \I__9472\ : InMux
    port map (
            O => \N__44631\,
            I => n12560
        );

    \I__9471\ : InMux
    port map (
            O => \N__44628\,
            I => n12561
        );

    \I__9470\ : InMux
    port map (
            O => \N__44625\,
            I => n12562
        );

    \I__9469\ : InMux
    port map (
            O => \N__44622\,
            I => \N__44619\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__44619\,
            I => \N__44616\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__44616\,
            I => \N__44613\
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__44613\,
            I => n13
        );

    \I__9465\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44607\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__44607\,
            I => \N__44602\
        );

    \I__9463\ : InMux
    port map (
            O => \N__44606\,
            I => \N__44599\
        );

    \I__9462\ : InMux
    port map (
            O => \N__44605\,
            I => \N__44596\
        );

    \I__9461\ : Span4Mux_v
    port map (
            O => \N__44602\,
            I => \N__44593\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__44599\,
            I => \N__44590\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__44596\,
            I => encoder0_position_20
        );

    \I__9458\ : Odrv4
    port map (
            O => \N__44593\,
            I => encoder0_position_20
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__44590\,
            I => encoder0_position_20
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__44583\,
            I => \N__44580\
        );

    \I__9455\ : InMux
    port map (
            O => \N__44580\,
            I => \N__44575\
        );

    \I__9454\ : InMux
    port map (
            O => \N__44579\,
            I => \N__44572\
        );

    \I__9453\ : InMux
    port map (
            O => \N__44578\,
            I => \N__44569\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__44575\,
            I => n1720
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__44572\,
            I => n1720
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__44569\,
            I => n1720
        );

    \I__9449\ : InMux
    port map (
            O => \N__44562\,
            I => \N__44559\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__44559\,
            I => \N__44556\
        );

    \I__9447\ : Odrv4
    port map (
            O => \N__44556\,
            I => n1787
        );

    \I__9446\ : InMux
    port map (
            O => \N__44553\,
            I => n12590
        );

    \I__9445\ : InMux
    port map (
            O => \N__44550\,
            I => \N__44547\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__44547\,
            I => \N__44544\
        );

    \I__9443\ : Span4Mux_v
    port map (
            O => \N__44544\,
            I => \N__44540\
        );

    \I__9442\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44537\
        );

    \I__9441\ : Span4Mux_h
    port map (
            O => \N__44540\,
            I => \N__44534\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__44537\,
            I => \N__44531\
        );

    \I__9439\ : Odrv4
    port map (
            O => \N__44534\,
            I => n15622
        );

    \I__9438\ : Odrv4
    port map (
            O => \N__44531\,
            I => n15622
        );

    \I__9437\ : InMux
    port map (
            O => \N__44526\,
            I => n12591
        );

    \I__9436\ : InMux
    port map (
            O => \N__44523\,
            I => \N__44520\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__44520\,
            I => \N__44515\
        );

    \I__9434\ : InMux
    port map (
            O => \N__44519\,
            I => \N__44512\
        );

    \I__9433\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44509\
        );

    \I__9432\ : Span4Mux_v
    port map (
            O => \N__44515\,
            I => \N__44504\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__44512\,
            I => \N__44504\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__44509\,
            I => n1818
        );

    \I__9429\ : Odrv4
    port map (
            O => \N__44504\,
            I => n1818
        );

    \I__9428\ : InMux
    port map (
            O => \N__44499\,
            I => \bfn_13_19_0_\
        );

    \I__9427\ : InMux
    port map (
            O => \N__44496\,
            I => n12550
        );

    \I__9426\ : InMux
    port map (
            O => \N__44493\,
            I => n12551
        );

    \I__9425\ : InMux
    port map (
            O => \N__44490\,
            I => n12552
        );

    \I__9424\ : InMux
    port map (
            O => \N__44487\,
            I => n12553
        );

    \I__9423\ : InMux
    port map (
            O => \N__44484\,
            I => n12554
        );

    \I__9422\ : InMux
    port map (
            O => \N__44481\,
            I => n12555
        );

    \I__9421\ : InMux
    port map (
            O => \N__44478\,
            I => \N__44475\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__44475\,
            I => \N__44472\
        );

    \I__9419\ : Odrv4
    port map (
            O => \N__44472\,
            I => n1795
        );

    \I__9418\ : InMux
    port map (
            O => \N__44469\,
            I => n12582
        );

    \I__9417\ : CascadeMux
    port map (
            O => \N__44466\,
            I => \N__44463\
        );

    \I__9416\ : InMux
    port map (
            O => \N__44463\,
            I => \N__44460\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__44460\,
            I => \N__44457\
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__44457\,
            I => n1794
        );

    \I__9413\ : InMux
    port map (
            O => \N__44454\,
            I => n12583
        );

    \I__9412\ : InMux
    port map (
            O => \N__44451\,
            I => \N__44448\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__44448\,
            I => \N__44445\
        );

    \I__9410\ : Odrv4
    port map (
            O => \N__44445\,
            I => n1793
        );

    \I__9409\ : InMux
    port map (
            O => \N__44442\,
            I => \bfn_13_18_0_\
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__44439\,
            I => \N__44436\
        );

    \I__9407\ : InMux
    port map (
            O => \N__44436\,
            I => \N__44433\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__44433\,
            I => \N__44430\
        );

    \I__9405\ : Odrv4
    port map (
            O => \N__44430\,
            I => n1792
        );

    \I__9404\ : InMux
    port map (
            O => \N__44427\,
            I => n12585
        );

    \I__9403\ : InMux
    port map (
            O => \N__44424\,
            I => \N__44421\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__44421\,
            I => \N__44418\
        );

    \I__9401\ : Odrv4
    port map (
            O => \N__44418\,
            I => n1791
        );

    \I__9400\ : InMux
    port map (
            O => \N__44415\,
            I => n12586
        );

    \I__9399\ : InMux
    port map (
            O => \N__44412\,
            I => \N__44409\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__44409\,
            I => \N__44406\
        );

    \I__9397\ : Span4Mux_v
    port map (
            O => \N__44406\,
            I => \N__44403\
        );

    \I__9396\ : Odrv4
    port map (
            O => \N__44403\,
            I => n1790
        );

    \I__9395\ : InMux
    port map (
            O => \N__44400\,
            I => n12587
        );

    \I__9394\ : CascadeMux
    port map (
            O => \N__44397\,
            I => \N__44394\
        );

    \I__9393\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44390\
        );

    \I__9392\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44387\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__44390\,
            I => n1722
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__44387\,
            I => n1722
        );

    \I__9389\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44379\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__44379\,
            I => n1789
        );

    \I__9387\ : InMux
    port map (
            O => \N__44376\,
            I => n12588
        );

    \I__9386\ : InMux
    port map (
            O => \N__44373\,
            I => \N__44368\
        );

    \I__9385\ : InMux
    port map (
            O => \N__44372\,
            I => \N__44365\
        );

    \I__9384\ : InMux
    port map (
            O => \N__44371\,
            I => \N__44362\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__44368\,
            I => n1721
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__44365\,
            I => n1721
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__44362\,
            I => n1721
        );

    \I__9380\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44352\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__44352\,
            I => \N__44349\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__44349\,
            I => \N__44346\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__44346\,
            I => n1788
        );

    \I__9376\ : InMux
    port map (
            O => \N__44343\,
            I => n12589
        );

    \I__9375\ : SRMux
    port map (
            O => \N__44340\,
            I => \N__44336\
        );

    \I__9374\ : InMux
    port map (
            O => \N__44339\,
            I => \N__44333\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__44336\,
            I => \N__44330\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__44333\,
            I => \N__44327\
        );

    \I__9371\ : Odrv12
    port map (
            O => \N__44330\,
            I => \pwm_setpoint_23__N_195\
        );

    \I__9370\ : Odrv4
    port map (
            O => \N__44327\,
            I => \pwm_setpoint_23__N_195\
        );

    \I__9369\ : InMux
    port map (
            O => \N__44322\,
            I => \N__44319\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__44319\,
            I => \N__44316\
        );

    \I__9367\ : Odrv12
    port map (
            O => \N__44316\,
            I => \pwm_setpoint_23_N_171_21\
        );

    \I__9366\ : InMux
    port map (
            O => \N__44313\,
            I => \N__44307\
        );

    \I__9365\ : InMux
    port map (
            O => \N__44312\,
            I => \N__44307\
        );

    \I__9364\ : LocalMux
    port map (
            O => \N__44307\,
            I => \N__44304\
        );

    \I__9363\ : Odrv12
    port map (
            O => \N__44304\,
            I => duty_21
        );

    \I__9362\ : InMux
    port map (
            O => \N__44301\,
            I => \N__44298\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__44298\,
            I => \N__44295\
        );

    \I__9360\ : Span4Mux_v
    port map (
            O => \N__44295\,
            I => \N__44292\
        );

    \I__9359\ : Span4Mux_h
    port map (
            O => \N__44292\,
            I => \N__44289\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__44289\,
            I => n1801
        );

    \I__9357\ : InMux
    port map (
            O => \N__44286\,
            I => \bfn_13_17_0_\
        );

    \I__9356\ : CascadeMux
    port map (
            O => \N__44283\,
            I => \N__44280\
        );

    \I__9355\ : InMux
    port map (
            O => \N__44280\,
            I => \N__44277\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__44277\,
            I => \N__44274\
        );

    \I__9353\ : Span4Mux_v
    port map (
            O => \N__44274\,
            I => \N__44271\
        );

    \I__9352\ : Odrv4
    port map (
            O => \N__44271\,
            I => n1800
        );

    \I__9351\ : InMux
    port map (
            O => \N__44268\,
            I => n12577
        );

    \I__9350\ : InMux
    port map (
            O => \N__44265\,
            I => \N__44262\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__44262\,
            I => \N__44259\
        );

    \I__9348\ : Span4Mux_v
    port map (
            O => \N__44259\,
            I => \N__44256\
        );

    \I__9347\ : Odrv4
    port map (
            O => \N__44256\,
            I => n1799
        );

    \I__9346\ : InMux
    port map (
            O => \N__44253\,
            I => n12578
        );

    \I__9345\ : InMux
    port map (
            O => \N__44250\,
            I => \N__44247\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__44247\,
            I => \N__44244\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__44244\,
            I => n1798
        );

    \I__9342\ : InMux
    port map (
            O => \N__44241\,
            I => n12579
        );

    \I__9341\ : InMux
    port map (
            O => \N__44238\,
            I => \N__44235\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__9339\ : Odrv4
    port map (
            O => \N__44232\,
            I => n1797
        );

    \I__9338\ : InMux
    port map (
            O => \N__44229\,
            I => n12580
        );

    \I__9337\ : CascadeMux
    port map (
            O => \N__44226\,
            I => \N__44223\
        );

    \I__9336\ : InMux
    port map (
            O => \N__44223\,
            I => \N__44220\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__44220\,
            I => \N__44217\
        );

    \I__9334\ : Span4Mux_v
    port map (
            O => \N__44217\,
            I => \N__44214\
        );

    \I__9333\ : Odrv4
    port map (
            O => \N__44214\,
            I => n1796
        );

    \I__9332\ : InMux
    port map (
            O => \N__44211\,
            I => n12581
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__44208\,
            I => \n8_adj_657_cascade_\
        );

    \I__9330\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44202\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__44202\,
            I => \N__44199\
        );

    \I__9328\ : Odrv12
    port map (
            O => \N__44199\,
            I => n15180
        );

    \I__9327\ : CascadeMux
    port map (
            O => \N__44196\,
            I => \n15219_cascade_\
        );

    \I__9326\ : InMux
    port map (
            O => \N__44193\,
            I => \N__44190\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__44190\,
            I => n24_adj_669
        );

    \I__9324\ : InMux
    port map (
            O => \N__44187\,
            I => \N__44181\
        );

    \I__9323\ : InMux
    port map (
            O => \N__44186\,
            I => \N__44181\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__44181\,
            I => \N__44178\
        );

    \I__9321\ : Span4Mux_h
    port map (
            O => \N__44178\,
            I => \N__44175\
        );

    \I__9320\ : Odrv4
    port map (
            O => \N__44175\,
            I => pwm_setpoint_22
        );

    \I__9319\ : InMux
    port map (
            O => \N__44172\,
            I => \N__44169\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__44169\,
            I => n15274
        );

    \I__9317\ : InMux
    port map (
            O => \N__44166\,
            I => \N__44160\
        );

    \I__9316\ : InMux
    port map (
            O => \N__44165\,
            I => \N__44153\
        );

    \I__9315\ : InMux
    port map (
            O => \N__44164\,
            I => \N__44153\
        );

    \I__9314\ : InMux
    port map (
            O => \N__44163\,
            I => \N__44153\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__44160\,
            I => n45
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__44153\,
            I => n45
        );

    \I__9311\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44145\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__44145\,
            I => n15255
        );

    \I__9309\ : CascadeMux
    port map (
            O => \N__44142\,
            I => \n40_cascade_\
        );

    \I__9308\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44135\
        );

    \I__9307\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44132\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__44135\,
            I => \N__44127\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__44132\,
            I => \N__44127\
        );

    \I__9304\ : Span4Mux_s2_v
    port map (
            O => \N__44127\,
            I => \N__44124\
        );

    \I__9303\ : Odrv4
    port map (
            O => \N__44124\,
            I => duty_20
        );

    \I__9302\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44118\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__44118\,
            I => \N__44115\
        );

    \I__9300\ : Odrv4
    port map (
            O => \N__44115\,
            I => \pwm_setpoint_23_N_171_20\
        );

    \I__9299\ : CascadeMux
    port map (
            O => \N__44112\,
            I => \N__44109\
        );

    \I__9298\ : InMux
    port map (
            O => \N__44109\,
            I => \N__44106\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__44106\,
            I => \N__44103\
        );

    \I__9296\ : Odrv12
    port map (
            O => \N__44103\,
            I => n4_adj_584
        );

    \I__9295\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44097\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__44097\,
            I => n16_adj_664
        );

    \I__9293\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44090\
        );

    \I__9292\ : InMux
    port map (
            O => \N__44093\,
            I => \N__44087\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__44090\,
            I => \N__44084\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__44087\,
            I => \N__44079\
        );

    \I__9289\ : Span4Mux_h
    port map (
            O => \N__44084\,
            I => \N__44079\
        );

    \I__9288\ : Odrv4
    port map (
            O => \N__44079\,
            I => duty_12
        );

    \I__9287\ : InMux
    port map (
            O => \N__44076\,
            I => \N__44073\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__44073\,
            I => \N__44070\
        );

    \I__9285\ : Span4Mux_h
    port map (
            O => \N__44070\,
            I => \N__44067\
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__44067\,
            I => \pwm_setpoint_23_N_171_12\
        );

    \I__9283\ : InMux
    port map (
            O => \N__44064\,
            I => \N__44058\
        );

    \I__9282\ : InMux
    port map (
            O => \N__44063\,
            I => \N__44058\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__44058\,
            I => n37
        );

    \I__9280\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44051\
        );

    \I__9279\ : InMux
    port map (
            O => \N__44054\,
            I => \N__44048\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__44051\,
            I => \N__44045\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__44048\,
            I => \N__44042\
        );

    \I__9276\ : Span4Mux_h
    port map (
            O => \N__44045\,
            I => \N__44039\
        );

    \I__9275\ : Span4Mux_h
    port map (
            O => \N__44042\,
            I => \N__44036\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__44039\,
            I => pwm_setpoint_18
        );

    \I__9273\ : Odrv4
    port map (
            O => \N__44036\,
            I => pwm_setpoint_18
        );

    \I__9272\ : InMux
    port map (
            O => \N__44031\,
            I => \N__44028\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__44028\,
            I => \N__44025\
        );

    \I__9270\ : Odrv4
    port map (
            O => \N__44025\,
            I => n15277
        );

    \I__9269\ : InMux
    port map (
            O => \N__44022\,
            I => \N__44019\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__44019\,
            I => \N__44016\
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__44016\,
            I => n6_adj_656
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__44013\,
            I => \n15235_cascade_\
        );

    \I__9265\ : CascadeMux
    port map (
            O => \N__44010\,
            I => \n15236_cascade_\
        );

    \I__9264\ : InMux
    port map (
            O => \N__44007\,
            I => \N__44003\
        );

    \I__9263\ : InMux
    port map (
            O => \N__44006\,
            I => \N__44000\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__44003\,
            I => \N__43997\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__44000\,
            I => \N__43994\
        );

    \I__9260\ : Span4Mux_v
    port map (
            O => \N__43997\,
            I => \N__43991\
        );

    \I__9259\ : Odrv4
    port map (
            O => \N__43994\,
            I => duty_11
        );

    \I__9258\ : Odrv4
    port map (
            O => \N__43991\,
            I => duty_11
        );

    \I__9257\ : InMux
    port map (
            O => \N__43986\,
            I => \N__43983\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__43983\,
            I => \N__43980\
        );

    \I__9255\ : Span4Mux_v
    port map (
            O => \N__43980\,
            I => \N__43977\
        );

    \I__9254\ : Odrv4
    port map (
            O => \N__43977\,
            I => \pwm_setpoint_23_N_171_11\
        );

    \I__9253\ : InMux
    port map (
            O => \N__43974\,
            I => \N__43970\
        );

    \I__9252\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43967\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__43970\,
            I => \N__43964\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__43967\,
            I => \N__43961\
        );

    \I__9249\ : Span4Mux_s2_v
    port map (
            O => \N__43964\,
            I => \N__43958\
        );

    \I__9248\ : Odrv4
    port map (
            O => \N__43961\,
            I => duty_17
        );

    \I__9247\ : Odrv4
    port map (
            O => \N__43958\,
            I => duty_17
        );

    \I__9246\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43950\
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__43950\,
            I => \N__43947\
        );

    \I__9244\ : Span4Mux_h
    port map (
            O => \N__43947\,
            I => \N__43944\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__43944\,
            I => \pwm_setpoint_23_N_171_17\
        );

    \I__9242\ : InMux
    port map (
            O => \N__43941\,
            I => \N__43938\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__43938\,
            I => \N__43935\
        );

    \I__9240\ : Span4Mux_h
    port map (
            O => \N__43935\,
            I => \N__43931\
        );

    \I__9239\ : InMux
    port map (
            O => \N__43934\,
            I => \N__43928\
        );

    \I__9238\ : Odrv4
    port map (
            O => \N__43931\,
            I => pwm_setpoint_17
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__43928\,
            I => pwm_setpoint_17
        );

    \I__9236\ : InMux
    port map (
            O => \N__43923\,
            I => \N__43920\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__43920\,
            I => n15278
        );

    \I__9234\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43914\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__43914\,
            I => \N__43911\
        );

    \I__9232\ : Odrv12
    port map (
            O => \N__43911\,
            I => n6_adj_577
        );

    \I__9231\ : InMux
    port map (
            O => \N__43908\,
            I => \N__43904\
        );

    \I__9230\ : InMux
    port map (
            O => \N__43907\,
            I => \N__43901\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__43904\,
            I => \N__43898\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__43901\,
            I => \N__43895\
        );

    \I__9227\ : Span4Mux_s3_v
    port map (
            O => \N__43898\,
            I => \N__43890\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__43895\,
            I => \N__43890\
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__43890\,
            I => duty_19
        );

    \I__9224\ : InMux
    port map (
            O => \N__43887\,
            I => n12477
        );

    \I__9223\ : CascadeMux
    port map (
            O => \N__43884\,
            I => \N__43881\
        );

    \I__9222\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__43878\,
            I => n5_adj_578
        );

    \I__9220\ : InMux
    port map (
            O => \N__43875\,
            I => n12478
        );

    \I__9219\ : InMux
    port map (
            O => \N__43872\,
            I => \N__43869\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__43869\,
            I => \N__43866\
        );

    \I__9217\ : Odrv12
    port map (
            O => \N__43866\,
            I => n4_adj_579
        );

    \I__9216\ : InMux
    port map (
            O => \N__43863\,
            I => n12479
        );

    \I__9215\ : InMux
    port map (
            O => \N__43860\,
            I => \N__43857\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__43857\,
            I => \N__43854\
        );

    \I__9213\ : Span4Mux_v
    port map (
            O => \N__43854\,
            I => \N__43851\
        );

    \I__9212\ : Odrv4
    port map (
            O => \N__43851\,
            I => n3_adj_580
        );

    \I__9211\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43842\
        );

    \I__9210\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43842\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__43842\,
            I => \N__43839\
        );

    \I__9208\ : Span12Mux_s4_v
    port map (
            O => \N__43839\,
            I => \N__43836\
        );

    \I__9207\ : Odrv12
    port map (
            O => \N__43836\,
            I => duty_22
        );

    \I__9206\ : InMux
    port map (
            O => \N__43833\,
            I => n12480
        );

    \I__9205\ : InMux
    port map (
            O => \N__43830\,
            I => \N__43827\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__43827\,
            I => n2_adj_581
        );

    \I__9203\ : InMux
    port map (
            O => \N__43824\,
            I => n12481
        );

    \I__9202\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43812\
        );

    \I__9201\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43812\
        );

    \I__9200\ : InMux
    port map (
            O => \N__43819\,
            I => \N__43812\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__43812\,
            I => \N__43809\
        );

    \I__9198\ : Odrv4
    port map (
            O => \N__43809\,
            I => n35
        );

    \I__9197\ : InMux
    port map (
            O => \N__43806\,
            I => \N__43803\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__43803\,
            I => \N__43800\
        );

    \I__9195\ : Span4Mux_h
    port map (
            O => \N__43800\,
            I => \N__43797\
        );

    \I__9194\ : Odrv4
    port map (
            O => \N__43797\,
            I => n33_adj_675
        );

    \I__9193\ : CascadeMux
    port map (
            O => \N__43794\,
            I => \n35_cascade_\
        );

    \I__9192\ : InMux
    port map (
            O => \N__43791\,
            I => \N__43788\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__43788\,
            I => \N__43785\
        );

    \I__9190\ : Odrv12
    port map (
            O => \N__43785\,
            I => n15225
        );

    \I__9189\ : InMux
    port map (
            O => \N__43782\,
            I => \N__43778\
        );

    \I__9188\ : InMux
    port map (
            O => \N__43781\,
            I => \N__43775\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__43778\,
            I => \N__43772\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__43775\,
            I => pwm_setpoint_13
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__43772\,
            I => pwm_setpoint_13
        );

    \I__9184\ : CascadeMux
    port map (
            O => \N__43767\,
            I => \N__43764\
        );

    \I__9183\ : InMux
    port map (
            O => \N__43764\,
            I => \N__43759\
        );

    \I__9182\ : InMux
    port map (
            O => \N__43763\,
            I => \N__43756\
        );

    \I__9181\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43753\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__43759\,
            I => \N__43750\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__43756\,
            I => \N__43745\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__43753\,
            I => \N__43745\
        );

    \I__9177\ : Sp12to4
    port map (
            O => \N__43750\,
            I => \N__43742\
        );

    \I__9176\ : Span4Mux_h
    port map (
            O => \N__43745\,
            I => \N__43739\
        );

    \I__9175\ : Odrv12
    port map (
            O => \N__43742\,
            I => n27_adj_671
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__43739\,
            I => n27_adj_671
        );

    \I__9173\ : InMux
    port map (
            O => \N__43734\,
            I => \N__43731\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__43731\,
            I => n14_adj_569
        );

    \I__9171\ : InMux
    port map (
            O => \N__43728\,
            I => n12469
        );

    \I__9170\ : InMux
    port map (
            O => \N__43725\,
            I => \N__43722\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__43722\,
            I => \N__43719\
        );

    \I__9168\ : Odrv12
    port map (
            O => \N__43719\,
            I => n13_adj_570
        );

    \I__9167\ : InMux
    port map (
            O => \N__43716\,
            I => n12470
        );

    \I__9166\ : InMux
    port map (
            O => \N__43713\,
            I => \N__43710\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__43710\,
            I => \N__43707\
        );

    \I__9164\ : Span4Mux_v
    port map (
            O => \N__43707\,
            I => \N__43704\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__43704\,
            I => n12_adj_571
        );

    \I__9162\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43698\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__43698\,
            I => \N__43694\
        );

    \I__9160\ : InMux
    port map (
            O => \N__43697\,
            I => \N__43691\
        );

    \I__9159\ : Span4Mux_v
    port map (
            O => \N__43694\,
            I => \N__43688\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__43691\,
            I => duty_13
        );

    \I__9157\ : Odrv4
    port map (
            O => \N__43688\,
            I => duty_13
        );

    \I__9156\ : InMux
    port map (
            O => \N__43683\,
            I => n12471
        );

    \I__9155\ : InMux
    port map (
            O => \N__43680\,
            I => \N__43677\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__43677\,
            I => n11_adj_572
        );

    \I__9153\ : InMux
    port map (
            O => \N__43674\,
            I => \N__43670\
        );

    \I__9152\ : InMux
    port map (
            O => \N__43673\,
            I => \N__43667\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__43670\,
            I => \N__43662\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__43667\,
            I => \N__43662\
        );

    \I__9149\ : Span4Mux_v
    port map (
            O => \N__43662\,
            I => \N__43659\
        );

    \I__9148\ : Odrv4
    port map (
            O => \N__43659\,
            I => duty_14
        );

    \I__9147\ : InMux
    port map (
            O => \N__43656\,
            I => n12472
        );

    \I__9146\ : CascadeMux
    port map (
            O => \N__43653\,
            I => \N__43650\
        );

    \I__9145\ : InMux
    port map (
            O => \N__43650\,
            I => \N__43647\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__43647\,
            I => \N__43644\
        );

    \I__9143\ : Span4Mux_v
    port map (
            O => \N__43644\,
            I => \N__43641\
        );

    \I__9142\ : Sp12to4
    port map (
            O => \N__43641\,
            I => \N__43638\
        );

    \I__9141\ : Odrv12
    port map (
            O => \N__43638\,
            I => n10_adj_573
        );

    \I__9140\ : InMux
    port map (
            O => \N__43635\,
            I => \N__43631\
        );

    \I__9139\ : InMux
    port map (
            O => \N__43634\,
            I => \N__43628\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__43631\,
            I => \N__43625\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__43628\,
            I => \N__43622\
        );

    \I__9136\ : Span4Mux_v
    port map (
            O => \N__43625\,
            I => \N__43619\
        );

    \I__9135\ : Span4Mux_h
    port map (
            O => \N__43622\,
            I => \N__43616\
        );

    \I__9134\ : Odrv4
    port map (
            O => \N__43619\,
            I => duty_15
        );

    \I__9133\ : Odrv4
    port map (
            O => \N__43616\,
            I => duty_15
        );

    \I__9132\ : InMux
    port map (
            O => \N__43611\,
            I => n12473
        );

    \I__9131\ : InMux
    port map (
            O => \N__43608\,
            I => \N__43605\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__43605\,
            I => \N__43602\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__43602\,
            I => n9_adj_574
        );

    \I__9128\ : InMux
    port map (
            O => \N__43599\,
            I => \N__43595\
        );

    \I__9127\ : InMux
    port map (
            O => \N__43598\,
            I => \N__43592\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__43595\,
            I => \N__43589\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__43592\,
            I => \N__43586\
        );

    \I__9124\ : Span4Mux_h
    port map (
            O => \N__43589\,
            I => \N__43581\
        );

    \I__9123\ : Span4Mux_v
    port map (
            O => \N__43586\,
            I => \N__43581\
        );

    \I__9122\ : Odrv4
    port map (
            O => \N__43581\,
            I => duty_16
        );

    \I__9121\ : InMux
    port map (
            O => \N__43578\,
            I => \bfn_12_28_0_\
        );

    \I__9120\ : InMux
    port map (
            O => \N__43575\,
            I => \N__43572\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__43572\,
            I => \N__43569\
        );

    \I__9118\ : Span4Mux_h
    port map (
            O => \N__43569\,
            I => \N__43566\
        );

    \I__9117\ : Odrv4
    port map (
            O => \N__43566\,
            I => n8_adj_575
        );

    \I__9116\ : InMux
    port map (
            O => \N__43563\,
            I => n12475
        );

    \I__9115\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43557\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__43557\,
            I => n7_adj_576
        );

    \I__9113\ : InMux
    port map (
            O => \N__43554\,
            I => \N__43550\
        );

    \I__9112\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43547\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__43550\,
            I => \N__43544\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__43547\,
            I => \N__43541\
        );

    \I__9109\ : Span4Mux_v
    port map (
            O => \N__43544\,
            I => \N__43538\
        );

    \I__9108\ : Span4Mux_h
    port map (
            O => \N__43541\,
            I => \N__43535\
        );

    \I__9107\ : Odrv4
    port map (
            O => \N__43538\,
            I => duty_18
        );

    \I__9106\ : Odrv4
    port map (
            O => \N__43535\,
            I => duty_18
        );

    \I__9105\ : InMux
    port map (
            O => \N__43530\,
            I => n12476
        );

    \I__9104\ : InMux
    port map (
            O => \N__43527\,
            I => \N__43524\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__43524\,
            I => \N__43521\
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__43521\,
            I => n22_adj_555
        );

    \I__9101\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43515\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__43515\,
            I => \N__43511\
        );

    \I__9099\ : InMux
    port map (
            O => \N__43514\,
            I => \N__43508\
        );

    \I__9098\ : Span4Mux_h
    port map (
            O => \N__43511\,
            I => \N__43505\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__43508\,
            I => duty_3
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__43505\,
            I => duty_3
        );

    \I__9095\ : InMux
    port map (
            O => \N__43500\,
            I => n12461
        );

    \I__9094\ : CascadeMux
    port map (
            O => \N__43497\,
            I => \N__43494\
        );

    \I__9093\ : InMux
    port map (
            O => \N__43494\,
            I => \N__43491\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__43491\,
            I => \N__43488\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__43488\,
            I => n21_adj_556
        );

    \I__9090\ : InMux
    port map (
            O => \N__43485\,
            I => \N__43482\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__43482\,
            I => \N__43479\
        );

    \I__9088\ : Span4Mux_s2_v
    port map (
            O => \N__43479\,
            I => \N__43475\
        );

    \I__9087\ : InMux
    port map (
            O => \N__43478\,
            I => \N__43472\
        );

    \I__9086\ : Sp12to4
    port map (
            O => \N__43475\,
            I => \N__43467\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__43472\,
            I => \N__43467\
        );

    \I__9084\ : Span12Mux_s11_h
    port map (
            O => \N__43467\,
            I => \N__43464\
        );

    \I__9083\ : Odrv12
    port map (
            O => \N__43464\,
            I => duty_4
        );

    \I__9082\ : InMux
    port map (
            O => \N__43461\,
            I => n12462
        );

    \I__9081\ : InMux
    port map (
            O => \N__43458\,
            I => \N__43455\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__43455\,
            I => \N__43452\
        );

    \I__9079\ : Odrv12
    port map (
            O => \N__43452\,
            I => n20_adj_557
        );

    \I__9078\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43443\
        );

    \I__9077\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43443\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__43443\,
            I => \N__43440\
        );

    \I__9075\ : Span4Mux_v
    port map (
            O => \N__43440\,
            I => \N__43437\
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__43437\,
            I => duty_5
        );

    \I__9073\ : InMux
    port map (
            O => \N__43434\,
            I => n12463
        );

    \I__9072\ : InMux
    port map (
            O => \N__43431\,
            I => \N__43428\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__43428\,
            I => n19_adj_558
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__43425\,
            I => \N__43422\
        );

    \I__9069\ : InMux
    port map (
            O => \N__43422\,
            I => \N__43416\
        );

    \I__9068\ : InMux
    port map (
            O => \N__43421\,
            I => \N__43416\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__43416\,
            I => \N__43413\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__43413\,
            I => \N__43410\
        );

    \I__9065\ : Odrv4
    port map (
            O => \N__43410\,
            I => duty_6
        );

    \I__9064\ : InMux
    port map (
            O => \N__43407\,
            I => n12464
        );

    \I__9063\ : CascadeMux
    port map (
            O => \N__43404\,
            I => \N__43401\
        );

    \I__9062\ : InMux
    port map (
            O => \N__43401\,
            I => \N__43398\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__43398\,
            I => \N__43395\
        );

    \I__9060\ : Odrv12
    port map (
            O => \N__43395\,
            I => n18_adj_559
        );

    \I__9059\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43388\
        );

    \I__9058\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43385\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__43388\,
            I => \N__43382\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__43385\,
            I => \N__43377\
        );

    \I__9055\ : Span4Mux_h
    port map (
            O => \N__43382\,
            I => \N__43377\
        );

    \I__9054\ : Odrv4
    port map (
            O => \N__43377\,
            I => duty_7
        );

    \I__9053\ : InMux
    port map (
            O => \N__43374\,
            I => n12465
        );

    \I__9052\ : InMux
    port map (
            O => \N__43371\,
            I => \N__43368\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__43368\,
            I => \N__43365\
        );

    \I__9050\ : Odrv12
    port map (
            O => \N__43365\,
            I => n17_adj_560
        );

    \I__9049\ : InMux
    port map (
            O => \N__43362\,
            I => \bfn_12_27_0_\
        );

    \I__9048\ : InMux
    port map (
            O => \N__43359\,
            I => \N__43356\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__43356\,
            I => n16_adj_563
        );

    \I__9046\ : InMux
    port map (
            O => \N__43353\,
            I => \N__43349\
        );

    \I__9045\ : InMux
    port map (
            O => \N__43352\,
            I => \N__43346\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__43349\,
            I => \N__43341\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__43346\,
            I => \N__43341\
        );

    \I__9042\ : Span4Mux_v
    port map (
            O => \N__43341\,
            I => \N__43338\
        );

    \I__9041\ : Odrv4
    port map (
            O => \N__43338\,
            I => duty_9
        );

    \I__9040\ : InMux
    port map (
            O => \N__43335\,
            I => n12467
        );

    \I__9039\ : InMux
    port map (
            O => \N__43332\,
            I => \N__43329\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__43329\,
            I => n15_adj_568
        );

    \I__9037\ : InMux
    port map (
            O => \N__43326\,
            I => \N__43320\
        );

    \I__9036\ : InMux
    port map (
            O => \N__43325\,
            I => \N__43320\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__43320\,
            I => \N__43317\
        );

    \I__9034\ : Span4Mux_h
    port map (
            O => \N__43317\,
            I => \N__43314\
        );

    \I__9033\ : Odrv4
    port map (
            O => \N__43314\,
            I => duty_10
        );

    \I__9032\ : InMux
    port map (
            O => \N__43311\,
            I => n12468
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__43308\,
            I => \N__43305\
        );

    \I__9030\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43302\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__43302\,
            I => n404
        );

    \I__9028\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43296\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__43296\,
            I => n2539
        );

    \I__9026\ : InMux
    port map (
            O => \N__43293\,
            I => n12484
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__43290\,
            I => \N__43287\
        );

    \I__9024\ : InMux
    port map (
            O => \N__43287\,
            I => \N__43284\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__43284\,
            I => \N__43281\
        );

    \I__9022\ : Odrv4
    port map (
            O => \N__43281\,
            I => n403
        );

    \I__9021\ : InMux
    port map (
            O => \N__43278\,
            I => \N__43275\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__43275\,
            I => n2538
        );

    \I__9019\ : InMux
    port map (
            O => \N__43272\,
            I => n12485
        );

    \I__9018\ : CascadeMux
    port map (
            O => \N__43269\,
            I => \N__43266\
        );

    \I__9017\ : InMux
    port map (
            O => \N__43266\,
            I => \N__43263\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__43263\,
            I => \N__43260\
        );

    \I__9015\ : Odrv12
    port map (
            O => \N__43260\,
            I => n402
        );

    \I__9014\ : InMux
    port map (
            O => \N__43257\,
            I => n12486
        );

    \I__9013\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43251\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__43251\,
            I => n2537
        );

    \I__9011\ : InMux
    port map (
            O => \N__43248\,
            I => \N__43245\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__43245\,
            I => \N__43242\
        );

    \I__9009\ : Span4Mux_h
    port map (
            O => \N__43242\,
            I => \N__43239\
        );

    \I__9008\ : Span4Mux_h
    port map (
            O => \N__43239\,
            I => \N__43236\
        );

    \I__9007\ : Odrv4
    port map (
            O => \N__43236\,
            I => encoder0_position_scaled_6
        );

    \I__9006\ : InMux
    port map (
            O => \N__43233\,
            I => \N__43230\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__43230\,
            I => \N__43227\
        );

    \I__9004\ : Span4Mux_h
    port map (
            O => \N__43227\,
            I => \N__43222\
        );

    \I__9003\ : InMux
    port map (
            O => \N__43226\,
            I => \N__43219\
        );

    \I__9002\ : InMux
    port map (
            O => \N__43225\,
            I => \N__43216\
        );

    \I__9001\ : Span4Mux_v
    port map (
            O => \N__43222\,
            I => \N__43213\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__43219\,
            I => \N__43208\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__43216\,
            I => \N__43208\
        );

    \I__8998\ : Span4Mux_h
    port map (
            O => \N__43213\,
            I => \N__43205\
        );

    \I__8997\ : Span4Mux_v
    port map (
            O => \N__43208\,
            I => \N__43202\
        );

    \I__8996\ : Odrv4
    port map (
            O => \N__43205\,
            I => n3109
        );

    \I__8995\ : Odrv4
    port map (
            O => \N__43202\,
            I => n3109
        );

    \I__8994\ : CascadeMux
    port map (
            O => \N__43197\,
            I => \N__43194\
        );

    \I__8993\ : InMux
    port map (
            O => \N__43194\,
            I => \N__43191\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__43191\,
            I => \N__43188\
        );

    \I__8991\ : Span4Mux_v
    port map (
            O => \N__43188\,
            I => \N__43185\
        );

    \I__8990\ : Span4Mux_h
    port map (
            O => \N__43185\,
            I => \N__43182\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__43182\,
            I => n3176
        );

    \I__8988\ : InMux
    port map (
            O => \N__43179\,
            I => \N__43175\
        );

    \I__8987\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43163\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__43175\,
            I => \N__43160\
        );

    \I__8985\ : CascadeMux
    port map (
            O => \N__43174\,
            I => \N__43157\
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__43173\,
            I => \N__43153\
        );

    \I__8983\ : CascadeMux
    port map (
            O => \N__43172\,
            I => \N__43143\
        );

    \I__8982\ : CascadeMux
    port map (
            O => \N__43171\,
            I => \N__43140\
        );

    \I__8981\ : CascadeMux
    port map (
            O => \N__43170\,
            I => \N__43135\
        );

    \I__8980\ : CascadeMux
    port map (
            O => \N__43169\,
            I => \N__43130\
        );

    \I__8979\ : CascadeMux
    port map (
            O => \N__43168\,
            I => \N__43126\
        );

    \I__8978\ : CascadeMux
    port map (
            O => \N__43167\,
            I => \N__43121\
        );

    \I__8977\ : CascadeMux
    port map (
            O => \N__43166\,
            I => \N__43118\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__43163\,
            I => \N__43114\
        );

    \I__8975\ : Span4Mux_h
    port map (
            O => \N__43160\,
            I => \N__43111\
        );

    \I__8974\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43106\
        );

    \I__8973\ : InMux
    port map (
            O => \N__43156\,
            I => \N__43106\
        );

    \I__8972\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43097\
        );

    \I__8971\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43097\
        );

    \I__8970\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43097\
        );

    \I__8969\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43097\
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__43149\,
            I => \N__43094\
        );

    \I__8967\ : CascadeMux
    port map (
            O => \N__43148\,
            I => \N__43090\
        );

    \I__8966\ : CascadeMux
    port map (
            O => \N__43147\,
            I => \N__43087\
        );

    \I__8965\ : InMux
    port map (
            O => \N__43146\,
            I => \N__43082\
        );

    \I__8964\ : InMux
    port map (
            O => \N__43143\,
            I => \N__43073\
        );

    \I__8963\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43073\
        );

    \I__8962\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43073\
        );

    \I__8961\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43073\
        );

    \I__8960\ : InMux
    port map (
            O => \N__43135\,
            I => \N__43066\
        );

    \I__8959\ : InMux
    port map (
            O => \N__43134\,
            I => \N__43066\
        );

    \I__8958\ : InMux
    port map (
            O => \N__43133\,
            I => \N__43066\
        );

    \I__8957\ : InMux
    port map (
            O => \N__43130\,
            I => \N__43057\
        );

    \I__8956\ : InMux
    port map (
            O => \N__43129\,
            I => \N__43057\
        );

    \I__8955\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43057\
        );

    \I__8954\ : InMux
    port map (
            O => \N__43125\,
            I => \N__43057\
        );

    \I__8953\ : InMux
    port map (
            O => \N__43124\,
            I => \N__43048\
        );

    \I__8952\ : InMux
    port map (
            O => \N__43121\,
            I => \N__43048\
        );

    \I__8951\ : InMux
    port map (
            O => \N__43118\,
            I => \N__43048\
        );

    \I__8950\ : InMux
    port map (
            O => \N__43117\,
            I => \N__43048\
        );

    \I__8949\ : Span4Mux_v
    port map (
            O => \N__43114\,
            I => \N__43039\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__43111\,
            I => \N__43039\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__43106\,
            I => \N__43039\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__43097\,
            I => \N__43039\
        );

    \I__8945\ : InMux
    port map (
            O => \N__43094\,
            I => \N__43026\
        );

    \I__8944\ : InMux
    port map (
            O => \N__43093\,
            I => \N__43026\
        );

    \I__8943\ : InMux
    port map (
            O => \N__43090\,
            I => \N__43026\
        );

    \I__8942\ : InMux
    port map (
            O => \N__43087\,
            I => \N__43026\
        );

    \I__8941\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43026\
        );

    \I__8940\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43026\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__43082\,
            I => n3138
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__43073\,
            I => n3138
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__43066\,
            I => n3138
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__43057\,
            I => n3138
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__43048\,
            I => n3138
        );

    \I__8934\ : Odrv4
    port map (
            O => \N__43039\,
            I => n3138
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__43026\,
            I => n3138
        );

    \I__8932\ : InMux
    port map (
            O => \N__43011\,
            I => \N__43007\
        );

    \I__8931\ : CascadeMux
    port map (
            O => \N__43010\,
            I => \N__43003\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__43007\,
            I => \N__43000\
        );

    \I__8929\ : InMux
    port map (
            O => \N__43006\,
            I => \N__42995\
        );

    \I__8928\ : InMux
    port map (
            O => \N__43003\,
            I => \N__42995\
        );

    \I__8927\ : Span4Mux_v
    port map (
            O => \N__43000\,
            I => \N__42992\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__42995\,
            I => \N__42989\
        );

    \I__8925\ : Span4Mux_h
    port map (
            O => \N__42992\,
            I => \N__42986\
        );

    \I__8924\ : Span4Mux_h
    port map (
            O => \N__42989\,
            I => \N__42983\
        );

    \I__8923\ : Odrv4
    port map (
            O => \N__42986\,
            I => n3208
        );

    \I__8922\ : Odrv4
    port map (
            O => \N__42983\,
            I => n3208
        );

    \I__8921\ : InMux
    port map (
            O => \N__42978\,
            I => \N__42975\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__42975\,
            I => \N__42972\
        );

    \I__8919\ : Odrv4
    port map (
            O => \N__42972\,
            I => n25_adj_552
        );

    \I__8918\ : InMux
    port map (
            O => \N__42969\,
            I => \N__42965\
        );

    \I__8917\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42962\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__42965\,
            I => \N__42959\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__42962\,
            I => \N__42956\
        );

    \I__8914\ : Span4Mux_h
    port map (
            O => \N__42959\,
            I => \N__42953\
        );

    \I__8913\ : Odrv12
    port map (
            O => \N__42956\,
            I => duty_0
        );

    \I__8912\ : Odrv4
    port map (
            O => \N__42953\,
            I => duty_0
        );

    \I__8911\ : InMux
    port map (
            O => \N__42948\,
            I => \bfn_12_26_0_\
        );

    \I__8910\ : InMux
    port map (
            O => \N__42945\,
            I => \N__42942\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__42942\,
            I => \N__42939\
        );

    \I__8908\ : Span4Mux_v
    port map (
            O => \N__42939\,
            I => \N__42936\
        );

    \I__8907\ : Odrv4
    port map (
            O => \N__42936\,
            I => n24_adj_553
        );

    \I__8906\ : InMux
    port map (
            O => \N__42933\,
            I => \N__42929\
        );

    \I__8905\ : InMux
    port map (
            O => \N__42932\,
            I => \N__42926\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__42929\,
            I => \N__42923\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__42926\,
            I => \N__42920\
        );

    \I__8902\ : Span4Mux_h
    port map (
            O => \N__42923\,
            I => \N__42917\
        );

    \I__8901\ : Odrv12
    port map (
            O => \N__42920\,
            I => duty_1
        );

    \I__8900\ : Odrv4
    port map (
            O => \N__42917\,
            I => duty_1
        );

    \I__8899\ : InMux
    port map (
            O => \N__42912\,
            I => n12459
        );

    \I__8898\ : CascadeMux
    port map (
            O => \N__42909\,
            I => \N__42906\
        );

    \I__8897\ : InMux
    port map (
            O => \N__42906\,
            I => \N__42903\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__42903\,
            I => \N__42900\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__42900\,
            I => n23_adj_554
        );

    \I__8894\ : InMux
    port map (
            O => \N__42897\,
            I => \N__42893\
        );

    \I__8893\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42890\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__42893\,
            I => \N__42887\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__42890\,
            I => \N__42884\
        );

    \I__8890\ : Span4Mux_v
    port map (
            O => \N__42887\,
            I => \N__42881\
        );

    \I__8889\ : Span4Mux_v
    port map (
            O => \N__42884\,
            I => \N__42878\
        );

    \I__8888\ : Odrv4
    port map (
            O => \N__42881\,
            I => duty_2
        );

    \I__8887\ : Odrv4
    port map (
            O => \N__42878\,
            I => duty_2
        );

    \I__8886\ : InMux
    port map (
            O => \N__42873\,
            I => n12460
        );

    \I__8885\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42867\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__42867\,
            I => \N__42862\
        );

    \I__8883\ : InMux
    port map (
            O => \N__42866\,
            I => \N__42859\
        );

    \I__8882\ : InMux
    port map (
            O => \N__42865\,
            I => \N__42856\
        );

    \I__8881\ : Odrv4
    port map (
            O => \N__42862\,
            I => n6
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__42859\,
            I => n6
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__42856\,
            I => n6
        );

    \I__8878\ : CascadeMux
    port map (
            O => \N__42849\,
            I => \N__42843\
        );

    \I__8877\ : CascadeMux
    port map (
            O => \N__42848\,
            I => \N__42840\
        );

    \I__8876\ : InMux
    port map (
            O => \N__42847\,
            I => \N__42837\
        );

    \I__8875\ : InMux
    port map (
            O => \N__42846\,
            I => \N__42834\
        );

    \I__8874\ : InMux
    port map (
            O => \N__42843\,
            I => \N__42829\
        );

    \I__8873\ : InMux
    port map (
            O => \N__42840\,
            I => \N__42829\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__42837\,
            I => n13641
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__42834\,
            I => n13641
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__42829\,
            I => n13641
        );

    \I__8869\ : CascadeMux
    port map (
            O => \N__42822\,
            I => \n13648_cascade_\
        );

    \I__8868\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42816\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__42816\,
            I => \N__42810\
        );

    \I__8866\ : CascadeMux
    port map (
            O => \N__42815\,
            I => \N__42807\
        );

    \I__8865\ : CascadeMux
    port map (
            O => \N__42814\,
            I => \N__42804\
        );

    \I__8864\ : InMux
    port map (
            O => \N__42813\,
            I => \N__42801\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__42810\,
            I => \N__42798\
        );

    \I__8862\ : InMux
    port map (
            O => \N__42807\,
            I => \N__42793\
        );

    \I__8861\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42793\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__42801\,
            I => encoder0_position_27
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__42798\,
            I => encoder0_position_27
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__42793\,
            I => encoder0_position_27
        );

    \I__8857\ : CascadeMux
    port map (
            O => \N__42786\,
            I => \N__42783\
        );

    \I__8856\ : InMux
    port map (
            O => \N__42783\,
            I => \N__42779\
        );

    \I__8855\ : InMux
    port map (
            O => \N__42782\,
            I => \N__42775\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__42779\,
            I => \N__42772\
        );

    \I__8853\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42769\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__42775\,
            I => n832
        );

    \I__8851\ : Odrv4
    port map (
            O => \N__42772\,
            I => n832
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__42769\,
            I => n832
        );

    \I__8849\ : InMux
    port map (
            O => \N__42762\,
            I => \N__42759\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__42759\,
            I => \N__42756\
        );

    \I__8847\ : Odrv4
    port map (
            O => \N__42756\,
            I => n999
        );

    \I__8846\ : CascadeMux
    port map (
            O => \N__42753\,
            I => \N__42749\
        );

    \I__8845\ : CascadeMux
    port map (
            O => \N__42752\,
            I => \N__42746\
        );

    \I__8844\ : InMux
    port map (
            O => \N__42749\,
            I => \N__42742\
        );

    \I__8843\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42739\
        );

    \I__8842\ : InMux
    port map (
            O => \N__42745\,
            I => \N__42736\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__42742\,
            I => n932
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__42739\,
            I => n932
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__42736\,
            I => n932
        );

    \I__8838\ : CascadeMux
    port map (
            O => \N__42729\,
            I => \N__42725\
        );

    \I__8837\ : InMux
    port map (
            O => \N__42728\,
            I => \N__42721\
        );

    \I__8836\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42718\
        );

    \I__8835\ : CascadeMux
    port map (
            O => \N__42724\,
            I => \N__42715\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__42721\,
            I => \N__42710\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__42718\,
            I => \N__42710\
        );

    \I__8832\ : InMux
    port map (
            O => \N__42715\,
            I => \N__42706\
        );

    \I__8831\ : Span4Mux_h
    port map (
            O => \N__42710\,
            I => \N__42703\
        );

    \I__8830\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42700\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__42706\,
            I => encoder0_position_26
        );

    \I__8828\ : Odrv4
    port map (
            O => \N__42703\,
            I => encoder0_position_26
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__42700\,
            I => encoder0_position_26
        );

    \I__8826\ : InMux
    port map (
            O => \N__42693\,
            I => \N__42690\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__42690\,
            I => n13650
        );

    \I__8824\ : CascadeMux
    port map (
            O => \N__42687\,
            I => \N__42684\
        );

    \I__8823\ : InMux
    port map (
            O => \N__42684\,
            I => \N__42679\
        );

    \I__8822\ : CascadeMux
    port map (
            O => \N__42683\,
            I => \N__42676\
        );

    \I__8821\ : InMux
    port map (
            O => \N__42682\,
            I => \N__42673\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__42679\,
            I => \N__42670\
        );

    \I__8819\ : InMux
    port map (
            O => \N__42676\,
            I => \N__42667\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__42673\,
            I => n833
        );

    \I__8817\ : Odrv4
    port map (
            O => \N__42670\,
            I => n833
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__42667\,
            I => n833
        );

    \I__8815\ : InMux
    port map (
            O => \N__42660\,
            I => \N__42657\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__42657\,
            I => \N__42654\
        );

    \I__8813\ : Span4Mux_h
    port map (
            O => \N__42654\,
            I => \N__42651\
        );

    \I__8812\ : Span4Mux_h
    port map (
            O => \N__42651\,
            I => \N__42648\
        );

    \I__8811\ : Odrv4
    port map (
            O => \N__42648\,
            I => encoder0_position_scaled_3
        );

    \I__8810\ : CascadeMux
    port map (
            O => \N__42645\,
            I => \N__42642\
        );

    \I__8809\ : InMux
    port map (
            O => \N__42642\,
            I => \N__42638\
        );

    \I__8808\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42635\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__42638\,
            I => n293
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__42635\,
            I => n293
        );

    \I__8805\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42627\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__42627\,
            I => n2542
        );

    \I__8803\ : InMux
    port map (
            O => \N__42624\,
            I => \bfn_12_25_0_\
        );

    \I__8802\ : CascadeMux
    port map (
            O => \N__42621\,
            I => \N__42618\
        );

    \I__8801\ : InMux
    port map (
            O => \N__42618\,
            I => \N__42615\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__42615\,
            I => \N__42612\
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__42612\,
            I => n292
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__42609\,
            I => \N__42606\
        );

    \I__8797\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42603\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__42603\,
            I => n2541
        );

    \I__8795\ : InMux
    port map (
            O => \N__42600\,
            I => n12482
        );

    \I__8794\ : CascadeMux
    port map (
            O => \N__42597\,
            I => \N__42594\
        );

    \I__8793\ : InMux
    port map (
            O => \N__42594\,
            I => \N__42591\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__42591\,
            I => n174
        );

    \I__8791\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42585\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__42585\,
            I => n2540
        );

    \I__8789\ : InMux
    port map (
            O => \N__42582\,
            I => n12483
        );

    \I__8788\ : InMux
    port map (
            O => \N__42579\,
            I => n12499
        );

    \I__8787\ : CascadeMux
    port map (
            O => \N__42576\,
            I => \N__42573\
        );

    \I__8786\ : InMux
    port map (
            O => \N__42573\,
            I => \N__42570\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__42570\,
            I => n1001
        );

    \I__8784\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42563\
        );

    \I__8783\ : InMux
    port map (
            O => \N__42566\,
            I => \N__42560\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__42563\,
            I => n927
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__42560\,
            I => n927
        );

    \I__8780\ : CascadeMux
    port map (
            O => \N__42555\,
            I => \n14466_cascade_\
        );

    \I__8779\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42549\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__42549\,
            I => n11940
        );

    \I__8777\ : CascadeMux
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__8776\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42540\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__42540\,
            I => \N__42535\
        );

    \I__8774\ : InMux
    port map (
            O => \N__42539\,
            I => \N__42530\
        );

    \I__8773\ : InMux
    port map (
            O => \N__42538\,
            I => \N__42530\
        );

    \I__8772\ : Odrv4
    port map (
            O => \N__42535\,
            I => n930
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__42530\,
            I => n930
        );

    \I__8770\ : CascadeMux
    port map (
            O => \N__42525\,
            I => \n960_cascade_\
        );

    \I__8769\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42519\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__42519\,
            I => n997
        );

    \I__8767\ : CascadeMux
    port map (
            O => \N__42516\,
            I => \N__42512\
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__42515\,
            I => \N__42508\
        );

    \I__8765\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42505\
        );

    \I__8764\ : InMux
    port map (
            O => \N__42511\,
            I => \N__42500\
        );

    \I__8763\ : InMux
    port map (
            O => \N__42508\,
            I => \N__42500\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__42505\,
            I => n929
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__42500\,
            I => n929
        );

    \I__8760\ : CascadeMux
    port map (
            O => \N__42495\,
            I => \N__42492\
        );

    \I__8759\ : InMux
    port map (
            O => \N__42492\,
            I => \N__42489\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__42489\,
            I => n996
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__42486\,
            I => \n1028_cascade_\
        );

    \I__8756\ : InMux
    port map (
            O => \N__42483\,
            I => \N__42480\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__42480\,
            I => n998
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__42477\,
            I => \N__42474\
        );

    \I__8753\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42470\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__42473\,
            I => \N__42467\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__42470\,
            I => \N__42464\
        );

    \I__8750\ : InMux
    port map (
            O => \N__42467\,
            I => \N__42461\
        );

    \I__8749\ : Odrv4
    port map (
            O => \N__42464\,
            I => n931
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__42461\,
            I => n931
        );

    \I__8747\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42453\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__42453\,
            I => \N__42450\
        );

    \I__8745\ : Span4Mux_h
    port map (
            O => \N__42450\,
            I => \N__42447\
        );

    \I__8744\ : Odrv4
    port map (
            O => \N__42447\,
            I => encoder0_position_scaled_8
        );

    \I__8743\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42438\
        );

    \I__8742\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42438\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__42438\,
            I => \N__42434\
        );

    \I__8740\ : InMux
    port map (
            O => \N__42437\,
            I => \N__42431\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__42434\,
            I => \N__42428\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__42431\,
            I => encoder0_position_15
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__42428\,
            I => encoder0_position_15
        );

    \I__8736\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__42420\,
            I => \N__42416\
        );

    \I__8734\ : InMux
    port map (
            O => \N__42419\,
            I => \N__42413\
        );

    \I__8733\ : Span4Mux_h
    port map (
            O => \N__42416\,
            I => \N__42410\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__42413\,
            I => \N__42407\
        );

    \I__8731\ : Sp12to4
    port map (
            O => \N__42410\,
            I => \N__42403\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__42407\,
            I => \N__42400\
        );

    \I__8729\ : InMux
    port map (
            O => \N__42406\,
            I => \N__42397\
        );

    \I__8728\ : Odrv12
    port map (
            O => \N__42403\,
            I => n304
        );

    \I__8727\ : Odrv4
    port map (
            O => \N__42400\,
            I => n304
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__42397\,
            I => n304
        );

    \I__8725\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42387\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__42387\,
            I => \N__42384\
        );

    \I__8723\ : Span12Mux_h
    port map (
            O => \N__42384\,
            I => \N__42381\
        );

    \I__8722\ : Odrv12
    port map (
            O => \N__42381\,
            I => n15
        );

    \I__8721\ : InMux
    port map (
            O => \N__42378\,
            I => \N__42375\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__42375\,
            I => \N__42370\
        );

    \I__8719\ : InMux
    port map (
            O => \N__42374\,
            I => \N__42367\
        );

    \I__8718\ : InMux
    port map (
            O => \N__42373\,
            I => \N__42364\
        );

    \I__8717\ : Span4Mux_h
    port map (
            O => \N__42370\,
            I => \N__42361\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__42367\,
            I => \N__42358\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__42364\,
            I => encoder0_position_18
        );

    \I__8714\ : Odrv4
    port map (
            O => \N__42361\,
            I => encoder0_position_18
        );

    \I__8713\ : Odrv4
    port map (
            O => \N__42358\,
            I => encoder0_position_18
        );

    \I__8712\ : InMux
    port map (
            O => \N__42351\,
            I => \bfn_12_22_0_\
        );

    \I__8711\ : InMux
    port map (
            O => \N__42348\,
            I => n12493
        );

    \I__8710\ : InMux
    port map (
            O => \N__42345\,
            I => n12494
        );

    \I__8709\ : InMux
    port map (
            O => \N__42342\,
            I => n12495
        );

    \I__8708\ : InMux
    port map (
            O => \N__42339\,
            I => n12496
        );

    \I__8707\ : InMux
    port map (
            O => \N__42336\,
            I => n12497
        );

    \I__8706\ : InMux
    port map (
            O => \N__42333\,
            I => n12498
        );

    \I__8705\ : InMux
    port map (
            O => \N__42330\,
            I => \N__42327\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__42327\,
            I => \N__42323\
        );

    \I__8703\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42320\
        );

    \I__8702\ : Span4Mux_h
    port map (
            O => \N__42323\,
            I => \N__42317\
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__42320\,
            I => \N__42311\
        );

    \I__8700\ : Span4Mux_v
    port map (
            O => \N__42317\,
            I => \N__42311\
        );

    \I__8699\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42308\
        );

    \I__8698\ : Odrv4
    port map (
            O => \N__42311\,
            I => n2
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__42308\,
            I => n2
        );

    \I__8696\ : InMux
    port map (
            O => \N__42303\,
            I => \N__42300\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__42300\,
            I => \N__42297\
        );

    \I__8694\ : Span4Mux_h
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__8693\ : Odrv4
    port map (
            O => \N__42294\,
            I => n16
        );

    \I__8692\ : InMux
    port map (
            O => \N__42291\,
            I => \N__42284\
        );

    \I__8691\ : InMux
    port map (
            O => \N__42290\,
            I => \N__42284\
        );

    \I__8690\ : CascadeMux
    port map (
            O => \N__42289\,
            I => \N__42281\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__42284\,
            I => \N__42278\
        );

    \I__8688\ : InMux
    port map (
            O => \N__42281\,
            I => \N__42275\
        );

    \I__8687\ : Span4Mux_h
    port map (
            O => \N__42278\,
            I => \N__42272\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__42275\,
            I => encoder0_position_17
        );

    \I__8685\ : Odrv4
    port map (
            O => \N__42272\,
            I => encoder0_position_17
        );

    \I__8684\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42264\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__42264\,
            I => \N__42261\
        );

    \I__8682\ : Span4Mux_h
    port map (
            O => \N__42261\,
            I => \N__42258\
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__42258\,
            I => n30
        );

    \I__8680\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42252\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__42252\,
            I => \N__42247\
        );

    \I__8678\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42244\
        );

    \I__8677\ : CascadeMux
    port map (
            O => \N__42250\,
            I => \N__42241\
        );

    \I__8676\ : Span4Mux_v
    port map (
            O => \N__42247\,
            I => \N__42236\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__42244\,
            I => \N__42236\
        );

    \I__8674\ : InMux
    port map (
            O => \N__42241\,
            I => \N__42233\
        );

    \I__8673\ : Span4Mux_h
    port map (
            O => \N__42236\,
            I => \N__42230\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__42233\,
            I => encoder0_position_3
        );

    \I__8671\ : Odrv4
    port map (
            O => \N__42230\,
            I => encoder0_position_3
        );

    \I__8670\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42221\
        );

    \I__8669\ : InMux
    port map (
            O => \N__42224\,
            I => \N__42217\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__42221\,
            I => \N__42214\
        );

    \I__8667\ : InMux
    port map (
            O => \N__42220\,
            I => \N__42211\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__42217\,
            I => \N__42204\
        );

    \I__8665\ : Span4Mux_h
    port map (
            O => \N__42214\,
            I => \N__42204\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__42211\,
            I => \N__42204\
        );

    \I__8663\ : Span4Mux_h
    port map (
            O => \N__42204\,
            I => \N__42201\
        );

    \I__8662\ : Sp12to4
    port map (
            O => \N__42201\,
            I => \N__42198\
        );

    \I__8661\ : Span12Mux_v
    port map (
            O => \N__42198\,
            I => \N__42195\
        );

    \I__8660\ : Odrv12
    port map (
            O => \N__42195\,
            I => n316
        );

    \I__8659\ : CascadeMux
    port map (
            O => \N__42192\,
            I => \N__42168\
        );

    \I__8658\ : CascadeMux
    port map (
            O => \N__42191\,
            I => \N__42165\
        );

    \I__8657\ : CascadeMux
    port map (
            O => \N__42190\,
            I => \N__42162\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__42189\,
            I => \N__42159\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__42188\,
            I => \N__42156\
        );

    \I__8654\ : CascadeMux
    port map (
            O => \N__42187\,
            I => \N__42153\
        );

    \I__8653\ : CascadeMux
    port map (
            O => \N__42186\,
            I => \N__42150\
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__42185\,
            I => \N__42147\
        );

    \I__8651\ : CascadeMux
    port map (
            O => \N__42184\,
            I => \N__42144\
        );

    \I__8650\ : CascadeMux
    port map (
            O => \N__42183\,
            I => \N__42141\
        );

    \I__8649\ : CascadeMux
    port map (
            O => \N__42182\,
            I => \N__42138\
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__42181\,
            I => \N__42135\
        );

    \I__8647\ : CascadeMux
    port map (
            O => \N__42180\,
            I => \N__42132\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__42179\,
            I => \N__42129\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__42178\,
            I => \N__42125\
        );

    \I__8644\ : CascadeMux
    port map (
            O => \N__42177\,
            I => \N__42122\
        );

    \I__8643\ : CascadeMux
    port map (
            O => \N__42176\,
            I => \N__42119\
        );

    \I__8642\ : CascadeMux
    port map (
            O => \N__42175\,
            I => \N__42116\
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__42174\,
            I => \N__42112\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__42173\,
            I => \N__42109\
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__42172\,
            I => \N__42106\
        );

    \I__8638\ : CascadeMux
    port map (
            O => \N__42171\,
            I => \N__42103\
        );

    \I__8637\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42093\
        );

    \I__8636\ : InMux
    port map (
            O => \N__42165\,
            I => \N__42093\
        );

    \I__8635\ : InMux
    port map (
            O => \N__42162\,
            I => \N__42093\
        );

    \I__8634\ : InMux
    port map (
            O => \N__42159\,
            I => \N__42093\
        );

    \I__8633\ : InMux
    port map (
            O => \N__42156\,
            I => \N__42084\
        );

    \I__8632\ : InMux
    port map (
            O => \N__42153\,
            I => \N__42084\
        );

    \I__8631\ : InMux
    port map (
            O => \N__42150\,
            I => \N__42084\
        );

    \I__8630\ : InMux
    port map (
            O => \N__42147\,
            I => \N__42084\
        );

    \I__8629\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42075\
        );

    \I__8628\ : InMux
    port map (
            O => \N__42141\,
            I => \N__42075\
        );

    \I__8627\ : InMux
    port map (
            O => \N__42138\,
            I => \N__42075\
        );

    \I__8626\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42075\
        );

    \I__8625\ : InMux
    port map (
            O => \N__42132\,
            I => \N__42066\
        );

    \I__8624\ : InMux
    port map (
            O => \N__42129\,
            I => \N__42066\
        );

    \I__8623\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42066\
        );

    \I__8622\ : InMux
    port map (
            O => \N__42125\,
            I => \N__42066\
        );

    \I__8621\ : InMux
    port map (
            O => \N__42122\,
            I => \N__42057\
        );

    \I__8620\ : InMux
    port map (
            O => \N__42119\,
            I => \N__42057\
        );

    \I__8619\ : InMux
    port map (
            O => \N__42116\,
            I => \N__42057\
        );

    \I__8618\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42057\
        );

    \I__8617\ : InMux
    port map (
            O => \N__42112\,
            I => \N__42048\
        );

    \I__8616\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42048\
        );

    \I__8615\ : InMux
    port map (
            O => \N__42106\,
            I => \N__42048\
        );

    \I__8614\ : InMux
    port map (
            O => \N__42103\,
            I => \N__42048\
        );

    \I__8613\ : CascadeMux
    port map (
            O => \N__42102\,
            I => \N__42045\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__42093\,
            I => \N__42040\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__42084\,
            I => \N__42040\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__42075\,
            I => \N__42033\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__42066\,
            I => \N__42033\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__42057\,
            I => \N__42033\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__42048\,
            I => \N__42030\
        );

    \I__8606\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42027\
        );

    \I__8605\ : Span4Mux_v
    port map (
            O => \N__42040\,
            I => \N__42022\
        );

    \I__8604\ : Span4Mux_v
    port map (
            O => \N__42033\,
            I => \N__42022\
        );

    \I__8603\ : Span4Mux_h
    port map (
            O => \N__42030\,
            I => \N__42017\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__42027\,
            I => \N__42017\
        );

    \I__8601\ : Span4Mux_h
    port map (
            O => \N__42022\,
            I => \N__42012\
        );

    \I__8600\ : Span4Mux_v
    port map (
            O => \N__42017\,
            I => \N__42012\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__42012\,
            I => n2_adj_623
        );

    \I__8598\ : InMux
    port map (
            O => \N__42009\,
            I => \N__42006\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__42006\,
            I => \N__42003\
        );

    \I__8596\ : Span4Mux_v
    port map (
            O => \N__42003\,
            I => \N__42000\
        );

    \I__8595\ : Span4Mux_h
    port map (
            O => \N__42000\,
            I => \N__41997\
        );

    \I__8594\ : Odrv4
    port map (
            O => \N__41997\,
            I => encoder0_position_scaled_7
        );

    \I__8593\ : InMux
    port map (
            O => \N__41994\,
            I => \N__41989\
        );

    \I__8592\ : InMux
    port map (
            O => \N__41993\,
            I => \N__41986\
        );

    \I__8591\ : CascadeMux
    port map (
            O => \N__41992\,
            I => \N__41983\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__41989\,
            I => \N__41980\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__41986\,
            I => \N__41977\
        );

    \I__8588\ : InMux
    port map (
            O => \N__41983\,
            I => \N__41974\
        );

    \I__8587\ : Span4Mux_h
    port map (
            O => \N__41980\,
            I => \N__41971\
        );

    \I__8586\ : Span4Mux_h
    port map (
            O => \N__41977\,
            I => \N__41968\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__41974\,
            I => encoder0_position_23
        );

    \I__8584\ : Odrv4
    port map (
            O => \N__41971\,
            I => encoder0_position_23
        );

    \I__8583\ : Odrv4
    port map (
            O => \N__41968\,
            I => encoder0_position_23
        );

    \I__8582\ : CascadeMux
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__8581\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__41955\,
            I => \N__41952\
        );

    \I__8579\ : Span4Mux_v
    port map (
            O => \N__41952\,
            I => \N__41949\
        );

    \I__8578\ : Odrv4
    port map (
            O => \N__41949\,
            I => n10_adj_631
        );

    \I__8577\ : CascadeMux
    port map (
            O => \N__41946\,
            I => \N__41943\
        );

    \I__8576\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__8574\ : Span4Mux_v
    port map (
            O => \N__41937\,
            I => \N__41934\
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__41934\,
            I => n18_adj_639
        );

    \I__8572\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41928\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41925\
        );

    \I__8570\ : Span4Mux_v
    port map (
            O => \N__41925\,
            I => \N__41922\
        );

    \I__8569\ : Odrv4
    port map (
            O => \N__41922\,
            I => n17
        );

    \I__8568\ : CascadeMux
    port map (
            O => \N__41919\,
            I => \N__41915\
        );

    \I__8567\ : InMux
    port map (
            O => \N__41918\,
            I => \N__41912\
        );

    \I__8566\ : InMux
    port map (
            O => \N__41915\,
            I => \N__41909\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__41912\,
            I => \N__41905\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__41909\,
            I => \N__41902\
        );

    \I__8563\ : InMux
    port map (
            O => \N__41908\,
            I => \N__41899\
        );

    \I__8562\ : Span4Mux_h
    port map (
            O => \N__41905\,
            I => \N__41896\
        );

    \I__8561\ : Span4Mux_v
    port map (
            O => \N__41902\,
            I => \N__41893\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__41899\,
            I => encoder0_position_16
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__41896\,
            I => encoder0_position_16
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__41893\,
            I => encoder0_position_16
        );

    \I__8557\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41883\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41880\
        );

    \I__8555\ : Span4Mux_h
    port map (
            O => \N__41880\,
            I => \N__41877\
        );

    \I__8554\ : Odrv4
    port map (
            O => \N__41877\,
            I => n18
        );

    \I__8553\ : InMux
    port map (
            O => \N__41874\,
            I => \bfn_12_19_0_\
        );

    \I__8552\ : CascadeMux
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__8551\ : InMux
    port map (
            O => \N__41868\,
            I => \N__41865\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__41865\,
            I => \N__41862\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__41862\,
            I => n1885
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__41859\,
            I => \n1722_cascade_\
        );

    \I__8547\ : InMux
    port map (
            O => \N__41856\,
            I => \N__41851\
        );

    \I__8546\ : InMux
    port map (
            O => \N__41855\,
            I => \N__41848\
        );

    \I__8545\ : InMux
    port map (
            O => \N__41854\,
            I => \N__41845\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__41851\,
            I => n1821
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__41848\,
            I => n1821
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__41845\,
            I => n1821
        );

    \I__8541\ : CascadeMux
    port map (
            O => \N__41838\,
            I => \N__41835\
        );

    \I__8540\ : InMux
    port map (
            O => \N__41835\,
            I => \N__41831\
        );

    \I__8539\ : CascadeMux
    port map (
            O => \N__41834\,
            I => \N__41828\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__41831\,
            I => \N__41824\
        );

    \I__8537\ : InMux
    port map (
            O => \N__41828\,
            I => \N__41821\
        );

    \I__8536\ : InMux
    port map (
            O => \N__41827\,
            I => \N__41818\
        );

    \I__8535\ : Span4Mux_h
    port map (
            O => \N__41824\,
            I => \N__41815\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__41821\,
            I => \N__41810\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__41818\,
            I => \N__41810\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__41815\,
            I => n1827
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__41810\,
            I => n1827
        );

    \I__8530\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41800\
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__41804\,
            I => \N__41797\
        );

    \I__8528\ : CascadeMux
    port map (
            O => \N__41803\,
            I => \N__41793\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__41800\,
            I => \N__41786\
        );

    \I__8526\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41780\
        );

    \I__8525\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41780\
        );

    \I__8524\ : InMux
    port map (
            O => \N__41793\,
            I => \N__41777\
        );

    \I__8523\ : CascadeMux
    port map (
            O => \N__41792\,
            I => \N__41774\
        );

    \I__8522\ : CascadeMux
    port map (
            O => \N__41791\,
            I => \N__41771\
        );

    \I__8521\ : CascadeMux
    port map (
            O => \N__41790\,
            I => \N__41764\
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__41789\,
            I => \N__41761\
        );

    \I__8519\ : Span12Mux_s10_h
    port map (
            O => \N__41786\,
            I => \N__41755\
        );

    \I__8518\ : InMux
    port map (
            O => \N__41785\,
            I => \N__41752\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__41780\,
            I => \N__41747\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__41777\,
            I => \N__41747\
        );

    \I__8515\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41738\
        );

    \I__8514\ : InMux
    port map (
            O => \N__41771\,
            I => \N__41738\
        );

    \I__8513\ : InMux
    port map (
            O => \N__41770\,
            I => \N__41738\
        );

    \I__8512\ : InMux
    port map (
            O => \N__41769\,
            I => \N__41738\
        );

    \I__8511\ : InMux
    port map (
            O => \N__41768\,
            I => \N__41727\
        );

    \I__8510\ : InMux
    port map (
            O => \N__41767\,
            I => \N__41727\
        );

    \I__8509\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41727\
        );

    \I__8508\ : InMux
    port map (
            O => \N__41761\,
            I => \N__41727\
        );

    \I__8507\ : InMux
    port map (
            O => \N__41760\,
            I => \N__41727\
        );

    \I__8506\ : InMux
    port map (
            O => \N__41759\,
            I => \N__41722\
        );

    \I__8505\ : InMux
    port map (
            O => \N__41758\,
            I => \N__41722\
        );

    \I__8504\ : Odrv12
    port map (
            O => \N__41755\,
            I => n1752
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__41752\,
            I => n1752
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__41747\,
            I => n1752
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__41738\,
            I => n1752
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__41727\,
            I => n1752
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__41722\,
            I => n1752
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__41709\,
            I => \N__41706\
        );

    \I__8497\ : InMux
    port map (
            O => \N__41706\,
            I => \N__41703\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__41703\,
            I => \N__41700\
        );

    \I__8495\ : Span4Mux_h
    port map (
            O => \N__41700\,
            I => \N__41697\
        );

    \I__8494\ : Odrv4
    port map (
            O => \N__41697\,
            I => n16_adj_637
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__41694\,
            I => \N__41690\
        );

    \I__8492\ : CascadeMux
    port map (
            O => \N__41693\,
            I => \N__41687\
        );

    \I__8491\ : InMux
    port map (
            O => \N__41690\,
            I => \N__41684\
        );

    \I__8490\ : InMux
    port map (
            O => \N__41687\,
            I => \N__41681\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__41684\,
            I => n1826
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__41681\,
            I => n1826
        );

    \I__8487\ : InMux
    port map (
            O => \N__41676\,
            I => \N__41673\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__41673\,
            I => \N__41670\
        );

    \I__8485\ : Span4Mux_h
    port map (
            O => \N__41670\,
            I => \N__41667\
        );

    \I__8484\ : Odrv4
    port map (
            O => \N__41667\,
            I => n1893
        );

    \I__8483\ : InMux
    port map (
            O => \N__41664\,
            I => \bfn_12_18_0_\
        );

    \I__8482\ : CascadeMux
    port map (
            O => \N__41661\,
            I => \N__41657\
        );

    \I__8481\ : InMux
    port map (
            O => \N__41660\,
            I => \N__41653\
        );

    \I__8480\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41650\
        );

    \I__8479\ : InMux
    port map (
            O => \N__41656\,
            I => \N__41647\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__41653\,
            I => n1825
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__41650\,
            I => n1825
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__41647\,
            I => n1825
        );

    \I__8475\ : InMux
    port map (
            O => \N__41640\,
            I => \N__41637\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__41637\,
            I => \N__41634\
        );

    \I__8473\ : Odrv4
    port map (
            O => \N__41634\,
            I => n1892
        );

    \I__8472\ : InMux
    port map (
            O => \N__41631\,
            I => n12600
        );

    \I__8471\ : CascadeMux
    port map (
            O => \N__41628\,
            I => \N__41623\
        );

    \I__8470\ : CascadeMux
    port map (
            O => \N__41627\,
            I => \N__41620\
        );

    \I__8469\ : InMux
    port map (
            O => \N__41626\,
            I => \N__41617\
        );

    \I__8468\ : InMux
    port map (
            O => \N__41623\,
            I => \N__41614\
        );

    \I__8467\ : InMux
    port map (
            O => \N__41620\,
            I => \N__41611\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__41617\,
            I => n1824
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__41614\,
            I => n1824
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__41611\,
            I => n1824
        );

    \I__8463\ : InMux
    port map (
            O => \N__41604\,
            I => \N__41601\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__41601\,
            I => \N__41598\
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__41598\,
            I => n1891
        );

    \I__8460\ : InMux
    port map (
            O => \N__41595\,
            I => n12601
        );

    \I__8459\ : CascadeMux
    port map (
            O => \N__41592\,
            I => \N__41588\
        );

    \I__8458\ : InMux
    port map (
            O => \N__41591\,
            I => \N__41584\
        );

    \I__8457\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41581\
        );

    \I__8456\ : InMux
    port map (
            O => \N__41587\,
            I => \N__41578\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__41584\,
            I => n1823
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__41581\,
            I => n1823
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__41578\,
            I => n1823
        );

    \I__8452\ : CascadeMux
    port map (
            O => \N__41571\,
            I => \N__41568\
        );

    \I__8451\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41565\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__41565\,
            I => \N__41562\
        );

    \I__8449\ : Span4Mux_h
    port map (
            O => \N__41562\,
            I => \N__41559\
        );

    \I__8448\ : Odrv4
    port map (
            O => \N__41559\,
            I => n1890
        );

    \I__8447\ : InMux
    port map (
            O => \N__41556\,
            I => n12602
        );

    \I__8446\ : InMux
    port map (
            O => \N__41553\,
            I => \N__41549\
        );

    \I__8445\ : CascadeMux
    port map (
            O => \N__41552\,
            I => \N__41546\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__41549\,
            I => \N__41543\
        );

    \I__8443\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41540\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__41543\,
            I => \N__41536\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__41540\,
            I => \N__41533\
        );

    \I__8440\ : InMux
    port map (
            O => \N__41539\,
            I => \N__41530\
        );

    \I__8439\ : Odrv4
    port map (
            O => \N__41536\,
            I => n1822
        );

    \I__8438\ : Odrv4
    port map (
            O => \N__41533\,
            I => n1822
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__41530\,
            I => n1822
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__41523\,
            I => \N__41520\
        );

    \I__8435\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41517\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__41517\,
            I => \N__41514\
        );

    \I__8433\ : Odrv12
    port map (
            O => \N__41514\,
            I => n1889
        );

    \I__8432\ : InMux
    port map (
            O => \N__41511\,
            I => n12603
        );

    \I__8431\ : InMux
    port map (
            O => \N__41508\,
            I => \N__41505\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__41505\,
            I => n1888
        );

    \I__8429\ : InMux
    port map (
            O => \N__41502\,
            I => n12604
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__41499\,
            I => \N__41496\
        );

    \I__8427\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41492\
        );

    \I__8426\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41489\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__41492\,
            I => \N__41486\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__41489\,
            I => n1820
        );

    \I__8423\ : Odrv4
    port map (
            O => \N__41486\,
            I => n1820
        );

    \I__8422\ : InMux
    port map (
            O => \N__41481\,
            I => \N__41478\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__41478\,
            I => n1887
        );

    \I__8420\ : InMux
    port map (
            O => \N__41475\,
            I => n12605
        );

    \I__8419\ : CascadeMux
    port map (
            O => \N__41472\,
            I => \N__41468\
        );

    \I__8418\ : InMux
    port map (
            O => \N__41471\,
            I => \N__41465\
        );

    \I__8417\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41462\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__41465\,
            I => n1819
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__41462\,
            I => n1819
        );

    \I__8414\ : InMux
    port map (
            O => \N__41457\,
            I => \N__41454\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__41454\,
            I => n1886
        );

    \I__8412\ : InMux
    port map (
            O => \N__41451\,
            I => n12606
        );

    \I__8411\ : InMux
    port map (
            O => \N__41448\,
            I => \N__41445\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__41445\,
            I => \N__41442\
        );

    \I__8409\ : Odrv4
    port map (
            O => \N__41442\,
            I => n1901
        );

    \I__8408\ : InMux
    port map (
            O => \N__41439\,
            I => \bfn_12_17_0_\
        );

    \I__8407\ : CascadeMux
    port map (
            O => \N__41436\,
            I => \N__41433\
        );

    \I__8406\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41428\
        );

    \I__8405\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41425\
        );

    \I__8404\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41422\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__41428\,
            I => \N__41419\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__41425\,
            I => n1833
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__41422\,
            I => n1833
        );

    \I__8400\ : Odrv4
    port map (
            O => \N__41419\,
            I => n1833
        );

    \I__8399\ : InMux
    port map (
            O => \N__41412\,
            I => \N__41409\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__41409\,
            I => \N__41406\
        );

    \I__8397\ : Span4Mux_v
    port map (
            O => \N__41406\,
            I => \N__41403\
        );

    \I__8396\ : Odrv4
    port map (
            O => \N__41403\,
            I => n1900
        );

    \I__8395\ : InMux
    port map (
            O => \N__41400\,
            I => n12592
        );

    \I__8394\ : CascadeMux
    port map (
            O => \N__41397\,
            I => \N__41393\
        );

    \I__8393\ : CascadeMux
    port map (
            O => \N__41396\,
            I => \N__41390\
        );

    \I__8392\ : InMux
    port map (
            O => \N__41393\,
            I => \N__41387\
        );

    \I__8391\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41384\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__41387\,
            I => \N__41381\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__41384\,
            I => n1832
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__41381\,
            I => n1832
        );

    \I__8387\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41373\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__41373\,
            I => \N__41370\
        );

    \I__8385\ : Odrv4
    port map (
            O => \N__41370\,
            I => n1899
        );

    \I__8384\ : InMux
    port map (
            O => \N__41367\,
            I => n12593
        );

    \I__8383\ : CascadeMux
    port map (
            O => \N__41364\,
            I => \N__41360\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__41363\,
            I => \N__41357\
        );

    \I__8381\ : InMux
    port map (
            O => \N__41360\,
            I => \N__41354\
        );

    \I__8380\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41350\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__41354\,
            I => \N__41347\
        );

    \I__8378\ : InMux
    port map (
            O => \N__41353\,
            I => \N__41344\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__41350\,
            I => n1831
        );

    \I__8376\ : Odrv4
    port map (
            O => \N__41347\,
            I => n1831
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__41344\,
            I => n1831
        );

    \I__8374\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41334\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__41334\,
            I => \N__41331\
        );

    \I__8372\ : Span4Mux_v
    port map (
            O => \N__41331\,
            I => \N__41328\
        );

    \I__8371\ : Odrv4
    port map (
            O => \N__41328\,
            I => n1898
        );

    \I__8370\ : InMux
    port map (
            O => \N__41325\,
            I => n12594
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__41322\,
            I => \N__41317\
        );

    \I__8368\ : InMux
    port map (
            O => \N__41321\,
            I => \N__41312\
        );

    \I__8367\ : InMux
    port map (
            O => \N__41320\,
            I => \N__41312\
        );

    \I__8366\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41309\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__41312\,
            I => \N__41304\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__41309\,
            I => \N__41304\
        );

    \I__8363\ : Odrv4
    port map (
            O => \N__41304\,
            I => n1830
        );

    \I__8362\ : InMux
    port map (
            O => \N__41301\,
            I => \N__41298\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__41298\,
            I => n1897
        );

    \I__8360\ : InMux
    port map (
            O => \N__41295\,
            I => n12595
        );

    \I__8359\ : CascadeMux
    port map (
            O => \N__41292\,
            I => \N__41287\
        );

    \I__8358\ : InMux
    port map (
            O => \N__41291\,
            I => \N__41282\
        );

    \I__8357\ : InMux
    port map (
            O => \N__41290\,
            I => \N__41282\
        );

    \I__8356\ : InMux
    port map (
            O => \N__41287\,
            I => \N__41279\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__41282\,
            I => n1829
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__41279\,
            I => n1829
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__41274\,
            I => \N__41271\
        );

    \I__8352\ : InMux
    port map (
            O => \N__41271\,
            I => \N__41268\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__41268\,
            I => n1896
        );

    \I__8350\ : InMux
    port map (
            O => \N__41265\,
            I => n12596
        );

    \I__8349\ : CascadeMux
    port map (
            O => \N__41262\,
            I => \N__41258\
        );

    \I__8348\ : InMux
    port map (
            O => \N__41261\,
            I => \N__41254\
        );

    \I__8347\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41251\
        );

    \I__8346\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41248\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__41254\,
            I => n1828
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__41251\,
            I => n1828
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__41248\,
            I => n1828
        );

    \I__8342\ : CascadeMux
    port map (
            O => \N__41241\,
            I => \N__41238\
        );

    \I__8341\ : InMux
    port map (
            O => \N__41238\,
            I => \N__41235\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__41235\,
            I => \N__41232\
        );

    \I__8339\ : Odrv4
    port map (
            O => \N__41232\,
            I => n1895
        );

    \I__8338\ : InMux
    port map (
            O => \N__41229\,
            I => n12597
        );

    \I__8337\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41223\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41220\
        );

    \I__8335\ : Odrv4
    port map (
            O => \N__41220\,
            I => n1894
        );

    \I__8334\ : InMux
    port map (
            O => \N__41217\,
            I => n12598
        );

    \I__8333\ : InMux
    port map (
            O => \N__41214\,
            I => \N__41211\
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__41211\,
            I => n6_adj_677
        );

    \I__8331\ : InMux
    port map (
            O => \N__41208\,
            I => n13106
        );

    \I__8330\ : CascadeMux
    port map (
            O => \N__41205\,
            I => \N__41201\
        );

    \I__8329\ : CascadeMux
    port map (
            O => \N__41204\,
            I => \N__41198\
        );

    \I__8328\ : InMux
    port map (
            O => \N__41201\,
            I => \N__41192\
        );

    \I__8327\ : InMux
    port map (
            O => \N__41198\,
            I => \N__41192\
        );

    \I__8326\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41189\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__41192\,
            I => blink_counter_21
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__41189\,
            I => blink_counter_21
        );

    \I__8323\ : InMux
    port map (
            O => \N__41184\,
            I => n13107
        );

    \I__8322\ : InMux
    port map (
            O => \N__41181\,
            I => \N__41174\
        );

    \I__8321\ : InMux
    port map (
            O => \N__41180\,
            I => \N__41174\
        );

    \I__8320\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41171\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__41174\,
            I => blink_counter_22
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__41171\,
            I => blink_counter_22
        );

    \I__8317\ : InMux
    port map (
            O => \N__41166\,
            I => n13108
        );

    \I__8316\ : InMux
    port map (
            O => \N__41163\,
            I => \N__41156\
        );

    \I__8315\ : InMux
    port map (
            O => \N__41162\,
            I => \N__41156\
        );

    \I__8314\ : InMux
    port map (
            O => \N__41161\,
            I => \N__41153\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__41156\,
            I => blink_counter_23
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__41153\,
            I => blink_counter_23
        );

    \I__8311\ : InMux
    port map (
            O => \N__41148\,
            I => n13109
        );

    \I__8310\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41138\
        );

    \I__8309\ : InMux
    port map (
            O => \N__41144\,
            I => \N__41138\
        );

    \I__8308\ : InMux
    port map (
            O => \N__41143\,
            I => \N__41135\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__41138\,
            I => blink_counter_24
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__41135\,
            I => blink_counter_24
        );

    \I__8305\ : InMux
    port map (
            O => \N__41130\,
            I => \bfn_11_32_0_\
        );

    \I__8304\ : InMux
    port map (
            O => \N__41127\,
            I => n13111
        );

    \I__8303\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41121\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__41121\,
            I => \N__41117\
        );

    \I__8301\ : InMux
    port map (
            O => \N__41120\,
            I => \N__41114\
        );

    \I__8300\ : Odrv4
    port map (
            O => \N__41117\,
            I => blink_counter_25
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__41114\,
            I => blink_counter_25
        );

    \I__8298\ : InMux
    port map (
            O => \N__41109\,
            I => \N__41106\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__41103\
        );

    \I__8296\ : Odrv4
    port map (
            O => \N__41103\,
            I => \pwm_setpoint_23_N_171_19\
        );

    \I__8295\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41097\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__41097\,
            I => \N__41094\
        );

    \I__8293\ : Odrv4
    port map (
            O => \N__41094\,
            I => n8_adj_588
        );

    \I__8292\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41088\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__41088\,
            I => \N__41085\
        );

    \I__8290\ : Odrv4
    port map (
            O => \N__41085\,
            I => n5_adj_585
        );

    \I__8289\ : InMux
    port map (
            O => \N__41082\,
            I => \N__41079\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__41079\,
            I => n14_adj_685
        );

    \I__8287\ : InMux
    port map (
            O => \N__41076\,
            I => n13098
        );

    \I__8286\ : InMux
    port map (
            O => \N__41073\,
            I => \N__41070\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__41070\,
            I => n13_adj_684
        );

    \I__8284\ : InMux
    port map (
            O => \N__41067\,
            I => n13099
        );

    \I__8283\ : InMux
    port map (
            O => \N__41064\,
            I => \N__41061\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__41061\,
            I => n12_adj_683
        );

    \I__8281\ : InMux
    port map (
            O => \N__41058\,
            I => n13100
        );

    \I__8280\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41052\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__41052\,
            I => n11_adj_682
        );

    \I__8278\ : InMux
    port map (
            O => \N__41049\,
            I => n13101
        );

    \I__8277\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41043\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__41043\,
            I => n10_adj_681
        );

    \I__8275\ : InMux
    port map (
            O => \N__41040\,
            I => \bfn_11_31_0_\
        );

    \I__8274\ : InMux
    port map (
            O => \N__41037\,
            I => \N__41034\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__41034\,
            I => n9_adj_680
        );

    \I__8272\ : InMux
    port map (
            O => \N__41031\,
            I => n13103
        );

    \I__8271\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__41025\,
            I => n8_adj_679
        );

    \I__8269\ : InMux
    port map (
            O => \N__41022\,
            I => n13104
        );

    \I__8268\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41016\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__41016\,
            I => n7_adj_678
        );

    \I__8266\ : InMux
    port map (
            O => \N__41013\,
            I => n13105
        );

    \I__8265\ : InMux
    port map (
            O => \N__41010\,
            I => \N__41007\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__41007\,
            I => n23_adj_694
        );

    \I__8263\ : InMux
    port map (
            O => \N__41004\,
            I => n13089
        );

    \I__8262\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40998\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__40998\,
            I => n22_adj_693
        );

    \I__8260\ : InMux
    port map (
            O => \N__40995\,
            I => n13090
        );

    \I__8259\ : InMux
    port map (
            O => \N__40992\,
            I => \N__40989\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__40989\,
            I => n21_adj_692
        );

    \I__8257\ : InMux
    port map (
            O => \N__40986\,
            I => n13091
        );

    \I__8256\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40980\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__40980\,
            I => n20_adj_691
        );

    \I__8254\ : InMux
    port map (
            O => \N__40977\,
            I => n13092
        );

    \I__8253\ : InMux
    port map (
            O => \N__40974\,
            I => \N__40971\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__40971\,
            I => n19_adj_690
        );

    \I__8251\ : InMux
    port map (
            O => \N__40968\,
            I => n13093
        );

    \I__8250\ : InMux
    port map (
            O => \N__40965\,
            I => \N__40962\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__40962\,
            I => n18_adj_689
        );

    \I__8248\ : InMux
    port map (
            O => \N__40959\,
            I => \bfn_11_30_0_\
        );

    \I__8247\ : InMux
    port map (
            O => \N__40956\,
            I => \N__40953\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__40953\,
            I => n17_adj_688
        );

    \I__8245\ : InMux
    port map (
            O => \N__40950\,
            I => n13095
        );

    \I__8244\ : InMux
    port map (
            O => \N__40947\,
            I => \N__40944\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__40944\,
            I => n16_adj_687
        );

    \I__8242\ : InMux
    port map (
            O => \N__40941\,
            I => n13096
        );

    \I__8241\ : InMux
    port map (
            O => \N__40938\,
            I => \N__40935\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__40935\,
            I => n15_adj_686
        );

    \I__8239\ : InMux
    port map (
            O => \N__40932\,
            I => n13097
        );

    \I__8238\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40926\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__40926\,
            I => n12_adj_661
        );

    \I__8236\ : InMux
    port map (
            O => \N__40923\,
            I => \N__40920\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__40920\,
            I => \N__40917\
        );

    \I__8234\ : Span4Mux_h
    port map (
            O => \N__40917\,
            I => \N__40914\
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__40914\,
            I => \pwm_setpoint_23_N_171_7\
        );

    \I__8232\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40906\
        );

    \I__8231\ : InMux
    port map (
            O => \N__40910\,
            I => \N__40901\
        );

    \I__8230\ : InMux
    port map (
            O => \N__40909\,
            I => \N__40901\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__40906\,
            I => pwm_setpoint_16
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__40901\,
            I => pwm_setpoint_16
        );

    \I__8227\ : InMux
    port map (
            O => \N__40896\,
            I => \N__40891\
        );

    \I__8226\ : InMux
    port map (
            O => \N__40895\,
            I => \N__40886\
        );

    \I__8225\ : InMux
    port map (
            O => \N__40894\,
            I => \N__40886\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__40891\,
            I => pwm_setpoint_7
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__40886\,
            I => pwm_setpoint_7
        );

    \I__8222\ : InMux
    port map (
            O => \N__40881\,
            I => \N__40878\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__40878\,
            I => n15119
        );

    \I__8220\ : InMux
    port map (
            O => \N__40875\,
            I => \N__40872\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__40872\,
            I => \N__40869\
        );

    \I__8218\ : Span4Mux_h
    port map (
            O => \N__40869\,
            I => \N__40866\
        );

    \I__8217\ : Span4Mux_v
    port map (
            O => \N__40866\,
            I => \N__40863\
        );

    \I__8216\ : Odrv4
    port map (
            O => \N__40863\,
            I => encoder0_position_scaled_9
        );

    \I__8215\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40857\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__40857\,
            I => n26_adj_697
        );

    \I__8213\ : InMux
    port map (
            O => \N__40854\,
            I => \bfn_11_29_0_\
        );

    \I__8212\ : InMux
    port map (
            O => \N__40851\,
            I => \N__40848\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__40848\,
            I => n25_adj_696
        );

    \I__8210\ : InMux
    port map (
            O => \N__40845\,
            I => n13087
        );

    \I__8209\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__40839\,
            I => n24_adj_695
        );

    \I__8207\ : InMux
    port map (
            O => \N__40836\,
            I => n13088
        );

    \I__8206\ : InMux
    port map (
            O => \N__40833\,
            I => \N__40830\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__40830\,
            I => \N__40827\
        );

    \I__8204\ : Span4Mux_v
    port map (
            O => \N__40827\,
            I => \N__40824\
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__40824\,
            I => encoder0_position_scaled_10
        );

    \I__8202\ : InMux
    port map (
            O => \N__40821\,
            I => \N__40818\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__40818\,
            I => \N__40815\
        );

    \I__8200\ : Span4Mux_v
    port map (
            O => \N__40815\,
            I => \N__40812\
        );

    \I__8199\ : Odrv4
    port map (
            O => \N__40812\,
            I => \pwm_setpoint_23_N_171_3\
        );

    \I__8198\ : InMux
    port map (
            O => \N__40809\,
            I => \N__40806\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__40806\,
            I => \N__40803\
        );

    \I__8196\ : Span4Mux_h
    port map (
            O => \N__40803\,
            I => \N__40800\
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__40800\,
            I => encoder0_position_scaled_11
        );

    \I__8194\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40794\
        );

    \I__8193\ : LocalMux
    port map (
            O => \N__40794\,
            I => \N__40791\
        );

    \I__8192\ : Span4Mux_h
    port map (
            O => \N__40791\,
            I => \N__40788\
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__40788\,
            I => \pwm_setpoint_23_N_171_13\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__40785\,
            I => \n15_adj_663_cascade_\
        );

    \I__8189\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40779\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__40779\,
            I => n15125
        );

    \I__8187\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40773\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__40773\,
            I => \N__40770\
        );

    \I__8185\ : Span4Mux_v
    port map (
            O => \N__40770\,
            I => \N__40767\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__40767\,
            I => encoder0_position_scaled_18
        );

    \I__8183\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40761\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__40761\,
            I => \N__40758\
        );

    \I__8181\ : Span4Mux_h
    port map (
            O => \N__40758\,
            I => \N__40755\
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__40755\,
            I => encoder0_position_scaled_20
        );

    \I__8179\ : InMux
    port map (
            O => \N__40752\,
            I => \N__40749\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__40749\,
            I => \N__40746\
        );

    \I__8177\ : Span4Mux_h
    port map (
            O => \N__40746\,
            I => \N__40743\
        );

    \I__8176\ : Odrv4
    port map (
            O => \N__40743\,
            I => encoder0_position_scaled_23
        );

    \I__8175\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40737\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__40737\,
            I => \N__40732\
        );

    \I__8173\ : InMux
    port map (
            O => \N__40736\,
            I => \N__40729\
        );

    \I__8172\ : InMux
    port map (
            O => \N__40735\,
            I => \N__40725\
        );

    \I__8171\ : Span4Mux_h
    port map (
            O => \N__40732\,
            I => \N__40722\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__40729\,
            I => \N__40719\
        );

    \I__8169\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40716\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__40725\,
            I => encoder0_position_29
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__40722\,
            I => encoder0_position_29
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__40719\,
            I => encoder0_position_29
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__40716\,
            I => encoder0_position_29
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__40707\,
            I => \N__40702\
        );

    \I__8163\ : InMux
    port map (
            O => \N__40706\,
            I => \N__40699\
        );

    \I__8162\ : InMux
    port map (
            O => \N__40705\,
            I => \N__40694\
        );

    \I__8161\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40694\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__40699\,
            I => n4
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__40694\,
            I => n4
        );

    \I__8158\ : CascadeMux
    port map (
            O => \N__40689\,
            I => \N__40685\
        );

    \I__8157\ : CascadeMux
    port map (
            O => \N__40688\,
            I => \N__40681\
        );

    \I__8156\ : InMux
    port map (
            O => \N__40685\,
            I => \N__40675\
        );

    \I__8155\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40675\
        );

    \I__8154\ : InMux
    port map (
            O => \N__40681\,
            I => \N__40670\
        );

    \I__8153\ : InMux
    port map (
            O => \N__40680\,
            I => \N__40670\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__40675\,
            I => n3
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__40670\,
            I => n3
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__40665\,
            I => \N__40660\
        );

    \I__8149\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40657\
        );

    \I__8148\ : CascadeMux
    port map (
            O => \N__40663\,
            I => \N__40654\
        );

    \I__8147\ : InMux
    port map (
            O => \N__40660\,
            I => \N__40650\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__40657\,
            I => \N__40647\
        );

    \I__8145\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40644\
        );

    \I__8144\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40641\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__40650\,
            I => encoder0_position_30
        );

    \I__8142\ : Odrv12
    port map (
            O => \N__40647\,
            I => encoder0_position_30
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__40644\,
            I => encoder0_position_30
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__40641\,
            I => encoder0_position_30
        );

    \I__8139\ : CascadeMux
    port map (
            O => \N__40632\,
            I => \n13642_cascade_\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__40629\,
            I => \N__40625\
        );

    \I__8137\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40622\
        );

    \I__8136\ : InMux
    port map (
            O => \N__40625\,
            I => \N__40619\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__40622\,
            I => \N__40615\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__40619\,
            I => \N__40612\
        );

    \I__8133\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40609\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__40615\,
            I => n829
        );

    \I__8131\ : Odrv12
    port map (
            O => \N__40612\,
            I => n829
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__40609\,
            I => n829
        );

    \I__8129\ : InMux
    port map (
            O => \N__40602\,
            I => \N__40599\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__40599\,
            I => \N__40596\
        );

    \I__8127\ : Span4Mux_v
    port map (
            O => \N__40596\,
            I => \N__40593\
        );

    \I__8126\ : Odrv4
    port map (
            O => \N__40593\,
            I => n32
        );

    \I__8125\ : InMux
    port map (
            O => \N__40590\,
            I => \N__40586\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__40589\,
            I => \N__40583\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__40586\,
            I => \N__40580\
        );

    \I__8122\ : InMux
    port map (
            O => \N__40583\,
            I => \N__40576\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__40580\,
            I => \N__40573\
        );

    \I__8120\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40570\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__40576\,
            I => encoder0_position_1
        );

    \I__8118\ : Odrv4
    port map (
            O => \N__40573\,
            I => encoder0_position_1
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__40570\,
            I => encoder0_position_1
        );

    \I__8116\ : CascadeMux
    port map (
            O => \N__40563\,
            I => \N__40560\
        );

    \I__8115\ : InMux
    port map (
            O => \N__40560\,
            I => \N__40555\
        );

    \I__8114\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40552\
        );

    \I__8113\ : InMux
    port map (
            O => \N__40558\,
            I => \N__40549\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__40555\,
            I => \N__40546\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__40552\,
            I => \N__40541\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__40549\,
            I => \N__40541\
        );

    \I__8109\ : Span4Mux_v
    port map (
            O => \N__40546\,
            I => \N__40538\
        );

    \I__8108\ : Span4Mux_v
    port map (
            O => \N__40541\,
            I => \N__40535\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__40538\,
            I => \N__40532\
        );

    \I__8106\ : Span4Mux_h
    port map (
            O => \N__40535\,
            I => \N__40529\
        );

    \I__8105\ : Odrv4
    port map (
            O => \N__40532\,
            I => n318
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__40529\,
            I => n318
        );

    \I__8103\ : InMux
    port map (
            O => \N__40524\,
            I => \N__40521\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__40521\,
            I => \N__40518\
        );

    \I__8101\ : Span4Mux_h
    port map (
            O => \N__40518\,
            I => \N__40515\
        );

    \I__8100\ : Odrv4
    port map (
            O => \N__40515\,
            I => encoder0_position_scaled_14
        );

    \I__8099\ : CascadeMux
    port map (
            O => \N__40512\,
            I => \n10_adj_606_cascade_\
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__40509\,
            I => \n15_adj_565_cascade_\
        );

    \I__8097\ : InMux
    port map (
            O => \N__40506\,
            I => \N__40503\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__40503\,
            I => n16_adj_564
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__40500\,
            I => \n13644_cascade_\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__40497\,
            I => \N__40494\
        );

    \I__8093\ : InMux
    port map (
            O => \N__40494\,
            I => \N__40490\
        );

    \I__8092\ : InMux
    port map (
            O => \N__40493\,
            I => \N__40486\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__40490\,
            I => \N__40483\
        );

    \I__8090\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40480\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__40486\,
            I => n830
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__40483\,
            I => n830
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__40480\,
            I => n830
        );

    \I__8086\ : InMux
    port map (
            O => \N__40473\,
            I => \N__40467\
        );

    \I__8085\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40467\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__40467\,
            I => n7
        );

    \I__8083\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40461\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__40461\,
            I => n5_adj_676
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__40458\,
            I => \n5_adj_676_cascade_\
        );

    \I__8080\ : CascadeMux
    port map (
            O => \N__40455\,
            I => \n13641_cascade_\
        );

    \I__8079\ : CascadeMux
    port map (
            O => \N__40452\,
            I => \n13646_cascade_\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__40449\,
            I => \N__40446\
        );

    \I__8077\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40443\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__40443\,
            I => \N__40438\
        );

    \I__8075\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40433\
        );

    \I__8074\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40433\
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__40438\,
            I => n831
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__40433\,
            I => n831
        );

    \I__8071\ : CascadeMux
    port map (
            O => \N__40428\,
            I => \N__40423\
        );

    \I__8070\ : InMux
    port map (
            O => \N__40427\,
            I => \N__40420\
        );

    \I__8069\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40417\
        );

    \I__8068\ : InMux
    port map (
            O => \N__40423\,
            I => \N__40413\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__40420\,
            I => \N__40408\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__40417\,
            I => \N__40408\
        );

    \I__8065\ : InMux
    port map (
            O => \N__40416\,
            I => \N__40405\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__40413\,
            I => encoder0_position_28
        );

    \I__8063\ : Odrv4
    port map (
            O => \N__40408\,
            I => encoder0_position_28
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__40405\,
            I => encoder0_position_28
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__40398\,
            I => \N__40394\
        );

    \I__8060\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40386\
        );

    \I__8059\ : InMux
    port map (
            O => \N__40394\,
            I => \N__40386\
        );

    \I__8058\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40386\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__40386\,
            I => n5
        );

    \I__8056\ : CascadeMux
    port map (
            O => \N__40383\,
            I => \n931_cascade_\
        );

    \I__8055\ : CascadeMux
    port map (
            O => \N__40380\,
            I => \N__40377\
        );

    \I__8054\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40374\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__40374\,
            I => n10
        );

    \I__8052\ : CascadeMux
    port map (
            O => \N__40371\,
            I => \N__40368\
        );

    \I__8051\ : InMux
    port map (
            O => \N__40368\,
            I => \N__40365\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__40365\,
            I => n897
        );

    \I__8049\ : CascadeMux
    port map (
            O => \N__40362\,
            I => \N__40359\
        );

    \I__8048\ : InMux
    port map (
            O => \N__40359\,
            I => \N__40356\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__40356\,
            I => \N__40352\
        );

    \I__8046\ : InMux
    port map (
            O => \N__40355\,
            I => \N__40348\
        );

    \I__8045\ : Span4Mux_h
    port map (
            O => \N__40352\,
            I => \N__40345\
        );

    \I__8044\ : InMux
    port map (
            O => \N__40351\,
            I => \N__40342\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__40348\,
            I => encoder0_position_25
        );

    \I__8042\ : Odrv4
    port map (
            O => \N__40345\,
            I => encoder0_position_25
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__40342\,
            I => encoder0_position_25
        );

    \I__8040\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40332\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__40332\,
            I => n8
        );

    \I__8038\ : CascadeMux
    port map (
            O => \N__40329\,
            I => \N__40324\
        );

    \I__8037\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40321\
        );

    \I__8036\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40318\
        );

    \I__8035\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40315\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__40321\,
            I => \N__40312\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__40318\,
            I => n294
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__40315\,
            I => n294
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__40312\,
            I => n294
        );

    \I__8030\ : CascadeMux
    port map (
            O => \N__40305\,
            I => \N__40302\
        );

    \I__8029\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40299\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__40299\,
            I => n14574
        );

    \I__8027\ : CascadeMux
    port map (
            O => \N__40296\,
            I => \N__40293\
        );

    \I__8026\ : InMux
    port map (
            O => \N__40293\,
            I => \N__40290\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__40290\,
            I => \N__40287\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__40287\,
            I => n828
        );

    \I__8023\ : CascadeMux
    port map (
            O => \N__40284\,
            I => \n828_cascade_\
        );

    \I__8022\ : InMux
    port map (
            O => \N__40281\,
            I => \N__40278\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__40278\,
            I => n12012
        );

    \I__8020\ : InMux
    port map (
            O => \N__40275\,
            I => \N__40270\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__40274\,
            I => \N__40267\
        );

    \I__8018\ : CascadeMux
    port map (
            O => \N__40273\,
            I => \N__40264\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__40270\,
            I => \N__40258\
        );

    \I__8016\ : InMux
    port map (
            O => \N__40267\,
            I => \N__40247\
        );

    \I__8015\ : InMux
    port map (
            O => \N__40264\,
            I => \N__40247\
        );

    \I__8014\ : InMux
    port map (
            O => \N__40263\,
            I => \N__40247\
        );

    \I__8013\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40247\
        );

    \I__8012\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40247\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__40258\,
            I => n861
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__40247\,
            I => n861
        );

    \I__8009\ : CascadeMux
    port map (
            O => \N__40242\,
            I => \n861_cascade_\
        );

    \I__8008\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40236\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__40236\,
            I => \N__40233\
        );

    \I__8006\ : Odrv4
    port map (
            O => \N__40233\,
            I => n898
        );

    \I__8005\ : InMux
    port map (
            O => \N__40230\,
            I => n12487
        );

    \I__8004\ : InMux
    port map (
            O => \N__40227\,
            I => n12488
        );

    \I__8003\ : InMux
    port map (
            O => \N__40224\,
            I => n12489
        );

    \I__8002\ : InMux
    port map (
            O => \N__40221\,
            I => n12490
        );

    \I__8001\ : InMux
    port map (
            O => \N__40218\,
            I => n12491
        );

    \I__8000\ : InMux
    port map (
            O => \N__40215\,
            I => n12492
        );

    \I__7999\ : CascadeMux
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__7998\ : InMux
    port map (
            O => \N__40209\,
            I => \N__40206\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__40206\,
            I => \N__40203\
        );

    \I__7996\ : Odrv12
    port map (
            O => \N__40203\,
            I => n901
        );

    \I__7995\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40197\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__40197\,
            I => n896
        );

    \I__7993\ : CascadeMux
    port map (
            O => \N__40194\,
            I => \N__40191\
        );

    \I__7992\ : InMux
    port map (
            O => \N__40191\,
            I => \N__40188\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__40188\,
            I => n900
        );

    \I__7990\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40182\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__40182\,
            I => n899
        );

    \I__7988\ : CascadeMux
    port map (
            O => \N__40179\,
            I => \n1820_cascade_\
        );

    \I__7987\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40173\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__40173\,
            I => \N__40170\
        );

    \I__7985\ : Odrv4
    port map (
            O => \N__40170\,
            I => n14538
        );

    \I__7984\ : CascadeMux
    port map (
            O => \N__40167\,
            I => \N__40164\
        );

    \I__7983\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40161\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__40161\,
            I => n30_adj_651
        );

    \I__7981\ : InMux
    port map (
            O => \N__40158\,
            I => \N__40155\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__40155\,
            I => n26
        );

    \I__7979\ : InMux
    port map (
            O => \N__40152\,
            I => \N__40148\
        );

    \I__7978\ : CascadeMux
    port map (
            O => \N__40151\,
            I => \N__40145\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__40148\,
            I => \N__40142\
        );

    \I__7976\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40138\
        );

    \I__7975\ : Span4Mux_h
    port map (
            O => \N__40142\,
            I => \N__40135\
        );

    \I__7974\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40132\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__40138\,
            I => encoder0_position_7
        );

    \I__7972\ : Odrv4
    port map (
            O => \N__40135\,
            I => encoder0_position_7
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__40132\,
            I => encoder0_position_7
        );

    \I__7970\ : InMux
    port map (
            O => \N__40125\,
            I => \N__40122\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__40122\,
            I => \N__40118\
        );

    \I__7968\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40114\
        );

    \I__7967\ : Span4Mux_v
    port map (
            O => \N__40118\,
            I => \N__40111\
        );

    \I__7966\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40108\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__40114\,
            I => \N__40105\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__40111\,
            I => \N__40100\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__40108\,
            I => \N__40100\
        );

    \I__7962\ : Span4Mux_h
    port map (
            O => \N__40105\,
            I => \N__40097\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__40100\,
            I => \N__40094\
        );

    \I__7960\ : Span4Mux_h
    port map (
            O => \N__40097\,
            I => \N__40091\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__40094\,
            I => n312
        );

    \I__7958\ : Odrv4
    port map (
            O => \N__40091\,
            I => n312
        );

    \I__7957\ : InMux
    port map (
            O => \N__40086\,
            I => \N__40083\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__40083\,
            I => n31
        );

    \I__7955\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40077\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__40077\,
            I => \N__40073\
        );

    \I__7953\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40069\
        );

    \I__7952\ : Span4Mux_h
    port map (
            O => \N__40073\,
            I => \N__40066\
        );

    \I__7951\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40063\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__40069\,
            I => encoder0_position_2
        );

    \I__7949\ : Odrv4
    port map (
            O => \N__40066\,
            I => encoder0_position_2
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__40063\,
            I => encoder0_position_2
        );

    \I__7947\ : InMux
    port map (
            O => \N__40056\,
            I => \N__40051\
        );

    \I__7946\ : InMux
    port map (
            O => \N__40055\,
            I => \N__40048\
        );

    \I__7945\ : InMux
    port map (
            O => \N__40054\,
            I => \N__40045\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__40051\,
            I => \N__40042\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__40048\,
            I => \N__40039\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__40045\,
            I => \N__40036\
        );

    \I__7941\ : Span4Mux_h
    port map (
            O => \N__40042\,
            I => \N__40033\
        );

    \I__7940\ : Span4Mux_v
    port map (
            O => \N__40039\,
            I => \N__40030\
        );

    \I__7939\ : Span4Mux_h
    port map (
            O => \N__40036\,
            I => \N__40027\
        );

    \I__7938\ : Span4Mux_v
    port map (
            O => \N__40033\,
            I => \N__40024\
        );

    \I__7937\ : Span4Mux_h
    port map (
            O => \N__40030\,
            I => \N__40021\
        );

    \I__7936\ : Span4Mux_v
    port map (
            O => \N__40027\,
            I => \N__40018\
        );

    \I__7935\ : Sp12to4
    port map (
            O => \N__40024\,
            I => \N__40015\
        );

    \I__7934\ : Odrv4
    port map (
            O => \N__40021\,
            I => n317
        );

    \I__7933\ : Odrv4
    port map (
            O => \N__40018\,
            I => n317
        );

    \I__7932\ : Odrv12
    port map (
            O => \N__40015\,
            I => n317
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__40008\,
            I => \N__40003\
        );

    \I__7930\ : InMux
    port map (
            O => \N__40007\,
            I => \N__40000\
        );

    \I__7929\ : InMux
    port map (
            O => \N__40006\,
            I => \N__39997\
        );

    \I__7928\ : InMux
    port map (
            O => \N__40003\,
            I => \N__39994\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__40000\,
            I => \N__39991\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__39997\,
            I => \N__39988\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__39994\,
            I => \N__39981\
        );

    \I__7924\ : Span4Mux_h
    port map (
            O => \N__39991\,
            I => \N__39981\
        );

    \I__7923\ : Span4Mux_v
    port map (
            O => \N__39988\,
            I => \N__39981\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__39981\,
            I => encoder0_position_10
        );

    \I__7921\ : CascadeMux
    port map (
            O => \N__39978\,
            I => \N__39975\
        );

    \I__7920\ : InMux
    port map (
            O => \N__39975\,
            I => \N__39972\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__39972\,
            I => n23_adj_644
        );

    \I__7918\ : InMux
    port map (
            O => \N__39969\,
            I => \N__39966\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__39966\,
            I => \N__39963\
        );

    \I__7916\ : Span4Mux_h
    port map (
            O => \N__39963\,
            I => \N__39960\
        );

    \I__7915\ : Odrv4
    port map (
            O => \N__39960\,
            I => encoder0_position_scaled_1
        );

    \I__7914\ : InMux
    port map (
            O => \N__39957\,
            I => \bfn_11_22_0_\
        );

    \I__7913\ : CascadeMux
    port map (
            O => \N__39954\,
            I => \N__39951\
        );

    \I__7912\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39947\
        );

    \I__7911\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39943\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__39947\,
            I => \N__39940\
        );

    \I__7909\ : InMux
    port map (
            O => \N__39946\,
            I => \N__39937\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__39943\,
            I => \N__39932\
        );

    \I__7907\ : Span4Mux_v
    port map (
            O => \N__39940\,
            I => \N__39932\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__39937\,
            I => n1931
        );

    \I__7905\ : Odrv4
    port map (
            O => \N__39932\,
            I => n1931
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__39927\,
            I => \N__39923\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__39926\,
            I => \N__39920\
        );

    \I__7902\ : InMux
    port map (
            O => \N__39923\,
            I => \N__39915\
        );

    \I__7901\ : InMux
    port map (
            O => \N__39920\,
            I => \N__39915\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__39915\,
            I => \N__39911\
        );

    \I__7899\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39908\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__39911\,
            I => n1918
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__39908\,
            I => n1918
        );

    \I__7896\ : CascadeMux
    port map (
            O => \N__39903\,
            I => \N__39900\
        );

    \I__7895\ : InMux
    port map (
            O => \N__39900\,
            I => \N__39897\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__39897\,
            I => n14520
        );

    \I__7893\ : CascadeMux
    port map (
            O => \N__39894\,
            I => \n14176_cascade_\
        );

    \I__7892\ : CascadeMux
    port map (
            O => \N__39891\,
            I => \n1752_cascade_\
        );

    \I__7891\ : InMux
    port map (
            O => \N__39888\,
            I => \N__39885\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__39885\,
            I => \N__39878\
        );

    \I__7889\ : CascadeMux
    port map (
            O => \N__39884\,
            I => \N__39875\
        );

    \I__7888\ : InMux
    port map (
            O => \N__39883\,
            I => \N__39869\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__39882\,
            I => \N__39864\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__39881\,
            I => \N__39861\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__39878\,
            I => \N__39856\
        );

    \I__7884\ : InMux
    port map (
            O => \N__39875\,
            I => \N__39853\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__39874\,
            I => \N__39849\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__39873\,
            I => \N__39846\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__39872\,
            I => \N__39842\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__39869\,
            I => \N__39835\
        );

    \I__7879\ : InMux
    port map (
            O => \N__39868\,
            I => \N__39830\
        );

    \I__7878\ : InMux
    port map (
            O => \N__39867\,
            I => \N__39830\
        );

    \I__7877\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39821\
        );

    \I__7876\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39821\
        );

    \I__7875\ : InMux
    port map (
            O => \N__39860\,
            I => \N__39821\
        );

    \I__7874\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39821\
        );

    \I__7873\ : Span4Mux_h
    port map (
            O => \N__39856\,
            I => \N__39816\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__39853\,
            I => \N__39816\
        );

    \I__7871\ : InMux
    port map (
            O => \N__39852\,
            I => \N__39807\
        );

    \I__7870\ : InMux
    port map (
            O => \N__39849\,
            I => \N__39807\
        );

    \I__7869\ : InMux
    port map (
            O => \N__39846\,
            I => \N__39807\
        );

    \I__7868\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39807\
        );

    \I__7867\ : InMux
    port map (
            O => \N__39842\,
            I => \N__39802\
        );

    \I__7866\ : InMux
    port map (
            O => \N__39841\,
            I => \N__39802\
        );

    \I__7865\ : InMux
    port map (
            O => \N__39840\,
            I => \N__39795\
        );

    \I__7864\ : InMux
    port map (
            O => \N__39839\,
            I => \N__39795\
        );

    \I__7863\ : InMux
    port map (
            O => \N__39838\,
            I => \N__39795\
        );

    \I__7862\ : Odrv12
    port map (
            O => \N__39835\,
            I => n1851
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__39830\,
            I => n1851
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__39821\,
            I => n1851
        );

    \I__7859\ : Odrv4
    port map (
            O => \N__39816\,
            I => n1851
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__39807\,
            I => n1851
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__39802\,
            I => n1851
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__39795\,
            I => n1851
        );

    \I__7855\ : InMux
    port map (
            O => \N__39780\,
            I => \N__39777\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__39777\,
            I => \N__39774\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__39774\,
            I => \N__39771\
        );

    \I__7852\ : Span4Mux_v
    port map (
            O => \N__39771\,
            I => \N__39768\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__39768\,
            I => n15644
        );

    \I__7850\ : CascadeMux
    port map (
            O => \N__39765\,
            I => \n1832_cascade_\
        );

    \I__7849\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39759\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__39759\,
            I => \N__39756\
        );

    \I__7847\ : Odrv4
    port map (
            O => \N__39756\,
            I => n11968
        );

    \I__7846\ : CascadeMux
    port map (
            O => \N__39753\,
            I => \n1819_cascade_\
        );

    \I__7845\ : InMux
    port map (
            O => \N__39750\,
            I => \N__39747\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__39747\,
            I => n14532
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__39744\,
            I => \n1851_cascade_\
        );

    \I__7842\ : InMux
    port map (
            O => \N__39741\,
            I => \N__39738\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__39738\,
            I => \N__39734\
        );

    \I__7840\ : InMux
    port map (
            O => \N__39737\,
            I => \N__39731\
        );

    \I__7839\ : Span4Mux_v
    port map (
            O => \N__39734\,
            I => \N__39725\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__39731\,
            I => \N__39725\
        );

    \I__7837\ : InMux
    port map (
            O => \N__39730\,
            I => \N__39722\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__39725\,
            I => n1920
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__39722\,
            I => n1920
        );

    \I__7834\ : InMux
    port map (
            O => \N__39717\,
            I => \N__39713\
        );

    \I__7833\ : InMux
    port map (
            O => \N__39716\,
            I => \N__39710\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__39713\,
            I => \N__39707\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__39710\,
            I => \N__39704\
        );

    \I__7830\ : Span4Mux_h
    port map (
            O => \N__39707\,
            I => \N__39698\
        );

    \I__7829\ : Span4Mux_v
    port map (
            O => \N__39704\,
            I => \N__39698\
        );

    \I__7828\ : InMux
    port map (
            O => \N__39703\,
            I => \N__39695\
        );

    \I__7827\ : Odrv4
    port map (
            O => \N__39698\,
            I => n1919
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__39695\,
            I => n1919
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__39690\,
            I => \N__39687\
        );

    \I__7824\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39683\
        );

    \I__7823\ : InMux
    port map (
            O => \N__39686\,
            I => \N__39680\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__39683\,
            I => \N__39677\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__39680\,
            I => \N__39674\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__39677\,
            I => \N__39671\
        );

    \I__7819\ : Odrv4
    port map (
            O => \N__39674\,
            I => n1930
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__39671\,
            I => n1930
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__39666\,
            I => \n1930_cascade_\
        );

    \I__7816\ : CascadeMux
    port map (
            O => \N__39663\,
            I => \N__39659\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__39662\,
            I => \N__39656\
        );

    \I__7814\ : InMux
    port map (
            O => \N__39659\,
            I => \N__39653\
        );

    \I__7813\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39649\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__39653\,
            I => \N__39646\
        );

    \I__7811\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39643\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__39649\,
            I => \N__39640\
        );

    \I__7809\ : Span4Mux_h
    port map (
            O => \N__39646\,
            I => \N__39635\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__39643\,
            I => \N__39635\
        );

    \I__7807\ : Odrv4
    port map (
            O => \N__39640\,
            I => n1929
        );

    \I__7806\ : Odrv4
    port map (
            O => \N__39635\,
            I => n1929
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__39630\,
            I => \N__39627\
        );

    \I__7804\ : InMux
    port map (
            O => \N__39627\,
            I => \N__39624\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__39624\,
            I => n14540
        );

    \I__7802\ : CascadeMux
    port map (
            O => \N__39621\,
            I => \n1826_cascade_\
        );

    \I__7801\ : CascadeMux
    port map (
            O => \N__39618\,
            I => \N__39614\
        );

    \I__7800\ : CascadeMux
    port map (
            O => \N__39617\,
            I => \N__39611\
        );

    \I__7799\ : InMux
    port map (
            O => \N__39614\,
            I => \N__39608\
        );

    \I__7798\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39604\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__39608\,
            I => \N__39601\
        );

    \I__7796\ : InMux
    port map (
            O => \N__39607\,
            I => \N__39598\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__39604\,
            I => n1928
        );

    \I__7794\ : Odrv4
    port map (
            O => \N__39601\,
            I => n1928
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__39598\,
            I => n1928
        );

    \I__7792\ : InMux
    port map (
            O => \N__39591\,
            I => \N__39588\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__39588\,
            I => n14526
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__39585\,
            I => \n14530_cascade_\
        );

    \I__7789\ : InMux
    port map (
            O => \N__39582\,
            I => \N__39579\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__39579\,
            I => n11_adj_591
        );

    \I__7787\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39573\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__39573\,
            I => \pwm_setpoint_23_N_171_18\
        );

    \I__7785\ : InMux
    port map (
            O => \N__39570\,
            I => \N__39567\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__39567\,
            I => n3_adj_583
        );

    \I__7783\ : InMux
    port map (
            O => \N__39564\,
            I => \N__39561\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__39561\,
            I => n9_adj_589
        );

    \I__7781\ : InMux
    port map (
            O => \N__39558\,
            I => \N__39555\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__39555\,
            I => \N__39551\
        );

    \I__7779\ : InMux
    port map (
            O => \N__39554\,
            I => \N__39548\
        );

    \I__7778\ : Odrv12
    port map (
            O => \N__39551\,
            I => \reg_B_2\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__39548\,
            I => \reg_B_2\
        );

    \I__7776\ : InMux
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__39540\,
            I => \N__39536\
        );

    \I__7774\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39533\
        );

    \I__7773\ : Span4Mux_s2_h
    port map (
            O => \N__39536\,
            I => \N__39530\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__39533\,
            I => \N__39527\
        );

    \I__7771\ : Span4Mux_v
    port map (
            O => \N__39530\,
            I => \N__39523\
        );

    \I__7770\ : Span4Mux_v
    port map (
            O => \N__39527\,
            I => \N__39520\
        );

    \I__7769\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39517\
        );

    \I__7768\ : Span4Mux_v
    port map (
            O => \N__39523\,
            I => \N__39513\
        );

    \I__7767\ : Sp12to4
    port map (
            O => \N__39520\,
            I => \N__39508\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__39517\,
            I => \N__39508\
        );

    \I__7765\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39505\
        );

    \I__7764\ : Odrv4
    port map (
            O => \N__39513\,
            I => n14125
        );

    \I__7763\ : Odrv12
    port map (
            O => \N__39508\,
            I => n14125
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__39505\,
            I => n14125
        );

    \I__7761\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39495\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__39495\,
            I => n14937
        );

    \I__7759\ : CascadeMux
    port map (
            O => \N__39492\,
            I => \n14936_cascade_\
        );

    \I__7758\ : IoInMux
    port map (
            O => \N__39489\,
            I => \N__39486\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__39486\,
            I => \N__39483\
        );

    \I__7756\ : Span4Mux_s0_v
    port map (
            O => \N__39483\,
            I => \N__39480\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__39480\,
            I => \N__39477\
        );

    \I__7754\ : Odrv4
    port map (
            O => \N__39477\,
            I => \LED_c\
        );

    \I__7753\ : InMux
    port map (
            O => \N__39474\,
            I => \N__39471\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__39471\,
            I => \pwm_setpoint_23_N_171_22\
        );

    \I__7751\ : InMux
    port map (
            O => \N__39468\,
            I => \N__39465\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__39465\,
            I => n19_adj_599
        );

    \I__7749\ : InMux
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__39459\,
            I => \pwm_setpoint_23_N_171_6\
        );

    \I__7747\ : InMux
    port map (
            O => \N__39456\,
            I => \N__39453\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__39453\,
            I => \pwm_setpoint_23_N_171_10\
        );

    \I__7745\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39447\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__39447\,
            I => \pwm_setpoint_23_N_171_9\
        );

    \I__7743\ : InMux
    port map (
            O => \N__39444\,
            I => \N__39441\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__39441\,
            I => \pwm_setpoint_23_N_171_4\
        );

    \I__7741\ : InMux
    port map (
            O => \N__39438\,
            I => \N__39435\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__39435\,
            I => n7_adj_587
        );

    \I__7739\ : InMux
    port map (
            O => \N__39432\,
            I => \N__39429\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__39429\,
            I => \pwm_setpoint_23_N_171_15\
        );

    \I__7737\ : InMux
    port map (
            O => \N__39426\,
            I => \N__39422\
        );

    \I__7736\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39419\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__39422\,
            I => \N__39416\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39413\
        );

    \I__7733\ : Span4Mux_v
    port map (
            O => \N__39416\,
            I => \N__39410\
        );

    \I__7732\ : Span12Mux_s3_v
    port map (
            O => \N__39413\,
            I => \N__39407\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__39410\,
            I => \N__39404\
        );

    \I__7730\ : Odrv12
    port map (
            O => \N__39407\,
            I => \reg_B_1\
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__39404\,
            I => \reg_B_1\
        );

    \I__7728\ : InMux
    port map (
            O => \N__39399\,
            I => \N__39396\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__39396\,
            I => \N__39392\
        );

    \I__7726\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39389\
        );

    \I__7725\ : Odrv4
    port map (
            O => \N__39392\,
            I => pwm_setpoint_15
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__39389\,
            I => pwm_setpoint_15
        );

    \I__7723\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39379\
        );

    \I__7722\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39374\
        );

    \I__7721\ : InMux
    port map (
            O => \N__39382\,
            I => \N__39374\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__39379\,
            I => \N__39369\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__39374\,
            I => \N__39369\
        );

    \I__7718\ : Odrv12
    port map (
            O => \N__39369\,
            I => n31_adj_674
        );

    \I__7717\ : InMux
    port map (
            O => \N__39366\,
            I => \N__39363\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__39363\,
            I => n15121
        );

    \I__7715\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39357\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__39357\,
            I => n15182
        );

    \I__7713\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39351\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__39351\,
            I => \N__39347\
        );

    \I__7711\ : InMux
    port map (
            O => \N__39350\,
            I => \N__39344\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__39347\,
            I => n29_adj_672
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__39344\,
            I => n29_adj_672
        );

    \I__7708\ : CascadeMux
    port map (
            O => \N__39339\,
            I => \n30_adj_673_cascade_\
        );

    \I__7707\ : InMux
    port map (
            O => \N__39336\,
            I => \N__39333\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__39333\,
            I => n10_adj_659
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__39330\,
            I => \N__39327\
        );

    \I__7704\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39324\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__39324\,
            I => n15267
        );

    \I__7702\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39318\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__39318\,
            I => n20_adj_600
        );

    \I__7700\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39312\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__39312\,
            I => n16_adj_596
        );

    \I__7698\ : InMux
    port map (
            O => \N__39309\,
            I => \N__39306\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__39306\,
            I => n15_adj_595
        );

    \I__7696\ : InMux
    port map (
            O => \N__39303\,
            I => \N__39300\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__39300\,
            I => n21_adj_601
        );

    \I__7694\ : InMux
    port map (
            O => \N__39297\,
            I => \N__39294\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__39294\,
            I => \pwm_setpoint_23_N_171_5\
        );

    \I__7692\ : CascadeMux
    port map (
            O => \N__39291\,
            I => \n29_adj_672_cascade_\
        );

    \I__7691\ : InMux
    port map (
            O => \N__39288\,
            I => \N__39285\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__39285\,
            I => n15233
        );

    \I__7689\ : InMux
    port map (
            O => \N__39282\,
            I => \N__39279\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__39279\,
            I => n15234
        );

    \I__7687\ : InMux
    port map (
            O => \N__39276\,
            I => \N__39273\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__39273\,
            I => \N__39270\
        );

    \I__7685\ : Span4Mux_v
    port map (
            O => \N__39270\,
            I => \N__39267\
        );

    \I__7684\ : Odrv4
    port map (
            O => \N__39267\,
            I => encoder0_position_scaled_16
        );

    \I__7683\ : CascadeMux
    port map (
            O => \N__39264\,
            I => \n33_adj_675_cascade_\
        );

    \I__7682\ : InMux
    port map (
            O => \N__39261\,
            I => \N__39258\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__39258\,
            I => \N__39255\
        );

    \I__7680\ : Odrv4
    port map (
            O => \N__39255\,
            I => n12_adj_592
        );

    \I__7679\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39249\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__39249\,
            I => \N__39246\
        );

    \I__7677\ : Span4Mux_h
    port map (
            O => \N__39246\,
            I => \N__39243\
        );

    \I__7676\ : Odrv4
    port map (
            O => \N__39243\,
            I => \pwm_setpoint_23_N_171_16\
        );

    \I__7675\ : CascadeMux
    port map (
            O => \N__39240\,
            I => \N__39237\
        );

    \I__7674\ : InMux
    port map (
            O => \N__39237\,
            I => \N__39234\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__39234\,
            I => \N__39231\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__39231\,
            I => \pwm_setpoint_23_N_171_2\
        );

    \I__7671\ : CascadeMux
    port map (
            O => \N__39228\,
            I => \N__39225\
        );

    \I__7670\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39222\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__39222\,
            I => \N__39219\
        );

    \I__7668\ : Span4Mux_v
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__7667\ : Odrv4
    port map (
            O => \N__39216\,
            I => \pwm_setpoint_23_N_171_14\
        );

    \I__7666\ : InMux
    port map (
            O => \N__39213\,
            I => \N__39207\
        );

    \I__7665\ : InMux
    port map (
            O => \N__39212\,
            I => \N__39207\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__39207\,
            I => \N__39204\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__39204\,
            I => pwm_setpoint_14
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__39201\,
            I => \N__39198\
        );

    \I__7661\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39195\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__7659\ : Odrv4
    port map (
            O => \N__39192\,
            I => n3_adj_624
        );

    \I__7658\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39186\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__7656\ : Span4Mux_h
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__7655\ : Odrv4
    port map (
            O => \N__39180\,
            I => encoder0_position_scaled_2
        );

    \I__7654\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__39174\,
            I => n4_adj_655
        );

    \I__7652\ : CascadeMux
    port map (
            O => \N__39171\,
            I => \N__39168\
        );

    \I__7651\ : InMux
    port map (
            O => \N__39168\,
            I => \N__39165\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__39165\,
            I => \quad_counter0.a_prev_N_543\
        );

    \I__7649\ : InMux
    port map (
            O => \N__39162\,
            I => \N__39152\
        );

    \I__7648\ : InMux
    port map (
            O => \N__39161\,
            I => \N__39152\
        );

    \I__7647\ : InMux
    port map (
            O => \N__39160\,
            I => \N__39152\
        );

    \I__7646\ : InMux
    port map (
            O => \N__39159\,
            I => \N__39149\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__39152\,
            I => \quad_counter0.b_new_1\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__39149\,
            I => \quad_counter0.b_new_1\
        );

    \I__7643\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39138\
        );

    \I__7642\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39138\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__39138\,
            I => \quad_counter0.a_prev\
        );

    \I__7640\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39130\
        );

    \I__7639\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39125\
        );

    \I__7638\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39125\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__39130\,
            I => \quad_counter0.debounce_cnt\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__39125\,
            I => \quad_counter0.debounce_cnt\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__39120\,
            I => \quad_counter0.direction_N_540_cascade_\
        );

    \I__7634\ : CEMux
    port map (
            O => \N__39117\,
            I => \N__39114\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__39114\,
            I => \N__39108\
        );

    \I__7632\ : CEMux
    port map (
            O => \N__39113\,
            I => \N__39105\
        );

    \I__7631\ : CEMux
    port map (
            O => \N__39112\,
            I => \N__39102\
        );

    \I__7630\ : CEMux
    port map (
            O => \N__39111\,
            I => \N__39099\
        );

    \I__7629\ : Span4Mux_h
    port map (
            O => \N__39108\,
            I => \N__39092\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__39105\,
            I => \N__39092\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__39102\,
            I => \N__39092\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__39099\,
            I => \N__39089\
        );

    \I__7625\ : Span4Mux_v
    port map (
            O => \N__39092\,
            I => \N__39086\
        );

    \I__7624\ : Odrv4
    port map (
            O => \N__39089\,
            I => \direction_N_537\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__39086\,
            I => \direction_N_537\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__39081\,
            I => \N__39077\
        );

    \I__7621\ : CascadeMux
    port map (
            O => \N__39080\,
            I => \N__39071\
        );

    \I__7620\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39067\
        );

    \I__7619\ : InMux
    port map (
            O => \N__39076\,
            I => \N__39060\
        );

    \I__7618\ : InMux
    port map (
            O => \N__39075\,
            I => \N__39060\
        );

    \I__7617\ : InMux
    port map (
            O => \N__39074\,
            I => \N__39060\
        );

    \I__7616\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39055\
        );

    \I__7615\ : InMux
    port map (
            O => \N__39070\,
            I => \N__39055\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__39067\,
            I => a_new_1
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__39060\,
            I => a_new_1
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__39055\,
            I => a_new_1
        );

    \I__7611\ : CascadeMux
    port map (
            O => \N__39048\,
            I => \direction_N_537_cascade_\
        );

    \I__7610\ : InMux
    port map (
            O => \N__39045\,
            I => \N__39039\
        );

    \I__7609\ : InMux
    port map (
            O => \N__39044\,
            I => \N__39034\
        );

    \I__7608\ : InMux
    port map (
            O => \N__39043\,
            I => \N__39034\
        );

    \I__7607\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39031\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__39039\,
            I => b_prev
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__39034\,
            I => b_prev
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__39031\,
            I => b_prev
        );

    \I__7603\ : InMux
    port map (
            O => \N__39024\,
            I => \N__39021\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__39021\,
            I => n1302
        );

    \I__7601\ : CascadeMux
    port map (
            O => \N__39018\,
            I => \N__39015\
        );

    \I__7600\ : InMux
    port map (
            O => \N__39015\,
            I => \N__39012\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__39012\,
            I => n4_adj_625
        );

    \I__7598\ : InMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__39006\,
            I => pwm_setpoint_1
        );

    \I__7596\ : InMux
    port map (
            O => \N__39003\,
            I => \N__39000\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__39000\,
            I => pwm_setpoint_0
        );

    \I__7594\ : InMux
    port map (
            O => \N__38997\,
            I => \N__38994\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__38994\,
            I => \N__38991\
        );

    \I__7592\ : Odrv12
    port map (
            O => \N__38991\,
            I => n28
        );

    \I__7591\ : InMux
    port map (
            O => \N__38988\,
            I => \N__38984\
        );

    \I__7590\ : CascadeMux
    port map (
            O => \N__38987\,
            I => \N__38981\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__38984\,
            I => \N__38978\
        );

    \I__7588\ : InMux
    port map (
            O => \N__38981\,
            I => \N__38974\
        );

    \I__7587\ : Span4Mux_v
    port map (
            O => \N__38978\,
            I => \N__38971\
        );

    \I__7586\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38968\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__38974\,
            I => encoder0_position_5
        );

    \I__7584\ : Odrv4
    port map (
            O => \N__38971\,
            I => encoder0_position_5
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__38968\,
            I => encoder0_position_5
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__38961\,
            I => \N__38958\
        );

    \I__7581\ : InMux
    port map (
            O => \N__38958\,
            I => \N__38953\
        );

    \I__7580\ : InMux
    port map (
            O => \N__38957\,
            I => \N__38950\
        );

    \I__7579\ : InMux
    port map (
            O => \N__38956\,
            I => \N__38947\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__38953\,
            I => \N__38942\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__38950\,
            I => \N__38942\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__38947\,
            I => \N__38937\
        );

    \I__7575\ : Span4Mux_v
    port map (
            O => \N__38942\,
            I => \N__38937\
        );

    \I__7574\ : Span4Mux_h
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__7573\ : Span4Mux_h
    port map (
            O => \N__38934\,
            I => \N__38931\
        );

    \I__7572\ : Odrv4
    port map (
            O => \N__38931\,
            I => n314
        );

    \I__7571\ : InMux
    port map (
            O => \N__38928\,
            I => \N__38923\
        );

    \I__7570\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38920\
        );

    \I__7569\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38917\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__38923\,
            I => \N__38914\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__38920\,
            I => \N__38909\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__38917\,
            I => \N__38909\
        );

    \I__7565\ : Span4Mux_v
    port map (
            O => \N__38914\,
            I => \N__38906\
        );

    \I__7564\ : Span4Mux_h
    port map (
            O => \N__38909\,
            I => \N__38903\
        );

    \I__7563\ : Span4Mux_h
    port map (
            O => \N__38906\,
            I => \N__38900\
        );

    \I__7562\ : Span4Mux_h
    port map (
            O => \N__38903\,
            I => \N__38897\
        );

    \I__7561\ : Odrv4
    port map (
            O => \N__38900\,
            I => \quad_counter0.b_new_0\
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__38897\,
            I => \quad_counter0.b_new_0\
        );

    \I__7559\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38889\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__38889\,
            I => \N__38886\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__38886\,
            I => \N__38883\
        );

    \I__7556\ : Odrv4
    port map (
            O => \N__38883\,
            I => encoder0_position_scaled_0
        );

    \I__7555\ : InMux
    port map (
            O => \N__38880\,
            I => \N__38877\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__38877\,
            I => \N__38874\
        );

    \I__7553\ : Span4Mux_v
    port map (
            O => \N__38874\,
            I => \N__38871\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__38871\,
            I => encoder0_position_scaled_15
        );

    \I__7551\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38865\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__38865\,
            I => \N__38862\
        );

    \I__7549\ : Span4Mux_h
    port map (
            O => \N__38862\,
            I => \N__38859\
        );

    \I__7548\ : Odrv4
    port map (
            O => \N__38859\,
            I => encoder0_position_scaled_13
        );

    \I__7547\ : InMux
    port map (
            O => \N__38856\,
            I => n12994
        );

    \I__7546\ : InMux
    port map (
            O => \N__38853\,
            I => n12995
        );

    \I__7545\ : InMux
    port map (
            O => \N__38850\,
            I => n12996
        );

    \I__7544\ : InMux
    port map (
            O => \N__38847\,
            I => n12997
        );

    \I__7543\ : InMux
    port map (
            O => \N__38844\,
            I => n12998
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__7541\ : InMux
    port map (
            O => \N__38838\,
            I => \N__38835\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__38835\,
            I => n5_adj_626
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__38832\,
            I => \N__38829\
        );

    \I__7538\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38826\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__38826\,
            I => n6_adj_627
        );

    \I__7536\ : CascadeMux
    port map (
            O => \N__38823\,
            I => \N__38820\
        );

    \I__7535\ : InMux
    port map (
            O => \N__38820\,
            I => \N__38817\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__38817\,
            I => n8_adj_629
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__38814\,
            I => \N__38811\
        );

    \I__7532\ : InMux
    port map (
            O => \N__38811\,
            I => \N__38808\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__38808\,
            I => n7_adj_628
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__38805\,
            I => \N__38802\
        );

    \I__7529\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38799\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38796\
        );

    \I__7527\ : Odrv4
    port map (
            O => \N__38796\,
            I => n15_adj_636
        );

    \I__7526\ : InMux
    port map (
            O => \N__38793\,
            I => n12985
        );

    \I__7525\ : InMux
    port map (
            O => \N__38790\,
            I => n12986
        );

    \I__7524\ : CascadeMux
    port map (
            O => \N__38787\,
            I => \N__38784\
        );

    \I__7523\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38781\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__38781\,
            I => \N__38778\
        );

    \I__7521\ : Odrv4
    port map (
            O => \N__38778\,
            I => n13_adj_634
        );

    \I__7520\ : InMux
    port map (
            O => \N__38775\,
            I => n12987
        );

    \I__7519\ : InMux
    port map (
            O => \N__38772\,
            I => n12988
        );

    \I__7518\ : InMux
    port map (
            O => \N__38769\,
            I => n12989
        );

    \I__7517\ : InMux
    port map (
            O => \N__38766\,
            I => n12990
        );

    \I__7516\ : InMux
    port map (
            O => \N__38763\,
            I => \bfn_10_24_0_\
        );

    \I__7515\ : InMux
    port map (
            O => \N__38760\,
            I => n12992
        );

    \I__7514\ : InMux
    port map (
            O => \N__38757\,
            I => n12993
        );

    \I__7513\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38751\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__38751\,
            I => \N__38748\
        );

    \I__7511\ : Span4Mux_h
    port map (
            O => \N__38748\,
            I => \N__38745\
        );

    \I__7510\ : Span4Mux_h
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__7509\ : Odrv4
    port map (
            O => \N__38742\,
            I => n23
        );

    \I__7508\ : InMux
    port map (
            O => \N__38739\,
            I => n12977
        );

    \I__7507\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38733\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__38733\,
            I => \N__38730\
        );

    \I__7505\ : Odrv4
    port map (
            O => \N__38730\,
            I => n22_adj_643
        );

    \I__7504\ : InMux
    port map (
            O => \N__38727\,
            I => \N__38724\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__38724\,
            I => \N__38721\
        );

    \I__7502\ : Odrv4
    port map (
            O => \N__38721\,
            I => n22
        );

    \I__7501\ : InMux
    port map (
            O => \N__38718\,
            I => n12978
        );

    \I__7500\ : CascadeMux
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__7499\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38709\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__38709\,
            I => \N__38706\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__38706\,
            I => \N__38703\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__38703\,
            I => \N__38700\
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__38700\,
            I => n21_adj_642
        );

    \I__7494\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__38694\,
            I => \N__38691\
        );

    \I__7492\ : Span4Mux_h
    port map (
            O => \N__38691\,
            I => \N__38688\
        );

    \I__7491\ : Span4Mux_h
    port map (
            O => \N__38688\,
            I => \N__38685\
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__38685\,
            I => n21
        );

    \I__7489\ : InMux
    port map (
            O => \N__38682\,
            I => n12979
        );

    \I__7488\ : CascadeMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__7487\ : InMux
    port map (
            O => \N__38676\,
            I => \N__38673\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__38673\,
            I => \N__38670\
        );

    \I__7485\ : Span4Mux_h
    port map (
            O => \N__38670\,
            I => \N__38667\
        );

    \I__7484\ : Span4Mux_h
    port map (
            O => \N__38667\,
            I => \N__38664\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__38664\,
            I => n20_adj_641
        );

    \I__7482\ : InMux
    port map (
            O => \N__38661\,
            I => \N__38658\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__38658\,
            I => \N__38655\
        );

    \I__7480\ : Span4Mux_v
    port map (
            O => \N__38655\,
            I => \N__38652\
        );

    \I__7479\ : Span4Mux_h
    port map (
            O => \N__38652\,
            I => \N__38649\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__38649\,
            I => n20
        );

    \I__7477\ : InMux
    port map (
            O => \N__38646\,
            I => n12980
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__38643\,
            I => \N__38640\
        );

    \I__7475\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38637\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__38637\,
            I => \N__38634\
        );

    \I__7473\ : Span4Mux_h
    port map (
            O => \N__38634\,
            I => \N__38631\
        );

    \I__7472\ : Odrv4
    port map (
            O => \N__38631\,
            I => n19_adj_640
        );

    \I__7471\ : InMux
    port map (
            O => \N__38628\,
            I => \N__38625\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__38625\,
            I => \N__38622\
        );

    \I__7469\ : Span4Mux_v
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__7468\ : Odrv4
    port map (
            O => \N__38619\,
            I => n19
        );

    \I__7467\ : InMux
    port map (
            O => \N__38616\,
            I => n12981
        );

    \I__7466\ : InMux
    port map (
            O => \N__38613\,
            I => n12982
        );

    \I__7465\ : CascadeMux
    port map (
            O => \N__38610\,
            I => \N__38607\
        );

    \I__7464\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38604\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__38604\,
            I => \N__38601\
        );

    \I__7462\ : Odrv12
    port map (
            O => \N__38601\,
            I => n17_adj_638
        );

    \I__7461\ : InMux
    port map (
            O => \N__38598\,
            I => \bfn_10_23_0_\
        );

    \I__7460\ : InMux
    port map (
            O => \N__38595\,
            I => n12984
        );

    \I__7459\ : CascadeMux
    port map (
            O => \N__38592\,
            I => \N__38589\
        );

    \I__7458\ : InMux
    port map (
            O => \N__38589\,
            I => \N__38586\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__38586\,
            I => n31_adj_652
        );

    \I__7456\ : InMux
    port map (
            O => \N__38583\,
            I => n12969
        );

    \I__7455\ : InMux
    port map (
            O => \N__38580\,
            I => n12970
        );

    \I__7454\ : CascadeMux
    port map (
            O => \N__38577\,
            I => \N__38574\
        );

    \I__7453\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38571\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__38571\,
            I => n29_adj_650
        );

    \I__7451\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38565\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__38565\,
            I => \N__38562\
        );

    \I__7449\ : Span4Mux_v
    port map (
            O => \N__38562\,
            I => \N__38559\
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__38559\,
            I => n29
        );

    \I__7447\ : InMux
    port map (
            O => \N__38556\,
            I => n12971
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__38553\,
            I => \N__38550\
        );

    \I__7445\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38547\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__38547\,
            I => n28_adj_649
        );

    \I__7443\ : InMux
    port map (
            O => \N__38544\,
            I => n12972
        );

    \I__7442\ : CascadeMux
    port map (
            O => \N__38541\,
            I => \N__38538\
        );

    \I__7441\ : InMux
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__38535\,
            I => n27_adj_648
        );

    \I__7439\ : InMux
    port map (
            O => \N__38532\,
            I => n12973
        );

    \I__7438\ : CascadeMux
    port map (
            O => \N__38529\,
            I => \N__38526\
        );

    \I__7437\ : InMux
    port map (
            O => \N__38526\,
            I => \N__38523\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__38523\,
            I => n26_adj_647
        );

    \I__7435\ : InMux
    port map (
            O => \N__38520\,
            I => n12974
        );

    \I__7434\ : CascadeMux
    port map (
            O => \N__38517\,
            I => \N__38514\
        );

    \I__7433\ : InMux
    port map (
            O => \N__38514\,
            I => \N__38511\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__38511\,
            I => \N__38508\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__38508\,
            I => \N__38505\
        );

    \I__7430\ : Span4Mux_h
    port map (
            O => \N__38505\,
            I => \N__38502\
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__38502\,
            I => n25_adj_646
        );

    \I__7428\ : InMux
    port map (
            O => \N__38499\,
            I => \N__38496\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__38496\,
            I => \N__38493\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__38493\,
            I => \N__38490\
        );

    \I__7425\ : Span4Mux_h
    port map (
            O => \N__38490\,
            I => \N__38487\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__38487\,
            I => n25_adj_551
        );

    \I__7423\ : InMux
    port map (
            O => \N__38484\,
            I => \bfn_10_22_0_\
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__38481\,
            I => \N__38478\
        );

    \I__7421\ : InMux
    port map (
            O => \N__38478\,
            I => \N__38475\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__38475\,
            I => \N__38472\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__38472\,
            I => n24_adj_645
        );

    \I__7418\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38466\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__38466\,
            I => \N__38463\
        );

    \I__7416\ : Odrv12
    port map (
            O => \N__38463\,
            I => n24
        );

    \I__7415\ : InMux
    port map (
            O => \N__38460\,
            I => n12976
        );

    \I__7414\ : CascadeMux
    port map (
            O => \N__38457\,
            I => \N__38453\
        );

    \I__7413\ : InMux
    port map (
            O => \N__38456\,
            I => \N__38450\
        );

    \I__7412\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38447\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__38450\,
            I => \N__38444\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__38447\,
            I => n1932
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__38444\,
            I => n1932
        );

    \I__7408\ : CascadeMux
    port map (
            O => \N__38439\,
            I => \n1932_cascade_\
        );

    \I__7407\ : InMux
    port map (
            O => \N__38436\,
            I => \N__38433\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__38433\,
            I => \N__38430\
        );

    \I__7405\ : Odrv4
    port map (
            O => \N__38430\,
            I => n1999
        );

    \I__7404\ : CascadeMux
    port map (
            O => \N__38427\,
            I => \N__38424\
        );

    \I__7403\ : InMux
    port map (
            O => \N__38424\,
            I => \N__38420\
        );

    \I__7402\ : InMux
    port map (
            O => \N__38423\,
            I => \N__38417\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__38420\,
            I => \N__38414\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__38417\,
            I => \N__38411\
        );

    \I__7399\ : Span4Mux_h
    port map (
            O => \N__38414\,
            I => \N__38408\
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__38411\,
            I => n2031
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__38408\,
            I => n2031
        );

    \I__7396\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38399\
        );

    \I__7395\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38395\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__38399\,
            I => \N__38392\
        );

    \I__7393\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38389\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__38395\,
            I => \N__38386\
        );

    \I__7391\ : Span4Mux_v
    port map (
            O => \N__38392\,
            I => \N__38383\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__38389\,
            I => \N__38378\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__38386\,
            I => \N__38378\
        );

    \I__7388\ : Span4Mux_h
    port map (
            O => \N__38383\,
            I => \N__38375\
        );

    \I__7387\ : Odrv4
    port map (
            O => \N__38378\,
            I => n306
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__38375\,
            I => n306
        );

    \I__7385\ : CascadeMux
    port map (
            O => \N__38370\,
            I => \n2031_cascade_\
        );

    \I__7384\ : InMux
    port map (
            O => \N__38367\,
            I => \N__38364\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__38364\,
            I => n11964
        );

    \I__7382\ : InMux
    port map (
            O => \N__38361\,
            I => \N__38354\
        );

    \I__7381\ : InMux
    port map (
            O => \N__38360\,
            I => \N__38354\
        );

    \I__7380\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38351\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__38354\,
            I => \N__38348\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__38351\,
            I => \N__38345\
        );

    \I__7377\ : Span4Mux_v
    port map (
            O => \N__38348\,
            I => \N__38342\
        );

    \I__7376\ : Sp12to4
    port map (
            O => \N__38345\,
            I => \N__38339\
        );

    \I__7375\ : Odrv4
    port map (
            O => \N__38342\,
            I => n305
        );

    \I__7374\ : Odrv12
    port map (
            O => \N__38339\,
            I => n305
        );

    \I__7373\ : InMux
    port map (
            O => \N__38334\,
            I => \N__38331\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__38331\,
            I => \N__38328\
        );

    \I__7371\ : Span4Mux_v
    port map (
            O => \N__38328\,
            I => \N__38325\
        );

    \I__7370\ : Odrv4
    port map (
            O => \N__38325\,
            I => n2001
        );

    \I__7369\ : CascadeMux
    port map (
            O => \N__38322\,
            I => \N__38318\
        );

    \I__7368\ : CascadeMux
    port map (
            O => \N__38321\,
            I => \N__38315\
        );

    \I__7367\ : InMux
    port map (
            O => \N__38318\,
            I => \N__38312\
        );

    \I__7366\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38309\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__38312\,
            I => \N__38306\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__38309\,
            I => \N__38303\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__38306\,
            I => \N__38297\
        );

    \I__7362\ : Span4Mux_v
    port map (
            O => \N__38303\,
            I => \N__38297\
        );

    \I__7361\ : InMux
    port map (
            O => \N__38302\,
            I => \N__38294\
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__38297\,
            I => n2033
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__38294\,
            I => n2033
        );

    \I__7358\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38286\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__38286\,
            I => \N__38283\
        );

    \I__7356\ : Odrv4
    port map (
            O => \N__38283\,
            I => n1996
        );

    \I__7355\ : CascadeMux
    port map (
            O => \N__38280\,
            I => \N__38276\
        );

    \I__7354\ : InMux
    port map (
            O => \N__38279\,
            I => \N__38273\
        );

    \I__7353\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38270\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__38273\,
            I => \N__38264\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__38270\,
            I => \N__38264\
        );

    \I__7350\ : CascadeMux
    port map (
            O => \N__38269\,
            I => \N__38261\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__38264\,
            I => \N__38258\
        );

    \I__7348\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38255\
        );

    \I__7347\ : Odrv4
    port map (
            O => \N__38258\,
            I => n2028
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__38255\,
            I => n2028
        );

    \I__7345\ : InMux
    port map (
            O => \N__38250\,
            I => \N__38247\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__38247\,
            I => \N__38244\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__38244\,
            I => \N__38241\
        );

    \I__7342\ : Odrv4
    port map (
            O => \N__38241\,
            I => n2000
        );

    \I__7341\ : CascadeMux
    port map (
            O => \N__38238\,
            I => \N__38235\
        );

    \I__7340\ : InMux
    port map (
            O => \N__38235\,
            I => \N__38228\
        );

    \I__7339\ : InMux
    port map (
            O => \N__38234\,
            I => \N__38228\
        );

    \I__7338\ : InMux
    port map (
            O => \N__38233\,
            I => \N__38225\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__38228\,
            I => \N__38222\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__38225\,
            I => n1933
        );

    \I__7335\ : Odrv4
    port map (
            O => \N__38222\,
            I => n1933
        );

    \I__7334\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38214\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__38214\,
            I => \N__38211\
        );

    \I__7332\ : Span4Mux_v
    port map (
            O => \N__38211\,
            I => \N__38202\
        );

    \I__7331\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38199\
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__38209\,
            I => \N__38192\
        );

    \I__7329\ : CascadeMux
    port map (
            O => \N__38208\,
            I => \N__38188\
        );

    \I__7328\ : CascadeMux
    port map (
            O => \N__38207\,
            I => \N__38185\
        );

    \I__7327\ : CascadeMux
    port map (
            O => \N__38206\,
            I => \N__38181\
        );

    \I__7326\ : CascadeMux
    port map (
            O => \N__38205\,
            I => \N__38175\
        );

    \I__7325\ : Span4Mux_v
    port map (
            O => \N__38202\,
            I => \N__38168\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__38199\,
            I => \N__38168\
        );

    \I__7323\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38161\
        );

    \I__7322\ : InMux
    port map (
            O => \N__38197\,
            I => \N__38161\
        );

    \I__7321\ : InMux
    port map (
            O => \N__38196\,
            I => \N__38161\
        );

    \I__7320\ : InMux
    port map (
            O => \N__38195\,
            I => \N__38148\
        );

    \I__7319\ : InMux
    port map (
            O => \N__38192\,
            I => \N__38148\
        );

    \I__7318\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38148\
        );

    \I__7317\ : InMux
    port map (
            O => \N__38188\,
            I => \N__38148\
        );

    \I__7316\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38148\
        );

    \I__7315\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38148\
        );

    \I__7314\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38143\
        );

    \I__7313\ : InMux
    port map (
            O => \N__38180\,
            I => \N__38143\
        );

    \I__7312\ : InMux
    port map (
            O => \N__38179\,
            I => \N__38134\
        );

    \I__7311\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38134\
        );

    \I__7310\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38134\
        );

    \I__7309\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38134\
        );

    \I__7308\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38131\
        );

    \I__7307\ : Odrv4
    port map (
            O => \N__38168\,
            I => n1950
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__38161\,
            I => n1950
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__38148\,
            I => n1950
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__38143\,
            I => n1950
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__38134\,
            I => n1950
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__38131\,
            I => n1950
        );

    \I__7301\ : CascadeMux
    port map (
            O => \N__38118\,
            I => \N__38114\
        );

    \I__7300\ : CascadeMux
    port map (
            O => \N__38117\,
            I => \N__38111\
        );

    \I__7299\ : InMux
    port map (
            O => \N__38114\,
            I => \N__38108\
        );

    \I__7298\ : InMux
    port map (
            O => \N__38111\,
            I => \N__38105\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__38108\,
            I => \N__38100\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__38105\,
            I => \N__38100\
        );

    \I__7295\ : Span4Mux_h
    port map (
            O => \N__38100\,
            I => \N__38096\
        );

    \I__7294\ : InMux
    port map (
            O => \N__38099\,
            I => \N__38093\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__38096\,
            I => n2032
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__38093\,
            I => n2032
        );

    \I__7291\ : CascadeMux
    port map (
            O => \N__38088\,
            I => \N__38085\
        );

    \I__7290\ : InMux
    port map (
            O => \N__38085\,
            I => \N__38082\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__38082\,
            I => n33_adj_654
        );

    \I__7288\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38076\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__38076\,
            I => \N__38073\
        );

    \I__7286\ : Span4Mux_h
    port map (
            O => \N__38073\,
            I => \N__38070\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__38070\,
            I => n33
        );

    \I__7284\ : InMux
    port map (
            O => \N__38067\,
            I => \bfn_10_21_0_\
        );

    \I__7283\ : CascadeMux
    port map (
            O => \N__38064\,
            I => \N__38061\
        );

    \I__7282\ : InMux
    port map (
            O => \N__38061\,
            I => \N__38058\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__38058\,
            I => n32_adj_653
        );

    \I__7280\ : InMux
    port map (
            O => \N__38055\,
            I => n12968
        );

    \I__7279\ : CascadeMux
    port map (
            O => \N__38052\,
            I => \N__38049\
        );

    \I__7278\ : InMux
    port map (
            O => \N__38049\,
            I => \N__38045\
        );

    \I__7277\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38042\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__38045\,
            I => n1922
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__38042\,
            I => n1922
        );

    \I__7274\ : InMux
    port map (
            O => \N__38037\,
            I => \N__38034\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__38034\,
            I => n1989
        );

    \I__7272\ : CascadeMux
    port map (
            O => \N__38031\,
            I => \n1922_cascade_\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__38028\,
            I => \N__38025\
        );

    \I__7270\ : InMux
    port map (
            O => \N__38025\,
            I => \N__38021\
        );

    \I__7269\ : InMux
    port map (
            O => \N__38024\,
            I => \N__38018\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__38021\,
            I => \N__38015\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__38018\,
            I => \N__38012\
        );

    \I__7266\ : Span4Mux_h
    port map (
            O => \N__38015\,
            I => \N__38006\
        );

    \I__7265\ : Span4Mux_v
    port map (
            O => \N__38012\,
            I => \N__38006\
        );

    \I__7264\ : InMux
    port map (
            O => \N__38011\,
            I => \N__38003\
        );

    \I__7263\ : Odrv4
    port map (
            O => \N__38006\,
            I => n2021
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__38003\,
            I => n2021
        );

    \I__7261\ : InMux
    port map (
            O => \N__37998\,
            I => \N__37995\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__37995\,
            I => n14416
        );

    \I__7259\ : CascadeMux
    port map (
            O => \N__37992\,
            I => \n14420_cascade_\
        );

    \I__7258\ : CascadeMux
    port map (
            O => \N__37989\,
            I => \n1950_cascade_\
        );

    \I__7257\ : InMux
    port map (
            O => \N__37986\,
            I => \N__37983\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37980\
        );

    \I__7255\ : Span4Mux_v
    port map (
            O => \N__37980\,
            I => \N__37977\
        );

    \I__7254\ : Odrv4
    port map (
            O => \N__37977\,
            I => n1998
        );

    \I__7253\ : CascadeMux
    port map (
            O => \N__37974\,
            I => \N__37970\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__37973\,
            I => \N__37967\
        );

    \I__7251\ : InMux
    port map (
            O => \N__37970\,
            I => \N__37963\
        );

    \I__7250\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37960\
        );

    \I__7249\ : InMux
    port map (
            O => \N__37966\,
            I => \N__37957\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__37963\,
            I => \N__37952\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__37960\,
            I => \N__37952\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__37957\,
            I => \N__37947\
        );

    \I__7245\ : Span4Mux_h
    port map (
            O => \N__37952\,
            I => \N__37947\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__37947\,
            I => n2030
        );

    \I__7243\ : InMux
    port map (
            O => \N__37944\,
            I => \N__37941\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__37941\,
            I => \N__37938\
        );

    \I__7241\ : Span12Mux_s9_h
    port map (
            O => \N__37938\,
            I => \N__37934\
        );

    \I__7240\ : InMux
    port map (
            O => \N__37937\,
            I => \N__37931\
        );

    \I__7239\ : Odrv12
    port map (
            O => \N__37934\,
            I => n15666
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__37931\,
            I => n15666
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__37926\,
            I => \N__37923\
        );

    \I__7236\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37919\
        );

    \I__7235\ : InMux
    port map (
            O => \N__37922\,
            I => \N__37916\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__37919\,
            I => n1917
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__37916\,
            I => n1917
        );

    \I__7232\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37908\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__37908\,
            I => n1988
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__37905\,
            I => \N__37901\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__37904\,
            I => \N__37898\
        );

    \I__7228\ : InMux
    port map (
            O => \N__37901\,
            I => \N__37895\
        );

    \I__7227\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37892\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__37895\,
            I => n1921
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__37892\,
            I => n1921
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__37887\,
            I => \N__37883\
        );

    \I__7223\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37880\
        );

    \I__7222\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37877\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__37880\,
            I => \N__37874\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__37877\,
            I => \N__37871\
        );

    \I__7219\ : Span4Mux_h
    port map (
            O => \N__37874\,
            I => \N__37867\
        );

    \I__7218\ : Span4Mux_h
    port map (
            O => \N__37871\,
            I => \N__37864\
        );

    \I__7217\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37861\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__37867\,
            I => n2020
        );

    \I__7215\ : Odrv4
    port map (
            O => \N__37864\,
            I => n2020
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__37861\,
            I => n2020
        );

    \I__7213\ : InMux
    port map (
            O => \N__37854\,
            I => \N__37851\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__37851\,
            I => n11966
        );

    \I__7211\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37844\
        );

    \I__7210\ : InMux
    port map (
            O => \N__37847\,
            I => \N__37841\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__37844\,
            I => \N__37837\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__37841\,
            I => \N__37834\
        );

    \I__7207\ : InMux
    port map (
            O => \N__37840\,
            I => \N__37831\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__37837\,
            I => \N__37828\
        );

    \I__7205\ : Span4Mux_v
    port map (
            O => \N__37834\,
            I => \N__37825\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__37831\,
            I => encoder0_position_9
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__37828\,
            I => encoder0_position_9
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__37825\,
            I => encoder0_position_9
        );

    \I__7201\ : InMux
    port map (
            O => \N__37818\,
            I => \N__37813\
        );

    \I__7200\ : InMux
    port map (
            O => \N__37817\,
            I => \N__37810\
        );

    \I__7199\ : InMux
    port map (
            O => \N__37816\,
            I => \N__37807\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__37813\,
            I => \N__37800\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__37810\,
            I => \N__37800\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__37807\,
            I => \N__37800\
        );

    \I__7195\ : Odrv12
    port map (
            O => \N__37800\,
            I => n310
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__37797\,
            I => \N__37794\
        );

    \I__7193\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37791\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__37791\,
            I => \N__37788\
        );

    \I__7191\ : Span4Mux_h
    port map (
            O => \N__37788\,
            I => \N__37783\
        );

    \I__7190\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37780\
        );

    \I__7189\ : InMux
    port map (
            O => \N__37786\,
            I => \N__37777\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__37783\,
            I => n1927
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__37780\,
            I => n1927
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__37777\,
            I => n1927
        );

    \I__7185\ : InMux
    port map (
            O => \N__37770\,
            I => \N__37766\
        );

    \I__7184\ : CascadeMux
    port map (
            O => \N__37769\,
            I => \N__37763\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__37766\,
            I => \N__37760\
        );

    \I__7182\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37757\
        );

    \I__7181\ : Odrv4
    port map (
            O => \N__37760\,
            I => n1923
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__37757\,
            I => n1923
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__37752\,
            I => \N__37749\
        );

    \I__7178\ : InMux
    port map (
            O => \N__37749\,
            I => \N__37745\
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__37748\,
            I => \N__37742\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37738\
        );

    \I__7175\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37735\
        );

    \I__7174\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37732\
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__37738\,
            I => n1926
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__37735\,
            I => n1926
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__37732\,
            I => n1926
        );

    \I__7170\ : CascadeMux
    port map (
            O => \N__37725\,
            I => \n1923_cascade_\
        );

    \I__7169\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37718\
        );

    \I__7168\ : CascadeMux
    port map (
            O => \N__37721\,
            I => \N__37715\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__37718\,
            I => \N__37711\
        );

    \I__7166\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37708\
        );

    \I__7165\ : InMux
    port map (
            O => \N__37714\,
            I => \N__37705\
        );

    \I__7164\ : Odrv4
    port map (
            O => \N__37711\,
            I => n1924
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__37708\,
            I => n1924
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__37705\,
            I => n1924
        );

    \I__7161\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37695\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__37695\,
            I => n14408
        );

    \I__7159\ : CascadeMux
    port map (
            O => \N__37692\,
            I => \n1921_cascade_\
        );

    \I__7158\ : InMux
    port map (
            O => \N__37689\,
            I => \N__37686\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__37686\,
            I => n14410
        );

    \I__7156\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37680\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__37680\,
            I => n1995
        );

    \I__7154\ : CascadeMux
    port map (
            O => \N__37677\,
            I => \N__37673\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__37676\,
            I => \N__37670\
        );

    \I__7152\ : InMux
    port map (
            O => \N__37673\,
            I => \N__37667\
        );

    \I__7151\ : InMux
    port map (
            O => \N__37670\,
            I => \N__37664\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__37667\,
            I => \N__37660\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37657\
        );

    \I__7148\ : InMux
    port map (
            O => \N__37663\,
            I => \N__37654\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__37660\,
            I => \N__37651\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__37657\,
            I => \N__37646\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__37654\,
            I => \N__37646\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__37651\,
            I => n2027
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__37646\,
            I => n2027
        );

    \I__7142\ : CascadeMux
    port map (
            O => \N__37641\,
            I => \N__37636\
        );

    \I__7141\ : CascadeMux
    port map (
            O => \N__37640\,
            I => \N__37633\
        );

    \I__7140\ : InMux
    port map (
            O => \N__37639\,
            I => \N__37630\
        );

    \I__7139\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37627\
        );

    \I__7138\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37624\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__37630\,
            I => n1925
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__37627\,
            I => n1925
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__37624\,
            I => n1925
        );

    \I__7134\ : InMux
    port map (
            O => \N__37617\,
            I => \N__37614\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__37614\,
            I => \N__37611\
        );

    \I__7132\ : Odrv12
    port map (
            O => \N__37611\,
            I => n6_adj_586
        );

    \I__7131\ : InMux
    port map (
            O => \N__37608\,
            I => n12430
        );

    \I__7130\ : InMux
    port map (
            O => \N__37605\,
            I => n12431
        );

    \I__7129\ : InMux
    port map (
            O => \N__37602\,
            I => n12432
        );

    \I__7128\ : InMux
    port map (
            O => \N__37599\,
            I => n12433
        );

    \I__7127\ : InMux
    port map (
            O => \N__37596\,
            I => n12434
        );

    \I__7126\ : InMux
    port map (
            O => \N__37593\,
            I => n12421
        );

    \I__7125\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37587\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__37587\,
            I => \N__37584\
        );

    \I__7123\ : Odrv4
    port map (
            O => \N__37584\,
            I => n14_adj_594
        );

    \I__7122\ : InMux
    port map (
            O => \N__37581\,
            I => n12422
        );

    \I__7121\ : InMux
    port map (
            O => \N__37578\,
            I => \N__37575\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__37575\,
            I => \N__37572\
        );

    \I__7119\ : Odrv4
    port map (
            O => \N__37572\,
            I => n13_adj_593
        );

    \I__7118\ : InMux
    port map (
            O => \N__37569\,
            I => n12423
        );

    \I__7117\ : InMux
    port map (
            O => \N__37566\,
            I => n12424
        );

    \I__7116\ : InMux
    port map (
            O => \N__37563\,
            I => n12425
        );

    \I__7115\ : InMux
    port map (
            O => \N__37560\,
            I => \N__37557\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__37557\,
            I => \N__37554\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__37554\,
            I => n10_adj_590
        );

    \I__7112\ : InMux
    port map (
            O => \N__37551\,
            I => n12426
        );

    \I__7111\ : InMux
    port map (
            O => \N__37548\,
            I => \bfn_9_32_0_\
        );

    \I__7110\ : InMux
    port map (
            O => \N__37545\,
            I => n12428
        );

    \I__7109\ : InMux
    port map (
            O => \N__37542\,
            I => n12429
        );

    \I__7108\ : InMux
    port map (
            O => \N__37539\,
            I => \N__37536\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__37536\,
            I => \N__37533\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__37533\,
            I => n24_adj_604
        );

    \I__7105\ : InMux
    port map (
            O => \N__37530\,
            I => \N__37527\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__37527\,
            I => \N__37524\
        );

    \I__7103\ : Odrv12
    port map (
            O => \N__37524\,
            I => \pwm_setpoint_23_N_171_1\
        );

    \I__7102\ : InMux
    port map (
            O => \N__37521\,
            I => n12412
        );

    \I__7101\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37515\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__37515\,
            I => \N__37512\
        );

    \I__7099\ : Odrv4
    port map (
            O => \N__37512\,
            I => n23_adj_603
        );

    \I__7098\ : InMux
    port map (
            O => \N__37509\,
            I => n12413
        );

    \I__7097\ : InMux
    port map (
            O => \N__37506\,
            I => \N__37503\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__37503\,
            I => n22_adj_602
        );

    \I__7095\ : InMux
    port map (
            O => \N__37500\,
            I => n12414
        );

    \I__7094\ : InMux
    port map (
            O => \N__37497\,
            I => n12415
        );

    \I__7093\ : InMux
    port map (
            O => \N__37494\,
            I => n12416
        );

    \I__7092\ : InMux
    port map (
            O => \N__37491\,
            I => n12417
        );

    \I__7091\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37485\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__37485\,
            I => \N__37482\
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__37482\,
            I => n18_adj_598
        );

    \I__7088\ : InMux
    port map (
            O => \N__37479\,
            I => n12418
        );

    \I__7087\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37473\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37470\
        );

    \I__7085\ : Odrv4
    port map (
            O => \N__37470\,
            I => n17_adj_597
        );

    \I__7084\ : InMux
    port map (
            O => \N__37467\,
            I => \bfn_9_31_0_\
        );

    \I__7083\ : InMux
    port map (
            O => \N__37464\,
            I => n12420
        );

    \I__7082\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37458\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__37458\,
            I => \N__37455\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__37455\,
            I => \N__37452\
        );

    \I__7079\ : Odrv4
    port map (
            O => \N__37452\,
            I => encoder0_position_scaled_19
        );

    \I__7078\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37446\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__37446\,
            I => \N__37443\
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__37443\,
            I => n25_adj_605
        );

    \I__7075\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37437\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__37437\,
            I => \N__37434\
        );

    \I__7073\ : Odrv12
    port map (
            O => \N__37434\,
            I => \pwm_setpoint_23_N_171_0\
        );

    \I__7072\ : InMux
    port map (
            O => \N__37431\,
            I => \bfn_9_30_0_\
        );

    \I__7071\ : CascadeMux
    port map (
            O => \N__37428\,
            I => \quad_counter0.a_prev_N_543_cascade_\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__37425\,
            I => \N__37408\
        );

    \I__7069\ : CascadeMux
    port map (
            O => \N__37424\,
            I => \N__37404\
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__37423\,
            I => \N__37400\
        );

    \I__7067\ : CascadeMux
    port map (
            O => \N__37422\,
            I => \N__37396\
        );

    \I__7066\ : CascadeMux
    port map (
            O => \N__37421\,
            I => \N__37393\
        );

    \I__7065\ : CascadeMux
    port map (
            O => \N__37420\,
            I => \N__37389\
        );

    \I__7064\ : CascadeMux
    port map (
            O => \N__37419\,
            I => \N__37385\
        );

    \I__7063\ : CascadeMux
    port map (
            O => \N__37418\,
            I => \N__37381\
        );

    \I__7062\ : CascadeMux
    port map (
            O => \N__37417\,
            I => \N__37376\
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__37416\,
            I => \N__37372\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__37415\,
            I => \N__37368\
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__37414\,
            I => \N__37362\
        );

    \I__7058\ : CascadeMux
    port map (
            O => \N__37413\,
            I => \N__37358\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__37412\,
            I => \N__37354\
        );

    \I__7056\ : InMux
    port map (
            O => \N__37411\,
            I => \N__37336\
        );

    \I__7055\ : InMux
    port map (
            O => \N__37408\,
            I => \N__37336\
        );

    \I__7054\ : InMux
    port map (
            O => \N__37407\,
            I => \N__37336\
        );

    \I__7053\ : InMux
    port map (
            O => \N__37404\,
            I => \N__37336\
        );

    \I__7052\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37336\
        );

    \I__7051\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37336\
        );

    \I__7050\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37336\
        );

    \I__7049\ : InMux
    port map (
            O => \N__37396\,
            I => \N__37336\
        );

    \I__7048\ : InMux
    port map (
            O => \N__37393\,
            I => \N__37319\
        );

    \I__7047\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37319\
        );

    \I__7046\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37319\
        );

    \I__7045\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37319\
        );

    \I__7044\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37319\
        );

    \I__7043\ : InMux
    port map (
            O => \N__37384\,
            I => \N__37319\
        );

    \I__7042\ : InMux
    port map (
            O => \N__37381\,
            I => \N__37319\
        );

    \I__7041\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37319\
        );

    \I__7040\ : InMux
    port map (
            O => \N__37379\,
            I => \N__37304\
        );

    \I__7039\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37304\
        );

    \I__7038\ : InMux
    port map (
            O => \N__37375\,
            I => \N__37304\
        );

    \I__7037\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37304\
        );

    \I__7036\ : InMux
    port map (
            O => \N__37371\,
            I => \N__37304\
        );

    \I__7035\ : InMux
    port map (
            O => \N__37368\,
            I => \N__37304\
        );

    \I__7034\ : InMux
    port map (
            O => \N__37367\,
            I => \N__37304\
        );

    \I__7033\ : InMux
    port map (
            O => \N__37366\,
            I => \N__37287\
        );

    \I__7032\ : InMux
    port map (
            O => \N__37365\,
            I => \N__37287\
        );

    \I__7031\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37287\
        );

    \I__7030\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37287\
        );

    \I__7029\ : InMux
    port map (
            O => \N__37358\,
            I => \N__37287\
        );

    \I__7028\ : InMux
    port map (
            O => \N__37357\,
            I => \N__37287\
        );

    \I__7027\ : InMux
    port map (
            O => \N__37354\,
            I => \N__37287\
        );

    \I__7026\ : InMux
    port map (
            O => \N__37353\,
            I => \N__37287\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__37336\,
            I => \N__37280\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37280\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__37304\,
            I => \N__37280\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__37287\,
            I => \N__37277\
        );

    \I__7021\ : Span4Mux_v
    port map (
            O => \N__37280\,
            I => \N__37274\
        );

    \I__7020\ : Odrv4
    port map (
            O => \N__37277\,
            I => \quad_counter0.direction_N_536\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__37274\,
            I => \quad_counter0.direction_N_536\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__37269\,
            I => \N__37266\
        );

    \I__7017\ : InMux
    port map (
            O => \N__37266\,
            I => \N__37262\
        );

    \I__7016\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37259\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__37262\,
            I => \N__37256\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__37259\,
            I => \N__37252\
        );

    \I__7013\ : Span4Mux_h
    port map (
            O => \N__37256\,
            I => \N__37249\
        );

    \I__7012\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37246\
        );

    \I__7011\ : Odrv12
    port map (
            O => \N__37252\,
            I => n3024
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__37249\,
            I => n3024
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__37246\,
            I => n3024
        );

    \I__7008\ : CascadeMux
    port map (
            O => \N__37239\,
            I => \N__37236\
        );

    \I__7007\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37233\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__37233\,
            I => \N__37230\
        );

    \I__7005\ : Span12Mux_h
    port map (
            O => \N__37230\,
            I => \N__37227\
        );

    \I__7004\ : Odrv12
    port map (
            O => \N__37227\,
            I => n3091
        );

    \I__7003\ : CascadeMux
    port map (
            O => \N__37224\,
            I => \N__37220\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__37223\,
            I => \N__37212\
        );

    \I__7001\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37207\
        );

    \I__7000\ : InMux
    port map (
            O => \N__37219\,
            I => \N__37200\
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__37218\,
            I => \N__37197\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__37217\,
            I => \N__37190\
        );

    \I__6997\ : InMux
    port map (
            O => \N__37216\,
            I => \N__37187\
        );

    \I__6996\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37184\
        );

    \I__6995\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37179\
        );

    \I__6994\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37179\
        );

    \I__6993\ : InMux
    port map (
            O => \N__37210\,
            I => \N__37176\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__37207\,
            I => \N__37173\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__37206\,
            I => \N__37166\
        );

    \I__6990\ : CascadeMux
    port map (
            O => \N__37205\,
            I => \N__37163\
        );

    \I__6989\ : CascadeMux
    port map (
            O => \N__37204\,
            I => \N__37159\
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__37203\,
            I => \N__37150\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__37200\,
            I => \N__37146\
        );

    \I__6986\ : InMux
    port map (
            O => \N__37197\,
            I => \N__37141\
        );

    \I__6985\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37141\
        );

    \I__6984\ : InMux
    port map (
            O => \N__37195\,
            I => \N__37132\
        );

    \I__6983\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37132\
        );

    \I__6982\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37132\
        );

    \I__6981\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37132\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__37187\,
            I => \N__37127\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__37184\,
            I => \N__37127\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__37179\,
            I => \N__37124\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__37176\,
            I => \N__37121\
        );

    \I__6976\ : Span12Mux_v
    port map (
            O => \N__37173\,
            I => \N__37118\
        );

    \I__6975\ : InMux
    port map (
            O => \N__37172\,
            I => \N__37113\
        );

    \I__6974\ : InMux
    port map (
            O => \N__37171\,
            I => \N__37113\
        );

    \I__6973\ : InMux
    port map (
            O => \N__37170\,
            I => \N__37110\
        );

    \I__6972\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37101\
        );

    \I__6971\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37101\
        );

    \I__6970\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37101\
        );

    \I__6969\ : InMux
    port map (
            O => \N__37162\,
            I => \N__37101\
        );

    \I__6968\ : InMux
    port map (
            O => \N__37159\,
            I => \N__37096\
        );

    \I__6967\ : InMux
    port map (
            O => \N__37158\,
            I => \N__37096\
        );

    \I__6966\ : InMux
    port map (
            O => \N__37157\,
            I => \N__37093\
        );

    \I__6965\ : InMux
    port map (
            O => \N__37156\,
            I => \N__37088\
        );

    \I__6964\ : InMux
    port map (
            O => \N__37155\,
            I => \N__37088\
        );

    \I__6963\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37079\
        );

    \I__6962\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37079\
        );

    \I__6961\ : InMux
    port map (
            O => \N__37150\,
            I => \N__37079\
        );

    \I__6960\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37079\
        );

    \I__6959\ : Span4Mux_h
    port map (
            O => \N__37146\,
            I => \N__37070\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__37141\,
            I => \N__37070\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__37132\,
            I => \N__37070\
        );

    \I__6956\ : Span4Mux_h
    port map (
            O => \N__37127\,
            I => \N__37070\
        );

    \I__6955\ : Span4Mux_h
    port map (
            O => \N__37124\,
            I => \N__37065\
        );

    \I__6954\ : Span4Mux_v
    port map (
            O => \N__37121\,
            I => \N__37065\
        );

    \I__6953\ : Odrv12
    port map (
            O => \N__37118\,
            I => n3039
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__37113\,
            I => n3039
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__37110\,
            I => n3039
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__37101\,
            I => n3039
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__37096\,
            I => n3039
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__37093\,
            I => n3039
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__37088\,
            I => n3039
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__37079\,
            I => n3039
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__37070\,
            I => n3039
        );

    \I__6944\ : Odrv4
    port map (
            O => \N__37065\,
            I => n3039
        );

    \I__6943\ : CascadeMux
    port map (
            O => \N__37044\,
            I => \N__37040\
        );

    \I__6942\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37036\
        );

    \I__6941\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37033\
        );

    \I__6940\ : InMux
    port map (
            O => \N__37039\,
            I => \N__37030\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__37036\,
            I => \N__37025\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__37033\,
            I => \N__37025\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__37030\,
            I => \N__37022\
        );

    \I__6936\ : Span4Mux_h
    port map (
            O => \N__37025\,
            I => \N__37019\
        );

    \I__6935\ : Span12Mux_s4_v
    port map (
            O => \N__37022\,
            I => \N__37016\
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__37019\,
            I => n3123
        );

    \I__6933\ : Odrv12
    port map (
            O => \N__37016\,
            I => n3123
        );

    \I__6932\ : InMux
    port map (
            O => \N__37011\,
            I => \N__37008\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__37008\,
            I => \N__37005\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__37005\,
            I => \N__37002\
        );

    \I__6929\ : IoSpan4Mux
    port map (
            O => \N__37002\,
            I => \N__36999\
        );

    \I__6928\ : IoSpan4Mux
    port map (
            O => \N__36999\,
            I => \N__36996\
        );

    \I__6927\ : Odrv4
    port map (
            O => \N__36996\,
            I => \ENCODER0_A_N\
        );

    \I__6926\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36984\
        );

    \I__6925\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36984\
        );

    \I__6924\ : InMux
    port map (
            O => \N__36991\,
            I => \N__36984\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__36984\,
            I => \quad_counter0.a_new_0\
        );

    \I__6922\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36978\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__36978\,
            I => \N__36975\
        );

    \I__6920\ : Span4Mux_v
    port map (
            O => \N__36975\,
            I => \N__36972\
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__36972\,
            I => encoder0_position_scaled_21
        );

    \I__6918\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36966\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__36966\,
            I => \N__36963\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__36963\,
            I => \N__36960\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__36960\,
            I => encoder0_position_scaled_4
        );

    \I__6914\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36954\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__36954\,
            I => \N__36951\
        );

    \I__6912\ : Span4Mux_h
    port map (
            O => \N__36951\,
            I => \N__36948\
        );

    \I__6911\ : Odrv4
    port map (
            O => \N__36948\,
            I => encoder0_position_scaled_5
        );

    \I__6910\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36942\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__36942\,
            I => \N__36939\
        );

    \I__6908\ : Span4Mux_h
    port map (
            O => \N__36939\,
            I => \N__36936\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__36936\,
            I => encoder0_position_scaled_22
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__36933\,
            I => \N__36929\
        );

    \I__6905\ : CascadeMux
    port map (
            O => \N__36932\,
            I => \N__36926\
        );

    \I__6904\ : InMux
    port map (
            O => \N__36929\,
            I => \N__36923\
        );

    \I__6903\ : InMux
    port map (
            O => \N__36926\,
            I => \N__36920\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__36923\,
            I => \N__36917\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__36920\,
            I => \N__36914\
        );

    \I__6900\ : Span4Mux_v
    port map (
            O => \N__36917\,
            I => \N__36909\
        );

    \I__6899\ : Span4Mux_h
    port map (
            O => \N__36914\,
            I => \N__36909\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__36909\,
            I => n3133
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__36906\,
            I => \N__36902\
        );

    \I__6896\ : InMux
    port map (
            O => \N__36905\,
            I => \N__36899\
        );

    \I__6895\ : InMux
    port map (
            O => \N__36902\,
            I => \N__36895\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__36899\,
            I => \N__36892\
        );

    \I__6893\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36889\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__36895\,
            I => \N__36886\
        );

    \I__6891\ : Span4Mux_h
    port map (
            O => \N__36892\,
            I => \N__36883\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__36889\,
            I => n3132
        );

    \I__6889\ : Odrv12
    port map (
            O => \N__36886\,
            I => n3132
        );

    \I__6888\ : Odrv4
    port map (
            O => \N__36883\,
            I => n3132
        );

    \I__6887\ : CascadeMux
    port map (
            O => \N__36876\,
            I => \N__36871\
        );

    \I__6886\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36868\
        );

    \I__6885\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36865\
        );

    \I__6884\ : InMux
    port map (
            O => \N__36871\,
            I => \N__36862\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36859\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36856\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36853\
        );

    \I__6880\ : Span4Mux_v
    port map (
            O => \N__36859\,
            I => \N__36850\
        );

    \I__6879\ : Span4Mux_h
    port map (
            O => \N__36856\,
            I => \N__36845\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__36853\,
            I => \N__36845\
        );

    \I__6877\ : Span4Mux_h
    port map (
            O => \N__36850\,
            I => \N__36842\
        );

    \I__6876\ : Odrv4
    port map (
            O => \N__36845\,
            I => n3129
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__36842\,
            I => n3129
        );

    \I__6874\ : InMux
    port map (
            O => \N__36837\,
            I => \N__36832\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__36836\,
            I => \N__36829\
        );

    \I__6872\ : InMux
    port map (
            O => \N__36835\,
            I => \N__36826\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__36832\,
            I => \N__36823\
        );

    \I__6870\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36820\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__36826\,
            I => \N__36817\
        );

    \I__6868\ : Span4Mux_h
    port map (
            O => \N__36823\,
            I => \N__36814\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__36820\,
            I => \N__36811\
        );

    \I__6866\ : Span4Mux_v
    port map (
            O => \N__36817\,
            I => \N__36808\
        );

    \I__6865\ : Odrv4
    port map (
            O => \N__36814\,
            I => n3130
        );

    \I__6864\ : Odrv12
    port map (
            O => \N__36811\,
            I => n3130
        );

    \I__6863\ : Odrv4
    port map (
            O => \N__36808\,
            I => n3130
        );

    \I__6862\ : CascadeMux
    port map (
            O => \N__36801\,
            I => \n11930_cascade_\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__36798\,
            I => \N__36795\
        );

    \I__6860\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36791\
        );

    \I__6859\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36788\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__36791\,
            I => \N__36784\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__36788\,
            I => \N__36781\
        );

    \I__6856\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36778\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__36784\,
            I => \N__36773\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__36781\,
            I => \N__36773\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__36778\,
            I => n3131
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__36773\,
            I => n3131
        );

    \I__6851\ : CascadeMux
    port map (
            O => \N__36768\,
            I => \N__36765\
        );

    \I__6850\ : InMux
    port map (
            O => \N__36765\,
            I => \N__36762\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__36762\,
            I => \N__36759\
        );

    \I__6848\ : Span4Mux_h
    port map (
            O => \N__36759\,
            I => \N__36756\
        );

    \I__6847\ : Odrv4
    port map (
            O => \N__36756\,
            I => n13819
        );

    \I__6846\ : InMux
    port map (
            O => \N__36753\,
            I => \quad_counter0.n13049\
        );

    \I__6845\ : InMux
    port map (
            O => \N__36750\,
            I => \quad_counter0.n13050\
        );

    \I__6844\ : InMux
    port map (
            O => \N__36747\,
            I => \quad_counter0.n13051\
        );

    \I__6843\ : InMux
    port map (
            O => \N__36744\,
            I => \quad_counter0.n13052\
        );

    \I__6842\ : InMux
    port map (
            O => \N__36741\,
            I => \quad_counter0.n13053\
        );

    \I__6841\ : InMux
    port map (
            O => \N__36738\,
            I => \quad_counter0.n13054\
        );

    \I__6840\ : InMux
    port map (
            O => \N__36735\,
            I => \quad_counter0.n13055\
        );

    \I__6839\ : InMux
    port map (
            O => \N__36732\,
            I => \N__36729\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__36729\,
            I => \N__36726\
        );

    \I__6837\ : Span4Mux_v
    port map (
            O => \N__36726\,
            I => \N__36723\
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__36723\,
            I => encoder0_position_scaled_17
        );

    \I__6835\ : CascadeMux
    port map (
            O => \N__36720\,
            I => \N__36715\
        );

    \I__6834\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36712\
        );

    \I__6833\ : InMux
    port map (
            O => \N__36718\,
            I => \N__36709\
        );

    \I__6832\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36706\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__36712\,
            I => \N__36703\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__36709\,
            I => \N__36700\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__36706\,
            I => encoder0_position_14
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__36703\,
            I => encoder0_position_14
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__36700\,
            I => encoder0_position_14
        );

    \I__6826\ : InMux
    port map (
            O => \N__36693\,
            I => \bfn_9_24_0_\
        );

    \I__6825\ : InMux
    port map (
            O => \N__36690\,
            I => \quad_counter0.n13041\
        );

    \I__6824\ : InMux
    port map (
            O => \N__36687\,
            I => \quad_counter0.n13042\
        );

    \I__6823\ : InMux
    port map (
            O => \N__36684\,
            I => \quad_counter0.n13043\
        );

    \I__6822\ : InMux
    port map (
            O => \N__36681\,
            I => \quad_counter0.n13044\
        );

    \I__6821\ : InMux
    port map (
            O => \N__36678\,
            I => \quad_counter0.n13045\
        );

    \I__6820\ : InMux
    port map (
            O => \N__36675\,
            I => \quad_counter0.n13046\
        );

    \I__6819\ : InMux
    port map (
            O => \N__36672\,
            I => \quad_counter0.n13047\
        );

    \I__6818\ : InMux
    port map (
            O => \N__36669\,
            I => \bfn_9_25_0_\
        );

    \I__6817\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36659\
        );

    \I__6816\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36659\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__36664\,
            I => \N__36656\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__36659\,
            I => \N__36653\
        );

    \I__6813\ : InMux
    port map (
            O => \N__36656\,
            I => \N__36650\
        );

    \I__6812\ : Span4Mux_h
    port map (
            O => \N__36653\,
            I => \N__36647\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__36650\,
            I => encoder0_position_8
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__36647\,
            I => encoder0_position_8
        );

    \I__6809\ : InMux
    port map (
            O => \N__36642\,
            I => \bfn_9_23_0_\
        );

    \I__6808\ : InMux
    port map (
            O => \N__36639\,
            I => \quad_counter0.n13033\
        );

    \I__6807\ : InMux
    port map (
            O => \N__36636\,
            I => \quad_counter0.n13034\
        );

    \I__6806\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36627\
        );

    \I__6805\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36627\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__36627\,
            I => \N__36623\
        );

    \I__6803\ : InMux
    port map (
            O => \N__36626\,
            I => \N__36620\
        );

    \I__6802\ : Span4Mux_h
    port map (
            O => \N__36623\,
            I => \N__36617\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__36620\,
            I => encoder0_position_11
        );

    \I__6800\ : Odrv4
    port map (
            O => \N__36617\,
            I => encoder0_position_11
        );

    \I__6799\ : InMux
    port map (
            O => \N__36612\,
            I => \quad_counter0.n13035\
        );

    \I__6798\ : InMux
    port map (
            O => \N__36609\,
            I => \N__36605\
        );

    \I__6797\ : InMux
    port map (
            O => \N__36608\,
            I => \N__36602\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36598\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__36602\,
            I => \N__36595\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__36601\,
            I => \N__36592\
        );

    \I__6793\ : Span4Mux_v
    port map (
            O => \N__36598\,
            I => \N__36589\
        );

    \I__6792\ : Span4Mux_h
    port map (
            O => \N__36595\,
            I => \N__36586\
        );

    \I__6791\ : InMux
    port map (
            O => \N__36592\,
            I => \N__36583\
        );

    \I__6790\ : Span4Mux_h
    port map (
            O => \N__36589\,
            I => \N__36578\
        );

    \I__6789\ : Span4Mux_v
    port map (
            O => \N__36586\,
            I => \N__36578\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__36583\,
            I => encoder0_position_12
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__36578\,
            I => encoder0_position_12
        );

    \I__6786\ : InMux
    port map (
            O => \N__36573\,
            I => \quad_counter0.n13036\
        );

    \I__6785\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36566\
        );

    \I__6784\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36562\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__36566\,
            I => \N__36559\
        );

    \I__6782\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36556\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__36562\,
            I => \N__36551\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__36559\,
            I => \N__36551\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__36556\,
            I => encoder0_position_13
        );

    \I__6778\ : Odrv4
    port map (
            O => \N__36551\,
            I => encoder0_position_13
        );

    \I__6777\ : InMux
    port map (
            O => \N__36546\,
            I => \quad_counter0.n13037\
        );

    \I__6776\ : InMux
    port map (
            O => \N__36543\,
            I => \quad_counter0.n13038\
        );

    \I__6775\ : InMux
    port map (
            O => \N__36540\,
            I => \quad_counter0.n13039\
        );

    \I__6774\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36533\
        );

    \I__6773\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36529\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__36533\,
            I => \N__36526\
        );

    \I__6771\ : InMux
    port map (
            O => \N__36532\,
            I => \N__36523\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__36529\,
            I => encoder0_position_0
        );

    \I__6769\ : Odrv4
    port map (
            O => \N__36526\,
            I => encoder0_position_0
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__36523\,
            I => encoder0_position_0
        );

    \I__6767\ : InMux
    port map (
            O => \N__36516\,
            I => \bfn_9_22_0_\
        );

    \I__6766\ : InMux
    port map (
            O => \N__36513\,
            I => \quad_counter0.n13025\
        );

    \I__6765\ : InMux
    port map (
            O => \N__36510\,
            I => \quad_counter0.n13026\
        );

    \I__6764\ : InMux
    port map (
            O => \N__36507\,
            I => \quad_counter0.n13027\
        );

    \I__6763\ : InMux
    port map (
            O => \N__36504\,
            I => \N__36500\
        );

    \I__6762\ : InMux
    port map (
            O => \N__36503\,
            I => \N__36496\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__36500\,
            I => \N__36493\
        );

    \I__6760\ : InMux
    port map (
            O => \N__36499\,
            I => \N__36490\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__36496\,
            I => encoder0_position_4
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__36493\,
            I => encoder0_position_4
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__36490\,
            I => encoder0_position_4
        );

    \I__6756\ : InMux
    port map (
            O => \N__36483\,
            I => \quad_counter0.n13028\
        );

    \I__6755\ : InMux
    port map (
            O => \N__36480\,
            I => \quad_counter0.n13029\
        );

    \I__6754\ : InMux
    port map (
            O => \N__36477\,
            I => \quad_counter0.n13030\
        );

    \I__6753\ : InMux
    port map (
            O => \N__36474\,
            I => \quad_counter0.n13031\
        );

    \I__6752\ : CascadeMux
    port map (
            O => \N__36471\,
            I => \n14558_cascade_\
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__36468\,
            I => \N__36465\
        );

    \I__6750\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36461\
        );

    \I__6749\ : InMux
    port map (
            O => \N__36464\,
            I => \N__36458\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__36461\,
            I => \N__36455\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__36458\,
            I => \N__36452\
        );

    \I__6746\ : Span4Mux_h
    port map (
            O => \N__36455\,
            I => \N__36448\
        );

    \I__6745\ : Span4Mux_h
    port map (
            O => \N__36452\,
            I => \N__36445\
        );

    \I__6744\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36442\
        );

    \I__6743\ : Odrv4
    port map (
            O => \N__36448\,
            I => n2019
        );

    \I__6742\ : Odrv4
    port map (
            O => \N__36445\,
            I => n2019
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__36442\,
            I => n2019
        );

    \I__6740\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__36432\,
            I => \N__36429\
        );

    \I__6738\ : Span4Mux_h
    port map (
            O => \N__36429\,
            I => \N__36426\
        );

    \I__6737\ : Odrv4
    port map (
            O => \N__36426\,
            I => n14564
        );

    \I__6736\ : InMux
    port map (
            O => \N__36423\,
            I => \N__36420\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__36420\,
            I => \N__36417\
        );

    \I__6734\ : Odrv4
    port map (
            O => \N__36417\,
            I => n1991
        );

    \I__6733\ : CascadeMux
    port map (
            O => \N__36414\,
            I => \N__36410\
        );

    \I__6732\ : CascadeMux
    port map (
            O => \N__36413\,
            I => \N__36407\
        );

    \I__6731\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36404\
        );

    \I__6730\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36401\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__36404\,
            I => \N__36398\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__36401\,
            I => \N__36394\
        );

    \I__6727\ : Span4Mux_h
    port map (
            O => \N__36398\,
            I => \N__36391\
        );

    \I__6726\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36388\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__36394\,
            I => n2023
        );

    \I__6724\ : Odrv4
    port map (
            O => \N__36391\,
            I => n2023
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__36388\,
            I => n2023
        );

    \I__6722\ : InMux
    port map (
            O => \N__36381\,
            I => \N__36378\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__36378\,
            I => \N__36375\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__36375\,
            I => n1994
        );

    \I__6719\ : CascadeMux
    port map (
            O => \N__36372\,
            I => \N__36368\
        );

    \I__6718\ : CascadeMux
    port map (
            O => \N__36371\,
            I => \N__36365\
        );

    \I__6717\ : InMux
    port map (
            O => \N__36368\,
            I => \N__36362\
        );

    \I__6716\ : InMux
    port map (
            O => \N__36365\,
            I => \N__36359\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__36362\,
            I => \N__36356\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__36359\,
            I => \N__36353\
        );

    \I__6713\ : Span4Mux_h
    port map (
            O => \N__36356\,
            I => \N__36349\
        );

    \I__6712\ : Span4Mux_h
    port map (
            O => \N__36353\,
            I => \N__36346\
        );

    \I__6711\ : InMux
    port map (
            O => \N__36352\,
            I => \N__36343\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__36349\,
            I => n2026
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__36346\,
            I => n2026
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__36343\,
            I => n2026
        );

    \I__6707\ : InMux
    port map (
            O => \N__36336\,
            I => \N__36333\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__36333\,
            I => n1993
        );

    \I__6705\ : InMux
    port map (
            O => \N__36330\,
            I => \N__36327\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__36327\,
            I => n1990
        );

    \I__6703\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36321\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__36321\,
            I => n1985
        );

    \I__6701\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36313\
        );

    \I__6700\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36308\
        );

    \I__6699\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36308\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__36313\,
            I => \N__36305\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__36308\,
            I => \N__36302\
        );

    \I__6696\ : Odrv4
    port map (
            O => \N__36305\,
            I => n2017
        );

    \I__6695\ : Odrv12
    port map (
            O => \N__36302\,
            I => n2017
        );

    \I__6694\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36294\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__36294\,
            I => n1992
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__36291\,
            I => \N__36288\
        );

    \I__6691\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36285\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__36285\,
            I => \N__36282\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__36282\,
            I => n1997
        );

    \I__6688\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36276\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__36276\,
            I => n1987
        );

    \I__6686\ : CascadeMux
    port map (
            O => \N__36273\,
            I => \N__36270\
        );

    \I__6685\ : InMux
    port map (
            O => \N__36270\,
            I => \N__36266\
        );

    \I__6684\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36263\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__36266\,
            I => \N__36260\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__36263\,
            I => \N__36256\
        );

    \I__6681\ : Span4Mux_h
    port map (
            O => \N__36260\,
            I => \N__36253\
        );

    \I__6680\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36250\
        );

    \I__6679\ : Odrv4
    port map (
            O => \N__36256\,
            I => n2025
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__36253\,
            I => n2025
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__36250\,
            I => n2025
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__36243\,
            I => \N__36239\
        );

    \I__6675\ : CascadeMux
    port map (
            O => \N__36242\,
            I => \N__36236\
        );

    \I__6674\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36233\
        );

    \I__6673\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36230\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__36233\,
            I => \N__36227\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__36230\,
            I => \N__36224\
        );

    \I__6670\ : Span4Mux_h
    port map (
            O => \N__36227\,
            I => \N__36220\
        );

    \I__6669\ : Span4Mux_h
    port map (
            O => \N__36224\,
            I => \N__36217\
        );

    \I__6668\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36214\
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__36220\,
            I => n2022
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__36217\,
            I => n2022
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__36214\,
            I => n2022
        );

    \I__6664\ : CascadeMux
    port map (
            O => \N__36207\,
            I => \N__36204\
        );

    \I__6663\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36200\
        );

    \I__6662\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36196\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__36200\,
            I => \N__36193\
        );

    \I__6660\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36190\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__36196\,
            I => \N__36187\
        );

    \I__6658\ : Span4Mux_h
    port map (
            O => \N__36193\,
            I => \N__36182\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__36190\,
            I => \N__36182\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__36187\,
            I => n2024
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__36182\,
            I => n2024
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__36177\,
            I => \n14550_cascade_\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__36174\,
            I => \N__36170\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__36173\,
            I => \N__36167\
        );

    \I__6651\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36164\
        );

    \I__6650\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36161\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__36164\,
            I => \N__36158\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__36161\,
            I => \N__36155\
        );

    \I__6647\ : Span4Mux_h
    port map (
            O => \N__36158\,
            I => \N__36151\
        );

    \I__6646\ : Span4Mux_h
    port map (
            O => \N__36155\,
            I => \N__36148\
        );

    \I__6645\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36145\
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__36151\,
            I => n2029
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__36148\,
            I => n2029
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__36145\,
            I => n2029
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__36138\,
            I => \n14556_cascade_\
        );

    \I__6640\ : InMux
    port map (
            O => \N__36135\,
            I => n12616
        );

    \I__6639\ : InMux
    port map (
            O => \N__36132\,
            I => n12617
        );

    \I__6638\ : InMux
    port map (
            O => \N__36129\,
            I => n12618
        );

    \I__6637\ : InMux
    port map (
            O => \N__36126\,
            I => n12619
        );

    \I__6636\ : InMux
    port map (
            O => \N__36123\,
            I => n12620
        );

    \I__6635\ : InMux
    port map (
            O => \N__36120\,
            I => n12621
        );

    \I__6634\ : CascadeMux
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__6633\ : InMux
    port map (
            O => \N__36114\,
            I => \N__36111\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__36111\,
            I => \N__36108\
        );

    \I__6631\ : Span4Mux_h
    port map (
            O => \N__36108\,
            I => \N__36105\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__36105\,
            I => n1986
        );

    \I__6629\ : InMux
    port map (
            O => \N__36102\,
            I => n12622
        );

    \I__6628\ : InMux
    port map (
            O => \N__36099\,
            I => \bfn_9_19_0_\
        );

    \I__6627\ : InMux
    port map (
            O => \N__36096\,
            I => n12624
        );

    \I__6626\ : InMux
    port map (
            O => \N__36093\,
            I => \N__36089\
        );

    \I__6625\ : InMux
    port map (
            O => \N__36092\,
            I => \N__36086\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__36089\,
            I => \N__36081\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__36086\,
            I => \N__36081\
        );

    \I__6622\ : Odrv12
    port map (
            O => \N__36081\,
            I => n2016
        );

    \I__6621\ : InMux
    port map (
            O => \N__36078\,
            I => \bfn_9_17_0_\
        );

    \I__6620\ : InMux
    port map (
            O => \N__36075\,
            I => n12608
        );

    \I__6619\ : InMux
    port map (
            O => \N__36072\,
            I => n12609
        );

    \I__6618\ : InMux
    port map (
            O => \N__36069\,
            I => n12610
        );

    \I__6617\ : InMux
    port map (
            O => \N__36066\,
            I => n12611
        );

    \I__6616\ : InMux
    port map (
            O => \N__36063\,
            I => n12612
        );

    \I__6615\ : InMux
    port map (
            O => \N__36060\,
            I => n12613
        );

    \I__6614\ : InMux
    port map (
            O => \N__36057\,
            I => n12614
        );

    \I__6613\ : InMux
    port map (
            O => \N__36054\,
            I => \bfn_9_18_0_\
        );

    \I__6612\ : InMux
    port map (
            O => \N__36051\,
            I => \N__36048\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__36048\,
            I => \N__36044\
        );

    \I__6610\ : InMux
    port map (
            O => \N__36047\,
            I => \N__36041\
        );

    \I__6609\ : Sp12to4
    port map (
            O => \N__36044\,
            I => \N__36036\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__36036\
        );

    \I__6607\ : Span12Mux_s5_v
    port map (
            O => \N__36036\,
            I => \N__36032\
        );

    \I__6606\ : InMux
    port map (
            O => \N__36035\,
            I => \N__36029\
        );

    \I__6605\ : Odrv12
    port map (
            O => \N__36032\,
            I => n3211
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__36029\,
            I => n3211
        );

    \I__6603\ : InMux
    port map (
            O => \N__36024\,
            I => \N__36021\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__36021\,
            I => n3278
        );

    \I__6601\ : InMux
    port map (
            O => \N__36018\,
            I => \bfn_7_32_0_\
        );

    \I__6600\ : InMux
    port map (
            O => \N__36015\,
            I => \N__36010\
        );

    \I__6599\ : InMux
    port map (
            O => \N__36014\,
            I => \N__36007\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__36013\,
            I => \N__36004\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__36010\,
            I => \N__36001\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__36007\,
            I => \N__35998\
        );

    \I__6595\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35995\
        );

    \I__6594\ : Span4Mux_s1_v
    port map (
            O => \N__36001\,
            I => \N__35992\
        );

    \I__6593\ : Span4Mux_s3_v
    port map (
            O => \N__35998\,
            I => \N__35987\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__35995\,
            I => \N__35987\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__35992\,
            I => n3210
        );

    \I__6590\ : Odrv4
    port map (
            O => \N__35987\,
            I => n3210
        );

    \I__6589\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35979\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__35979\,
            I => n3277
        );

    \I__6587\ : InMux
    port map (
            O => \N__35976\,
            I => n12931
        );

    \I__6586\ : InMux
    port map (
            O => \N__35973\,
            I => \N__35970\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__35970\,
            I => \N__35965\
        );

    \I__6584\ : InMux
    port map (
            O => \N__35969\,
            I => \N__35960\
        );

    \I__6583\ : InMux
    port map (
            O => \N__35968\,
            I => \N__35960\
        );

    \I__6582\ : Odrv12
    port map (
            O => \N__35965\,
            I => n3209
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__35960\,
            I => n3209
        );

    \I__6580\ : InMux
    port map (
            O => \N__35955\,
            I => \N__35952\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__35952\,
            I => \N__35949\
        );

    \I__6578\ : Span4Mux_v
    port map (
            O => \N__35949\,
            I => \N__35946\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__35946\,
            I => n3276
        );

    \I__6576\ : InMux
    port map (
            O => \N__35943\,
            I => n12932
        );

    \I__6575\ : InMux
    port map (
            O => \N__35940\,
            I => \N__35937\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__35937\,
            I => \N__35934\
        );

    \I__6573\ : Span4Mux_v
    port map (
            O => \N__35934\,
            I => \N__35931\
        );

    \I__6572\ : Odrv4
    port map (
            O => \N__35931\,
            I => n3275
        );

    \I__6571\ : InMux
    port map (
            O => \N__35928\,
            I => n12933
        );

    \I__6570\ : InMux
    port map (
            O => \N__35925\,
            I => \N__35922\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__6568\ : Span4Mux_s1_v
    port map (
            O => \N__35919\,
            I => \N__35914\
        );

    \I__6567\ : InMux
    port map (
            O => \N__35918\,
            I => \N__35909\
        );

    \I__6566\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35909\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__35914\,
            I => \N__35906\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__35909\,
            I => \N__35903\
        );

    \I__6563\ : Odrv4
    port map (
            O => \N__35906\,
            I => n3207
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__35903\,
            I => n3207
        );

    \I__6561\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35895\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__35895\,
            I => \N__35892\
        );

    \I__6559\ : Span4Mux_v
    port map (
            O => \N__35892\,
            I => \N__35889\
        );

    \I__6558\ : Span4Mux_v
    port map (
            O => \N__35889\,
            I => \N__35886\
        );

    \I__6557\ : Odrv4
    port map (
            O => \N__35886\,
            I => n3274
        );

    \I__6556\ : InMux
    port map (
            O => \N__35883\,
            I => n12934
        );

    \I__6555\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35876\
        );

    \I__6554\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35872\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__35876\,
            I => \N__35869\
        );

    \I__6552\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35866\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__35872\,
            I => \N__35863\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__35869\,
            I => \N__35860\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__35866\,
            I => \N__35857\
        );

    \I__6548\ : Odrv12
    port map (
            O => \N__35863\,
            I => n3206
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__35860\,
            I => n3206
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__35857\,
            I => n3206
        );

    \I__6545\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35847\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__35847\,
            I => n3273
        );

    \I__6543\ : InMux
    port map (
            O => \N__35844\,
            I => n12935
        );

    \I__6542\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35838\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__35838\,
            I => \N__35835\
        );

    \I__6540\ : Span4Mux_v
    port map (
            O => \N__35835\,
            I => \N__35830\
        );

    \I__6539\ : InMux
    port map (
            O => \N__35834\,
            I => \N__35825\
        );

    \I__6538\ : InMux
    port map (
            O => \N__35833\,
            I => \N__35825\
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__35830\,
            I => n3205
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__35825\,
            I => n3205
        );

    \I__6535\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35817\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__35817\,
            I => \N__35814\
        );

    \I__6533\ : Span4Mux_h
    port map (
            O => \N__35814\,
            I => \N__35811\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__35811\,
            I => \N__35808\
        );

    \I__6531\ : Odrv4
    port map (
            O => \N__35808\,
            I => n3272
        );

    \I__6530\ : InMux
    port map (
            O => \N__35805\,
            I => n12936
        );

    \I__6529\ : InMux
    port map (
            O => \N__35802\,
            I => \N__35798\
        );

    \I__6528\ : InMux
    port map (
            O => \N__35801\,
            I => \N__35795\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__35798\,
            I => \N__35792\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__35795\,
            I => \N__35789\
        );

    \I__6525\ : Span4Mux_s1_v
    port map (
            O => \N__35792\,
            I => \N__35786\
        );

    \I__6524\ : Odrv12
    port map (
            O => \N__35789\,
            I => n15450
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__35786\,
            I => n15450
        );

    \I__6522\ : CascadeMux
    port map (
            O => \N__35781\,
            I => \N__35778\
        );

    \I__6521\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35775\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35771\
        );

    \I__6519\ : InMux
    port map (
            O => \N__35774\,
            I => \N__35768\
        );

    \I__6518\ : Span4Mux_v
    port map (
            O => \N__35771\,
            I => \N__35765\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__35768\,
            I => \N__35762\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__35765\,
            I => n3204
        );

    \I__6515\ : Odrv4
    port map (
            O => \N__35762\,
            I => n3204
        );

    \I__6514\ : InMux
    port map (
            O => \N__35757\,
            I => n12937
        );

    \I__6513\ : InMux
    port map (
            O => \N__35754\,
            I => \N__35751\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__35751\,
            I => \N__35748\
        );

    \I__6511\ : Span4Mux_v
    port map (
            O => \N__35748\,
            I => \N__35745\
        );

    \I__6510\ : Span4Mux_v
    port map (
            O => \N__35745\,
            I => \N__35742\
        );

    \I__6509\ : Odrv4
    port map (
            O => \N__35742\,
            I => n14873
        );

    \I__6508\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35736\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__35736\,
            I => \N__35732\
        );

    \I__6506\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35729\
        );

    \I__6505\ : Span4Mux_h
    port map (
            O => \N__35732\,
            I => \N__35726\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__35729\,
            I => \N__35723\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__35726\,
            I => n3218
        );

    \I__6502\ : Odrv12
    port map (
            O => \N__35723\,
            I => n3218
        );

    \I__6501\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35715\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__35715\,
            I => n3285
        );

    \I__6499\ : InMux
    port map (
            O => \N__35712\,
            I => n12923
        );

    \I__6498\ : CascadeMux
    port map (
            O => \N__35709\,
            I => \N__35706\
        );

    \I__6497\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35701\
        );

    \I__6496\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35698\
        );

    \I__6495\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35695\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N__35692\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__35698\,
            I => \N__35689\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__35695\,
            I => \N__35686\
        );

    \I__6491\ : Odrv4
    port map (
            O => \N__35692\,
            I => n3217
        );

    \I__6490\ : Odrv4
    port map (
            O => \N__35689\,
            I => n3217
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__35686\,
            I => n3217
        );

    \I__6488\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35676\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__35676\,
            I => n3284
        );

    \I__6486\ : InMux
    port map (
            O => \N__35673\,
            I => n12924
        );

    \I__6485\ : InMux
    port map (
            O => \N__35670\,
            I => \N__35667\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__35667\,
            I => \N__35663\
        );

    \I__6483\ : InMux
    port map (
            O => \N__35666\,
            I => \N__35660\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__35663\,
            I => \N__35656\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__35660\,
            I => \N__35653\
        );

    \I__6480\ : InMux
    port map (
            O => \N__35659\,
            I => \N__35650\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__35656\,
            I => n3216
        );

    \I__6478\ : Odrv12
    port map (
            O => \N__35653\,
            I => n3216
        );

    \I__6477\ : LocalMux
    port map (
            O => \N__35650\,
            I => n3216
        );

    \I__6476\ : InMux
    port map (
            O => \N__35643\,
            I => \N__35640\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__35640\,
            I => n3283
        );

    \I__6474\ : InMux
    port map (
            O => \N__35637\,
            I => n12925
        );

    \I__6473\ : CascadeMux
    port map (
            O => \N__35634\,
            I => \N__35631\
        );

    \I__6472\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35627\
        );

    \I__6471\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35624\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__35627\,
            I => \N__35619\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__35624\,
            I => \N__35619\
        );

    \I__6468\ : Span4Mux_s3_v
    port map (
            O => \N__35619\,
            I => \N__35615\
        );

    \I__6467\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35612\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__35615\,
            I => n3215
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__35612\,
            I => n3215
        );

    \I__6464\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35604\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__35604\,
            I => n3282
        );

    \I__6462\ : InMux
    port map (
            O => \N__35601\,
            I => n12926
        );

    \I__6461\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35594\
        );

    \I__6460\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35591\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__35594\,
            I => \N__35588\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__35591\,
            I => \N__35585\
        );

    \I__6457\ : Span4Mux_v
    port map (
            O => \N__35588\,
            I => \N__35582\
        );

    \I__6456\ : Odrv12
    port map (
            O => \N__35585\,
            I => n3214
        );

    \I__6455\ : Odrv4
    port map (
            O => \N__35582\,
            I => n3214
        );

    \I__6454\ : InMux
    port map (
            O => \N__35577\,
            I => \N__35574\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__35574\,
            I => n3281
        );

    \I__6452\ : InMux
    port map (
            O => \N__35571\,
            I => n12927
        );

    \I__6451\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35564\
        );

    \I__6450\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35561\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__35564\,
            I => \N__35557\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35554\
        );

    \I__6447\ : InMux
    port map (
            O => \N__35560\,
            I => \N__35551\
        );

    \I__6446\ : Span4Mux_s1_v
    port map (
            O => \N__35557\,
            I => \N__35546\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__35554\,
            I => \N__35546\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35543\
        );

    \I__6443\ : Odrv4
    port map (
            O => \N__35546\,
            I => n3213
        );

    \I__6442\ : Odrv4
    port map (
            O => \N__35543\,
            I => n3213
        );

    \I__6441\ : CascadeMux
    port map (
            O => \N__35538\,
            I => \N__35535\
        );

    \I__6440\ : InMux
    port map (
            O => \N__35535\,
            I => \N__35532\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__35532\,
            I => n3280
        );

    \I__6438\ : InMux
    port map (
            O => \N__35529\,
            I => n12928
        );

    \I__6437\ : InMux
    port map (
            O => \N__35526\,
            I => \N__35521\
        );

    \I__6436\ : InMux
    port map (
            O => \N__35525\,
            I => \N__35518\
        );

    \I__6435\ : InMux
    port map (
            O => \N__35524\,
            I => \N__35515\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__35521\,
            I => \N__35512\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__35518\,
            I => \N__35509\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__35515\,
            I => \N__35506\
        );

    \I__6431\ : Span4Mux_s2_v
    port map (
            O => \N__35512\,
            I => \N__35503\
        );

    \I__6430\ : Span12Mux_s4_v
    port map (
            O => \N__35509\,
            I => \N__35500\
        );

    \I__6429\ : Span4Mux_h
    port map (
            O => \N__35506\,
            I => \N__35497\
        );

    \I__6428\ : Odrv4
    port map (
            O => \N__35503\,
            I => n3212
        );

    \I__6427\ : Odrv12
    port map (
            O => \N__35500\,
            I => n3212
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__35497\,
            I => n3212
        );

    \I__6425\ : InMux
    port map (
            O => \N__35490\,
            I => \N__35487\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__35487\,
            I => n3279
        );

    \I__6423\ : InMux
    port map (
            O => \N__35484\,
            I => n12929
        );

    \I__6422\ : InMux
    port map (
            O => \N__35481\,
            I => \N__35478\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__35478\,
            I => \N__35474\
        );

    \I__6420\ : InMux
    port map (
            O => \N__35477\,
            I => \N__35471\
        );

    \I__6419\ : Span4Mux_v
    port map (
            O => \N__35474\,
            I => \N__35465\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35465\
        );

    \I__6417\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35462\
        );

    \I__6416\ : Odrv4
    port map (
            O => \N__35465\,
            I => n3226
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__35462\,
            I => n3226
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__35457\,
            I => \N__35454\
        );

    \I__6413\ : InMux
    port map (
            O => \N__35454\,
            I => \N__35451\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__35451\,
            I => \N__35448\
        );

    \I__6411\ : Span4Mux_h
    port map (
            O => \N__35448\,
            I => \N__35445\
        );

    \I__6410\ : Span4Mux_v
    port map (
            O => \N__35445\,
            I => \N__35442\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__35442\,
            I => n3293
        );

    \I__6408\ : InMux
    port map (
            O => \N__35439\,
            I => n12915
        );

    \I__6407\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35432\
        );

    \I__6406\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35429\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__35432\,
            I => \N__35426\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35423\
        );

    \I__6403\ : Span4Mux_s3_v
    port map (
            O => \N__35426\,
            I => \N__35420\
        );

    \I__6402\ : Odrv4
    port map (
            O => \N__35423\,
            I => n3225
        );

    \I__6401\ : Odrv4
    port map (
            O => \N__35420\,
            I => n3225
        );

    \I__6400\ : InMux
    port map (
            O => \N__35415\,
            I => \N__35412\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__35412\,
            I => \N__35409\
        );

    \I__6398\ : Span4Mux_v
    port map (
            O => \N__35409\,
            I => \N__35406\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__35406\,
            I => n3292
        );

    \I__6396\ : InMux
    port map (
            O => \N__35403\,
            I => n12916
        );

    \I__6395\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35396\
        );

    \I__6394\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35393\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__35396\,
            I => \N__35389\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__35393\,
            I => \N__35386\
        );

    \I__6391\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35383\
        );

    \I__6390\ : Odrv4
    port map (
            O => \N__35389\,
            I => n3224
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__35386\,
            I => n3224
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__35383\,
            I => n3224
        );

    \I__6387\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35373\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__35373\,
            I => \N__35370\
        );

    \I__6385\ : Span4Mux_v
    port map (
            O => \N__35370\,
            I => \N__35367\
        );

    \I__6384\ : Span4Mux_v
    port map (
            O => \N__35367\,
            I => \N__35364\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__35364\,
            I => n3291
        );

    \I__6382\ : InMux
    port map (
            O => \N__35361\,
            I => n12917
        );

    \I__6381\ : InMux
    port map (
            O => \N__35358\,
            I => \N__35354\
        );

    \I__6380\ : InMux
    port map (
            O => \N__35357\,
            I => \N__35351\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__35354\,
            I => \N__35345\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__35351\,
            I => \N__35345\
        );

    \I__6377\ : InMux
    port map (
            O => \N__35350\,
            I => \N__35342\
        );

    \I__6376\ : Odrv4
    port map (
            O => \N__35345\,
            I => n3223
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__35342\,
            I => n3223
        );

    \I__6374\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35334\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__35334\,
            I => n3290
        );

    \I__6372\ : InMux
    port map (
            O => \N__35331\,
            I => n12918
        );

    \I__6371\ : InMux
    port map (
            O => \N__35328\,
            I => \N__35325\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__35325\,
            I => \N__35322\
        );

    \I__6369\ : Span4Mux_s3_v
    port map (
            O => \N__35322\,
            I => \N__35318\
        );

    \I__6368\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35315\
        );

    \I__6367\ : Odrv4
    port map (
            O => \N__35318\,
            I => n3222
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__35315\,
            I => n3222
        );

    \I__6365\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35307\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__35307\,
            I => \N__35304\
        );

    \I__6363\ : Span4Mux_h
    port map (
            O => \N__35304\,
            I => \N__35301\
        );

    \I__6362\ : Odrv4
    port map (
            O => \N__35301\,
            I => n3289
        );

    \I__6361\ : InMux
    port map (
            O => \N__35298\,
            I => n12919
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__35295\,
            I => \N__35292\
        );

    \I__6359\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35288\
        );

    \I__6358\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35285\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__35288\,
            I => \N__35282\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__35285\,
            I => n3221
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__35282\,
            I => n3221
        );

    \I__6354\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35274\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__35274\,
            I => \N__35271\
        );

    \I__6352\ : Odrv12
    port map (
            O => \N__35271\,
            I => n3288
        );

    \I__6351\ : InMux
    port map (
            O => \N__35268\,
            I => n12920
        );

    \I__6350\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35262\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__35262\,
            I => \N__35257\
        );

    \I__6348\ : InMux
    port map (
            O => \N__35261\,
            I => \N__35252\
        );

    \I__6347\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35252\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__35257\,
            I => n3220
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__35252\,
            I => n3220
        );

    \I__6344\ : CascadeMux
    port map (
            O => \N__35247\,
            I => \N__35244\
        );

    \I__6343\ : InMux
    port map (
            O => \N__35244\,
            I => \N__35241\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__35241\,
            I => \N__35238\
        );

    \I__6341\ : Odrv12
    port map (
            O => \N__35238\,
            I => n3287
        );

    \I__6340\ : InMux
    port map (
            O => \N__35235\,
            I => n12921
        );

    \I__6339\ : InMux
    port map (
            O => \N__35232\,
            I => \N__35228\
        );

    \I__6338\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35225\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__35228\,
            I => \N__35222\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__35225\,
            I => \N__35218\
        );

    \I__6335\ : Span4Mux_s3_v
    port map (
            O => \N__35222\,
            I => \N__35215\
        );

    \I__6334\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35212\
        );

    \I__6333\ : Odrv4
    port map (
            O => \N__35218\,
            I => n3219
        );

    \I__6332\ : Odrv4
    port map (
            O => \N__35215\,
            I => n3219
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__35212\,
            I => n3219
        );

    \I__6330\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35202\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__35202\,
            I => \N__35199\
        );

    \I__6328\ : Span4Mux_v
    port map (
            O => \N__35199\,
            I => \N__35196\
        );

    \I__6327\ : Odrv4
    port map (
            O => \N__35196\,
            I => n3286
        );

    \I__6326\ : InMux
    port map (
            O => \N__35193\,
            I => \bfn_7_31_0_\
        );

    \I__6325\ : InMux
    port map (
            O => \N__35190\,
            I => \N__35187\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__35187\,
            I => \N__35184\
        );

    \I__6323\ : Span4Mux_h
    port map (
            O => \N__35184\,
            I => \N__35181\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__35181\,
            I => n3301
        );

    \I__6321\ : InMux
    port map (
            O => \N__35178\,
            I => n12907
        );

    \I__6320\ : InMux
    port map (
            O => \N__35175\,
            I => \N__35171\
        );

    \I__6319\ : InMux
    port map (
            O => \N__35174\,
            I => \N__35168\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__35171\,
            I => n3233
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__35168\,
            I => n3233
        );

    \I__6316\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35160\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__35160\,
            I => n3300
        );

    \I__6314\ : InMux
    port map (
            O => \N__35157\,
            I => n12908
        );

    \I__6313\ : InMux
    port map (
            O => \N__35154\,
            I => \N__35151\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__35151\,
            I => \N__35147\
        );

    \I__6311\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35144\
        );

    \I__6310\ : Odrv12
    port map (
            O => \N__35147\,
            I => n3232
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__35144\,
            I => n3232
        );

    \I__6308\ : InMux
    port map (
            O => \N__35139\,
            I => \N__35136\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__35136\,
            I => \N__35133\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__35133\,
            I => n3299
        );

    \I__6305\ : InMux
    port map (
            O => \N__35130\,
            I => n12909
        );

    \I__6304\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35122\
        );

    \I__6303\ : InMux
    port map (
            O => \N__35126\,
            I => \N__35119\
        );

    \I__6302\ : InMux
    port map (
            O => \N__35125\,
            I => \N__35116\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__35122\,
            I => n3231
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__35119\,
            I => n3231
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__35116\,
            I => n3231
        );

    \I__6298\ : InMux
    port map (
            O => \N__35109\,
            I => n12910
        );

    \I__6297\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35103\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__35103\,
            I => n3298
        );

    \I__6295\ : InMux
    port map (
            O => \N__35100\,
            I => \N__35095\
        );

    \I__6294\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35092\
        );

    \I__6293\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35089\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__35095\,
            I => \N__35086\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__35092\,
            I => n3230
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__35089\,
            I => n3230
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__35086\,
            I => n3230
        );

    \I__6288\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35076\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__35076\,
            I => n15097
        );

    \I__6286\ : InMux
    port map (
            O => \N__35073\,
            I => n12911
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__35070\,
            I => \N__35066\
        );

    \I__6284\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35063\
        );

    \I__6283\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35060\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__35063\,
            I => n3229
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__35060\,
            I => n3229
        );

    \I__6280\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35052\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__35052\,
            I => n3296
        );

    \I__6278\ : InMux
    port map (
            O => \N__35049\,
            I => n12912
        );

    \I__6277\ : InMux
    port map (
            O => \N__35046\,
            I => \N__35043\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__35043\,
            I => \N__35038\
        );

    \I__6275\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35035\
        );

    \I__6274\ : InMux
    port map (
            O => \N__35041\,
            I => \N__35032\
        );

    \I__6273\ : Odrv4
    port map (
            O => \N__35038\,
            I => n3228
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__35035\,
            I => n3228
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__35032\,
            I => n3228
        );

    \I__6270\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__35022\,
            I => n3295
        );

    \I__6268\ : InMux
    port map (
            O => \N__35019\,
            I => n12913
        );

    \I__6267\ : InMux
    port map (
            O => \N__35016\,
            I => \N__35012\
        );

    \I__6266\ : InMux
    port map (
            O => \N__35015\,
            I => \N__35009\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__35012\,
            I => \N__35005\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__35002\
        );

    \I__6263\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34999\
        );

    \I__6262\ : Odrv4
    port map (
            O => \N__35005\,
            I => n3227
        );

    \I__6261\ : Odrv12
    port map (
            O => \N__35002\,
            I => n3227
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__34999\,
            I => n3227
        );

    \I__6259\ : CascadeMux
    port map (
            O => \N__34992\,
            I => \N__34989\
        );

    \I__6258\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34986\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__34986\,
            I => \N__34983\
        );

    \I__6256\ : Span4Mux_h
    port map (
            O => \N__34983\,
            I => \N__34980\
        );

    \I__6255\ : Span4Mux_v
    port map (
            O => \N__34980\,
            I => \N__34977\
        );

    \I__6254\ : Odrv4
    port map (
            O => \N__34977\,
            I => n3294
        );

    \I__6253\ : InMux
    port map (
            O => \N__34974\,
            I => \bfn_7_30_0_\
        );

    \I__6252\ : CascadeMux
    port map (
            O => \N__34971\,
            I => \N__34968\
        );

    \I__6251\ : InMux
    port map (
            O => \N__34968\,
            I => \N__34965\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__34965\,
            I => \N__34962\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__34962\,
            I => \N__34959\
        );

    \I__6248\ : Odrv4
    port map (
            O => \N__34959\,
            I => n3080
        );

    \I__6247\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34953\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__34953\,
            I => \N__34949\
        );

    \I__6245\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34945\
        );

    \I__6244\ : Span4Mux_v
    port map (
            O => \N__34949\,
            I => \N__34942\
        );

    \I__6243\ : InMux
    port map (
            O => \N__34948\,
            I => \N__34939\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__34945\,
            I => n3112
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__34942\,
            I => n3112
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__34939\,
            I => n3112
        );

    \I__6239\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34929\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__34929\,
            I => \N__34926\
        );

    \I__6237\ : Span4Mux_h
    port map (
            O => \N__34926\,
            I => \N__34923\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__34923\,
            I => n3192
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__34920\,
            I => \N__34917\
        );

    \I__6234\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34913\
        );

    \I__6233\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34910\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34907\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__34910\,
            I => \N__34903\
        );

    \I__6230\ : Span4Mux_v
    port map (
            O => \N__34907\,
            I => \N__34900\
        );

    \I__6229\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34897\
        );

    \I__6228\ : Odrv4
    port map (
            O => \N__34903\,
            I => n3125
        );

    \I__6227\ : Odrv4
    port map (
            O => \N__34900\,
            I => n3125
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__34897\,
            I => n3125
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__34890\,
            I => \N__34887\
        );

    \I__6224\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34884\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__34884\,
            I => \N__34881\
        );

    \I__6222\ : Span4Mux_h
    port map (
            O => \N__34881\,
            I => \N__34878\
        );

    \I__6221\ : Odrv4
    port map (
            O => \N__34878\,
            I => n3196
        );

    \I__6220\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34871\
        );

    \I__6219\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34868\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__34871\,
            I => \N__34865\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__34868\,
            I => \N__34860\
        );

    \I__6216\ : Span4Mux_h
    port map (
            O => \N__34865\,
            I => \N__34860\
        );

    \I__6215\ : Span4Mux_h
    port map (
            O => \N__34860\,
            I => \N__34857\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__34857\,
            I => \debounce.reg_A_0\
        );

    \I__6213\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34850\
        );

    \I__6212\ : CascadeMux
    port map (
            O => \N__34853\,
            I => \N__34847\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__34850\,
            I => \N__34844\
        );

    \I__6210\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34841\
        );

    \I__6209\ : Span4Mux_s3_h
    port map (
            O => \N__34844\,
            I => \N__34838\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__34841\,
            I => \N__34835\
        );

    \I__6207\ : Span4Mux_v
    port map (
            O => \N__34838\,
            I => \N__34832\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__34835\,
            I => \N__34829\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__34832\,
            I => \reg_B_0\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__34829\,
            I => \reg_B_0\
        );

    \I__6203\ : InMux
    port map (
            O => \N__34824\,
            I => \N__34820\
        );

    \I__6202\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34817\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34814\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__34817\,
            I => \debounce.reg_A_1\
        );

    \I__6199\ : Odrv12
    port map (
            O => \N__34814\,
            I => \debounce.reg_A_1\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__34809\,
            I => \N__34806\
        );

    \I__6197\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34803\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34800\
        );

    \I__6195\ : Span4Mux_v
    port map (
            O => \N__34800\,
            I => \N__34797\
        );

    \I__6194\ : Odrv4
    port map (
            O => \N__34797\,
            I => \debounce.n6\
        );

    \I__6193\ : InMux
    port map (
            O => \N__34794\,
            I => \N__34791\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__34791\,
            I => \N__34788\
        );

    \I__6191\ : Span4Mux_h
    port map (
            O => \N__34788\,
            I => \N__34785\
        );

    \I__6190\ : Odrv4
    port map (
            O => \N__34785\,
            I => n3185
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__34782\,
            I => \N__34777\
        );

    \I__6188\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34774\
        );

    \I__6187\ : InMux
    port map (
            O => \N__34780\,
            I => \N__34771\
        );

    \I__6186\ : InMux
    port map (
            O => \N__34777\,
            I => \N__34768\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__34774\,
            I => \N__34765\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34762\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34759\
        );

    \I__6182\ : Span4Mux_h
    port map (
            O => \N__34765\,
            I => \N__34752\
        );

    \I__6181\ : Span4Mux_v
    port map (
            O => \N__34762\,
            I => \N__34752\
        );

    \I__6180\ : Span4Mux_v
    port map (
            O => \N__34759\,
            I => \N__34752\
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__34752\,
            I => n3118
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__34749\,
            I => \N__34746\
        );

    \I__6177\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34743\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__34743\,
            I => \N__34740\
        );

    \I__6175\ : Span4Mux_h
    port map (
            O => \N__34740\,
            I => \N__34737\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__34737\,
            I => n3197
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__34734\,
            I => \n3229_cascade_\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__34731\,
            I => \N__34722\
        );

    \I__6171\ : CascadeMux
    port map (
            O => \N__34730\,
            I => \N__34717\
        );

    \I__6170\ : CascadeMux
    port map (
            O => \N__34729\,
            I => \N__34712\
        );

    \I__6169\ : CascadeMux
    port map (
            O => \N__34728\,
            I => \N__34709\
        );

    \I__6168\ : CascadeMux
    port map (
            O => \N__34727\,
            I => \N__34704\
        );

    \I__6167\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34696\
        );

    \I__6166\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34687\
        );

    \I__6165\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34687\
        );

    \I__6164\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34687\
        );

    \I__6163\ : InMux
    port map (
            O => \N__34720\,
            I => \N__34687\
        );

    \I__6162\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34678\
        );

    \I__6161\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34678\
        );

    \I__6160\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34678\
        );

    \I__6159\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34678\
        );

    \I__6158\ : InMux
    port map (
            O => \N__34709\,
            I => \N__34665\
        );

    \I__6157\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34665\
        );

    \I__6156\ : InMux
    port map (
            O => \N__34707\,
            I => \N__34665\
        );

    \I__6155\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34665\
        );

    \I__6154\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34665\
        );

    \I__6153\ : InMux
    port map (
            O => \N__34702\,
            I => \N__34665\
        );

    \I__6152\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34660\
        );

    \I__6151\ : CascadeMux
    port map (
            O => \N__34700\,
            I => \N__34657\
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__34699\,
            I => \N__34652\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__34696\,
            I => \N__34648\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__34687\,
            I => \N__34641\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__34678\,
            I => \N__34641\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__34665\,
            I => \N__34641\
        );

    \I__6145\ : InMux
    port map (
            O => \N__34664\,
            I => \N__34636\
        );

    \I__6144\ : InMux
    port map (
            O => \N__34663\,
            I => \N__34636\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__34660\,
            I => \N__34626\
        );

    \I__6142\ : InMux
    port map (
            O => \N__34657\,
            I => \N__34615\
        );

    \I__6141\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34615\
        );

    \I__6140\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34615\
        );

    \I__6139\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34615\
        );

    \I__6138\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34615\
        );

    \I__6137\ : Span4Mux_h
    port map (
            O => \N__34648\,
            I => \N__34608\
        );

    \I__6136\ : Span4Mux_v
    port map (
            O => \N__34641\,
            I => \N__34608\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34608\
        );

    \I__6134\ : InMux
    port map (
            O => \N__34635\,
            I => \N__34599\
        );

    \I__6133\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34599\
        );

    \I__6132\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34599\
        );

    \I__6131\ : InMux
    port map (
            O => \N__34632\,
            I => \N__34599\
        );

    \I__6130\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34594\
        );

    \I__6129\ : InMux
    port map (
            O => \N__34630\,
            I => \N__34594\
        );

    \I__6128\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34591\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__34626\,
            I => n3237
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__34615\,
            I => n3237
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__34608\,
            I => n3237
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__34599\,
            I => n3237
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__34594\,
            I => n3237
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__34591\,
            I => n3237
        );

    \I__6121\ : CascadeMux
    port map (
            O => \N__34578\,
            I => \N__34575\
        );

    \I__6120\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34572\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__34572\,
            I => \N__34569\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__34569\,
            I => n13_adj_709
        );

    \I__6117\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34562\
        );

    \I__6116\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34559\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__34562\,
            I => \N__34556\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__34559\,
            I => \N__34551\
        );

    \I__6113\ : Span4Mux_v
    port map (
            O => \N__34556\,
            I => \N__34551\
        );

    \I__6112\ : Odrv4
    port map (
            O => \N__34551\,
            I => n319
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__34548\,
            I => \n14780_cascade_\
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__34545\,
            I => \N__34541\
        );

    \I__6109\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34538\
        );

    \I__6108\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34535\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34531\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__34535\,
            I => \N__34528\
        );

    \I__6105\ : InMux
    port map (
            O => \N__34534\,
            I => \N__34525\
        );

    \I__6104\ : Span4Mux_h
    port map (
            O => \N__34531\,
            I => \N__34522\
        );

    \I__6103\ : Span4Mux_v
    port map (
            O => \N__34528\,
            I => \N__34517\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__34525\,
            I => \N__34517\
        );

    \I__6101\ : Odrv4
    port map (
            O => \N__34522\,
            I => n3128
        );

    \I__6100\ : Odrv4
    port map (
            O => \N__34517\,
            I => n3128
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__34512\,
            I => \N__34509\
        );

    \I__6098\ : InMux
    port map (
            O => \N__34509\,
            I => \N__34506\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__34506\,
            I => \N__34503\
        );

    \I__6096\ : Span4Mux_h
    port map (
            O => \N__34503\,
            I => \N__34500\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__34500\,
            I => n3195
        );

    \I__6094\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34493\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__34496\,
            I => \N__34490\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__34493\,
            I => \N__34487\
        );

    \I__6091\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34484\
        );

    \I__6090\ : Span4Mux_h
    port map (
            O => \N__34487\,
            I => \N__34481\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__34484\,
            I => \N__34478\
        );

    \I__6088\ : Span4Mux_v
    port map (
            O => \N__34481\,
            I => \N__34475\
        );

    \I__6087\ : Span4Mux_v
    port map (
            O => \N__34478\,
            I => \N__34472\
        );

    \I__6086\ : Odrv4
    port map (
            O => \N__34475\,
            I => n3117
        );

    \I__6085\ : Odrv4
    port map (
            O => \N__34472\,
            I => n3117
        );

    \I__6084\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34464\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__34464\,
            I => \N__34461\
        );

    \I__6082\ : Odrv4
    port map (
            O => \N__34461\,
            I => n3184
        );

    \I__6081\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34454\
        );

    \I__6080\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34451\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__34454\,
            I => \N__34448\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__34451\,
            I => \N__34445\
        );

    \I__6077\ : Span4Mux_h
    port map (
            O => \N__34448\,
            I => \N__34441\
        );

    \I__6076\ : Span4Mux_v
    port map (
            O => \N__34445\,
            I => \N__34438\
        );

    \I__6075\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34435\
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__34441\,
            I => n3119
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__34438\,
            I => n3119
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__34435\,
            I => n3119
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__34428\,
            I => \N__34425\
        );

    \I__6070\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34422\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__34422\,
            I => \N__34419\
        );

    \I__6068\ : Span4Mux_h
    port map (
            O => \N__34419\,
            I => \N__34416\
        );

    \I__6067\ : Odrv4
    port map (
            O => \N__34416\,
            I => n3186
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__34413\,
            I => \n3218_cascade_\
        );

    \I__6065\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34407\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__34407\,
            I => n14778
        );

    \I__6063\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34401\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__34401\,
            I => \N__34398\
        );

    \I__6061\ : Odrv4
    port map (
            O => \N__34398\,
            I => n12030
        );

    \I__6060\ : InMux
    port map (
            O => \N__34395\,
            I => \N__34392\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__34392\,
            I => n14786
        );

    \I__6058\ : InMux
    port map (
            O => \N__34389\,
            I => \N__34386\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__34386\,
            I => n14788
        );

    \I__6056\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34380\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__34380\,
            I => \N__34377\
        );

    \I__6054\ : Odrv4
    port map (
            O => \N__34377\,
            I => encoder0_position_scaled_12
        );

    \I__6053\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34371\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__34371\,
            I => \N__34368\
        );

    \I__6051\ : Span4Mux_h
    port map (
            O => \N__34368\,
            I => \N__34365\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__34365\,
            I => n3194
        );

    \I__6049\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34358\
        );

    \I__6048\ : CascadeMux
    port map (
            O => \N__34361\,
            I => \N__34355\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__34358\,
            I => \N__34352\
        );

    \I__6046\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34349\
        );

    \I__6045\ : Span4Mux_h
    port map (
            O => \N__34352\,
            I => \N__34346\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34343\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__34346\,
            I => n3127
        );

    \I__6042\ : Odrv12
    port map (
            O => \N__34343\,
            I => n3127
        );

    \I__6041\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34335\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__34335\,
            I => \N__34332\
        );

    \I__6039\ : Span4Mux_h
    port map (
            O => \N__34332\,
            I => \N__34327\
        );

    \I__6038\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34324\
        );

    \I__6037\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34321\
        );

    \I__6036\ : Odrv4
    port map (
            O => \N__34327\,
            I => n3013
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__34324\,
            I => n3013
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__34321\,
            I => n3013
        );

    \I__6033\ : InMux
    port map (
            O => \N__34314\,
            I => n12958
        );

    \I__6032\ : InMux
    port map (
            O => \N__34311\,
            I => n12959
        );

    \I__6031\ : InMux
    port map (
            O => \N__34308\,
            I => n12960
        );

    \I__6030\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34302\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__34302\,
            I => \N__34299\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__34299\,
            I => \N__34296\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__34296\,
            I => n3177
        );

    \I__6026\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34289\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__34292\,
            I => \N__34286\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__34289\,
            I => \N__34282\
        );

    \I__6023\ : InMux
    port map (
            O => \N__34286\,
            I => \N__34279\
        );

    \I__6022\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34276\
        );

    \I__6021\ : Span4Mux_h
    port map (
            O => \N__34282\,
            I => \N__34273\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__34279\,
            I => \N__34268\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__34276\,
            I => \N__34268\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__34273\,
            I => \N__34265\
        );

    \I__6017\ : Span4Mux_h
    port map (
            O => \N__34268\,
            I => \N__34262\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__34265\,
            I => n3110
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__34262\,
            I => n3110
        );

    \I__6014\ : CascadeMux
    port map (
            O => \N__34257\,
            I => \n31_adj_714_cascade_\
        );

    \I__6013\ : InMux
    port map (
            O => \N__34254\,
            I => \N__34251\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__34251\,
            I => \N__34248\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__34248\,
            I => n14232
        );

    \I__6010\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34240\
        );

    \I__6009\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34237\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__34243\,
            I => \N__34234\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__34240\,
            I => \N__34231\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__34237\,
            I => \N__34228\
        );

    \I__6005\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34225\
        );

    \I__6004\ : Span4Mux_s3_v
    port map (
            O => \N__34231\,
            I => \N__34222\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__34228\,
            I => n3126
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__34225\,
            I => n3126
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__34222\,
            I => n3126
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__34215\,
            I => \N__34212\
        );

    \I__5999\ : InMux
    port map (
            O => \N__34212\,
            I => \N__34209\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__34209\,
            I => \N__34206\
        );

    \I__5997\ : Odrv4
    port map (
            O => \N__34206\,
            I => n3193
        );

    \I__5996\ : CascadeMux
    port map (
            O => \N__34203\,
            I => \n3225_cascade_\
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__34200\,
            I => \n14776_cascade_\
        );

    \I__5994\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__34194\,
            I => n14764
        );

    \I__5992\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34188\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__34188\,
            I => \N__34185\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__34185\,
            I => \N__34181\
        );

    \I__5989\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34178\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__34181\,
            I => \N__34173\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__34178\,
            I => \N__34173\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__34173\,
            I => n15714
        );

    \I__5985\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34164\
        );

    \I__5984\ : CascadeMux
    port map (
            O => \N__34169\,
            I => \N__34156\
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__34168\,
            I => \N__34149\
        );

    \I__5982\ : CascadeMux
    port map (
            O => \N__34167\,
            I => \N__34145\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__34164\,
            I => \N__34141\
        );

    \I__5980\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34138\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__34162\,
            I => \N__34134\
        );

    \I__5978\ : CascadeMux
    port map (
            O => \N__34161\,
            I => \N__34130\
        );

    \I__5977\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34122\
        );

    \I__5976\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34122\
        );

    \I__5975\ : InMux
    port map (
            O => \N__34156\,
            I => \N__34119\
        );

    \I__5974\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34114\
        );

    \I__5973\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34114\
        );

    \I__5972\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34109\
        );

    \I__5971\ : InMux
    port map (
            O => \N__34152\,
            I => \N__34109\
        );

    \I__5970\ : InMux
    port map (
            O => \N__34149\,
            I => \N__34104\
        );

    \I__5969\ : InMux
    port map (
            O => \N__34148\,
            I => \N__34104\
        );

    \I__5968\ : InMux
    port map (
            O => \N__34145\,
            I => \N__34099\
        );

    \I__5967\ : InMux
    port map (
            O => \N__34144\,
            I => \N__34099\
        );

    \I__5966\ : Span4Mux_v
    port map (
            O => \N__34141\,
            I => \N__34094\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34094\
        );

    \I__5964\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34081\
        );

    \I__5963\ : InMux
    port map (
            O => \N__34134\,
            I => \N__34081\
        );

    \I__5962\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34081\
        );

    \I__5961\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34081\
        );

    \I__5960\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34081\
        );

    \I__5959\ : InMux
    port map (
            O => \N__34128\,
            I => \N__34081\
        );

    \I__5958\ : InMux
    port map (
            O => \N__34127\,
            I => \N__34078\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__34122\,
            I => \N__34075\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__34119\,
            I => \N__34070\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__34114\,
            I => \N__34070\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__34109\,
            I => n2148
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__34104\,
            I => n2148
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__34099\,
            I => n2148
        );

    \I__5951\ : Odrv4
    port map (
            O => \N__34094\,
            I => n2148
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__34081\,
            I => n2148
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__34078\,
            I => n2148
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__34075\,
            I => n2148
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__34070\,
            I => n2148
        );

    \I__5946\ : InMux
    port map (
            O => \N__34053\,
            I => n12949
        );

    \I__5945\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34047\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__34047\,
            I => \N__34043\
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__34046\,
            I => \N__34040\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__34043\,
            I => \N__34037\
        );

    \I__5941\ : InMux
    port map (
            O => \N__34040\,
            I => \N__34034\
        );

    \I__5940\ : Odrv4
    port map (
            O => \N__34037\,
            I => n15689
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__34034\,
            I => n15689
        );

    \I__5938\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34021\
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__34028\,
            I => \N__34012\
        );

    \I__5936\ : CascadeMux
    port map (
            O => \N__34027\,
            I => \N__34007\
        );

    \I__5935\ : CascadeMux
    port map (
            O => \N__34026\,
            I => \N__34004\
        );

    \I__5934\ : InMux
    port map (
            O => \N__34025\,
            I => \N__33997\
        );

    \I__5933\ : InMux
    port map (
            O => \N__34024\,
            I => \N__33997\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__34021\,
            I => \N__33994\
        );

    \I__5931\ : InMux
    port map (
            O => \N__34020\,
            I => \N__33989\
        );

    \I__5930\ : InMux
    port map (
            O => \N__34019\,
            I => \N__33989\
        );

    \I__5929\ : InMux
    port map (
            O => \N__34018\,
            I => \N__33986\
        );

    \I__5928\ : CascadeMux
    port map (
            O => \N__34017\,
            I => \N__33981\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__34016\,
            I => \N__33978\
        );

    \I__5926\ : InMux
    port map (
            O => \N__34015\,
            I => \N__33974\
        );

    \I__5925\ : InMux
    port map (
            O => \N__34012\,
            I => \N__33967\
        );

    \I__5924\ : InMux
    port map (
            O => \N__34011\,
            I => \N__33967\
        );

    \I__5923\ : InMux
    port map (
            O => \N__34010\,
            I => \N__33967\
        );

    \I__5922\ : InMux
    port map (
            O => \N__34007\,
            I => \N__33958\
        );

    \I__5921\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33958\
        );

    \I__5920\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33958\
        );

    \I__5919\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33958\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__33997\,
            I => \N__33955\
        );

    \I__5917\ : Span4Mux_v
    port map (
            O => \N__33994\,
            I => \N__33948\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__33989\,
            I => \N__33948\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__33986\,
            I => \N__33948\
        );

    \I__5914\ : InMux
    port map (
            O => \N__33985\,
            I => \N__33943\
        );

    \I__5913\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33943\
        );

    \I__5912\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33936\
        );

    \I__5911\ : InMux
    port map (
            O => \N__33978\,
            I => \N__33936\
        );

    \I__5910\ : InMux
    port map (
            O => \N__33977\,
            I => \N__33936\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__33974\,
            I => n2049
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__33967\,
            I => n2049
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__33958\,
            I => n2049
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__33955\,
            I => n2049
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__33948\,
            I => n2049
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__33943\,
            I => n2049
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__33936\,
            I => n2049
        );

    \I__5902\ : InMux
    port map (
            O => \N__33921\,
            I => n12950
        );

    \I__5901\ : InMux
    port map (
            O => \N__33918\,
            I => n12951
        );

    \I__5900\ : InMux
    port map (
            O => \N__33915\,
            I => n12952
        );

    \I__5899\ : InMux
    port map (
            O => \N__33912\,
            I => \bfn_7_25_0_\
        );

    \I__5898\ : InMux
    port map (
            O => \N__33909\,
            I => n12954
        );

    \I__5897\ : InMux
    port map (
            O => \N__33906\,
            I => n12955
        );

    \I__5896\ : InMux
    port map (
            O => \N__33903\,
            I => n12956
        );

    \I__5895\ : InMux
    port map (
            O => \N__33900\,
            I => n12957
        );

    \I__5894\ : InMux
    port map (
            O => \N__33897\,
            I => \N__33888\
        );

    \I__5893\ : InMux
    port map (
            O => \N__33896\,
            I => \N__33881\
        );

    \I__5892\ : InMux
    port map (
            O => \N__33895\,
            I => \N__33881\
        );

    \I__5891\ : InMux
    port map (
            O => \N__33894\,
            I => \N__33874\
        );

    \I__5890\ : InMux
    port map (
            O => \N__33893\,
            I => \N__33874\
        );

    \I__5889\ : InMux
    port map (
            O => \N__33892\,
            I => \N__33874\
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__33891\,
            I => \N__33868\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__33888\,
            I => \N__33859\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__33887\,
            I => \N__33855\
        );

    \I__5885\ : InMux
    port map (
            O => \N__33886\,
            I => \N__33851\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__33881\,
            I => \N__33846\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__33874\,
            I => \N__33841\
        );

    \I__5882\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33830\
        );

    \I__5881\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33830\
        );

    \I__5880\ : InMux
    port map (
            O => \N__33871\,
            I => \N__33830\
        );

    \I__5879\ : InMux
    port map (
            O => \N__33868\,
            I => \N__33830\
        );

    \I__5878\ : InMux
    port map (
            O => \N__33867\,
            I => \N__33830\
        );

    \I__5877\ : InMux
    port map (
            O => \N__33866\,
            I => \N__33825\
        );

    \I__5876\ : InMux
    port map (
            O => \N__33865\,
            I => \N__33825\
        );

    \I__5875\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33818\
        );

    \I__5874\ : InMux
    port map (
            O => \N__33863\,
            I => \N__33818\
        );

    \I__5873\ : InMux
    port map (
            O => \N__33862\,
            I => \N__33818\
        );

    \I__5872\ : Span4Mux_v
    port map (
            O => \N__33859\,
            I => \N__33815\
        );

    \I__5871\ : InMux
    port map (
            O => \N__33858\,
            I => \N__33808\
        );

    \I__5870\ : InMux
    port map (
            O => \N__33855\,
            I => \N__33808\
        );

    \I__5869\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33808\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__33851\,
            I => \N__33805\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__33850\,
            I => \N__33800\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__33849\,
            I => \N__33797\
        );

    \I__5865\ : Span4Mux_v
    port map (
            O => \N__33846\,
            I => \N__33792\
        );

    \I__5864\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33789\
        );

    \I__5863\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33786\
        );

    \I__5862\ : Span4Mux_s1_v
    port map (
            O => \N__33841\,
            I => \N__33777\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__33830\,
            I => \N__33777\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__33825\,
            I => \N__33777\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__33818\,
            I => \N__33777\
        );

    \I__5858\ : Span4Mux_h
    port map (
            O => \N__33815\,
            I => \N__33770\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__33808\,
            I => \N__33770\
        );

    \I__5856\ : Span4Mux_s3_h
    port map (
            O => \N__33805\,
            I => \N__33770\
        );

    \I__5855\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33759\
        );

    \I__5854\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33759\
        );

    \I__5853\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33759\
        );

    \I__5852\ : InMux
    port map (
            O => \N__33797\,
            I => \N__33759\
        );

    \I__5851\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33759\
        );

    \I__5850\ : InMux
    port map (
            O => \N__33795\,
            I => \N__33756\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__33792\,
            I => n2940
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__33789\,
            I => n2940
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__33786\,
            I => n2940
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__33777\,
            I => n2940
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__33770\,
            I => n2940
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__33759\,
            I => n2940
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__33756\,
            I => n2940
        );

    \I__5842\ : InMux
    port map (
            O => \N__33741\,
            I => n12941
        );

    \I__5841\ : InMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__5839\ : Span4Mux_v
    port map (
            O => \N__33732\,
            I => \N__33728\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__33731\,
            I => \N__33725\
        );

    \I__5837\ : Span4Mux_h
    port map (
            O => \N__33728\,
            I => \N__33722\
        );

    \I__5836\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33719\
        );

    \I__5835\ : Odrv4
    port map (
            O => \N__33722\,
            I => n15346
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__33719\,
            I => n15346
        );

    \I__5833\ : InMux
    port map (
            O => \N__33714\,
            I => \N__33710\
        );

    \I__5832\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33702\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__33710\,
            I => \N__33693\
        );

    \I__5830\ : InMux
    port map (
            O => \N__33709\,
            I => \N__33690\
        );

    \I__5829\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33683\
        );

    \I__5828\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33683\
        );

    \I__5827\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33683\
        );

    \I__5826\ : InMux
    port map (
            O => \N__33705\,
            I => \N__33680\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__33702\,
            I => \N__33677\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__33701\,
            I => \N__33673\
        );

    \I__5823\ : CascadeMux
    port map (
            O => \N__33700\,
            I => \N__33670\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__33699\,
            I => \N__33664\
        );

    \I__5821\ : CascadeMux
    port map (
            O => \N__33698\,
            I => \N__33658\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__33697\,
            I => \N__33652\
        );

    \I__5819\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33648\
        );

    \I__5818\ : Span4Mux_v
    port map (
            O => \N__33693\,
            I => \N__33642\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__33690\,
            I => \N__33639\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__33683\,
            I => \N__33636\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__33680\,
            I => \N__33633\
        );

    \I__5814\ : Span4Mux_s2_h
    port map (
            O => \N__33677\,
            I => \N__33630\
        );

    \I__5813\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33627\
        );

    \I__5812\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33616\
        );

    \I__5811\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33616\
        );

    \I__5810\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33616\
        );

    \I__5809\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33616\
        );

    \I__5808\ : InMux
    port map (
            O => \N__33667\,
            I => \N__33616\
        );

    \I__5807\ : InMux
    port map (
            O => \N__33664\,
            I => \N__33607\
        );

    \I__5806\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33607\
        );

    \I__5805\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33607\
        );

    \I__5804\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33607\
        );

    \I__5803\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33594\
        );

    \I__5802\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33594\
        );

    \I__5801\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33594\
        );

    \I__5800\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33594\
        );

    \I__5799\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33594\
        );

    \I__5798\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33594\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__33648\,
            I => \N__33591\
        );

    \I__5796\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33588\
        );

    \I__5795\ : InMux
    port map (
            O => \N__33646\,
            I => \N__33583\
        );

    \I__5794\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33583\
        );

    \I__5793\ : Span4Mux_h
    port map (
            O => \N__33642\,
            I => \N__33574\
        );

    \I__5792\ : Span4Mux_v
    port map (
            O => \N__33639\,
            I => \N__33574\
        );

    \I__5791\ : Span4Mux_s3_h
    port map (
            O => \N__33636\,
            I => \N__33574\
        );

    \I__5790\ : Span4Mux_s2_v
    port map (
            O => \N__33633\,
            I => \N__33574\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__33630\,
            I => n2841
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__33627\,
            I => n2841
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__33616\,
            I => n2841
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__33607\,
            I => n2841
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__33594\,
            I => n2841
        );

    \I__5784\ : Odrv12
    port map (
            O => \N__33591\,
            I => n2841
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__33588\,
            I => n2841
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__33583\,
            I => n2841
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__33574\,
            I => n2841
        );

    \I__5780\ : InMux
    port map (
            O => \N__33555\,
            I => n12942
        );

    \I__5779\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33548\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__33551\,
            I => \N__33545\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__33548\,
            I => \N__33542\
        );

    \I__5776\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33539\
        );

    \I__5775\ : Span4Mux_v
    port map (
            O => \N__33542\,
            I => \N__33536\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__33539\,
            I => \N__33533\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__33536\,
            I => n15310
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__33533\,
            I => n15310
        );

    \I__5771\ : InMux
    port map (
            O => \N__33528\,
            I => \N__33525\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__33525\,
            I => \N__33518\
        );

    \I__5769\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33507\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__33523\,
            I => \N__33499\
        );

    \I__5767\ : CascadeMux
    port map (
            O => \N__33522\,
            I => \N__33496\
        );

    \I__5766\ : CascadeMux
    port map (
            O => \N__33521\,
            I => \N__33493\
        );

    \I__5765\ : Span4Mux_h
    port map (
            O => \N__33518\,
            I => \N__33488\
        );

    \I__5764\ : InMux
    port map (
            O => \N__33517\,
            I => \N__33483\
        );

    \I__5763\ : InMux
    port map (
            O => \N__33516\,
            I => \N__33483\
        );

    \I__5762\ : CascadeMux
    port map (
            O => \N__33515\,
            I => \N__33480\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__33514\,
            I => \N__33477\
        );

    \I__5760\ : CascadeMux
    port map (
            O => \N__33513\,
            I => \N__33474\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__33512\,
            I => \N__33471\
        );

    \I__5758\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33465\
        );

    \I__5757\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33465\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__33507\,
            I => \N__33460\
        );

    \I__5755\ : CascadeMux
    port map (
            O => \N__33506\,
            I => \N__33457\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__33505\,
            I => \N__33453\
        );

    \I__5753\ : CascadeMux
    port map (
            O => \N__33504\,
            I => \N__33449\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__33503\,
            I => \N__33446\
        );

    \I__5751\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33432\
        );

    \I__5750\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33432\
        );

    \I__5749\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33432\
        );

    \I__5748\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33432\
        );

    \I__5747\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33432\
        );

    \I__5746\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33432\
        );

    \I__5745\ : Span4Mux_h
    port map (
            O => \N__33488\,
            I => \N__33427\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__33483\,
            I => \N__33427\
        );

    \I__5743\ : InMux
    port map (
            O => \N__33480\,
            I => \N__33416\
        );

    \I__5742\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33416\
        );

    \I__5741\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33416\
        );

    \I__5740\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33416\
        );

    \I__5739\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33416\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__33465\,
            I => \N__33413\
        );

    \I__5737\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33408\
        );

    \I__5736\ : InMux
    port map (
            O => \N__33463\,
            I => \N__33408\
        );

    \I__5735\ : Span4Mux_s3_v
    port map (
            O => \N__33460\,
            I => \N__33405\
        );

    \I__5734\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33400\
        );

    \I__5733\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33400\
        );

    \I__5732\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33389\
        );

    \I__5731\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33389\
        );

    \I__5730\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33389\
        );

    \I__5729\ : InMux
    port map (
            O => \N__33446\,
            I => \N__33389\
        );

    \I__5728\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33389\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__33432\,
            I => n2742
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__33427\,
            I => n2742
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__33416\,
            I => n2742
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__33413\,
            I => n2742
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__33408\,
            I => n2742
        );

    \I__5722\ : Odrv4
    port map (
            O => \N__33405\,
            I => n2742
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__33400\,
            I => n2742
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__33389\,
            I => n2742
        );

    \I__5719\ : InMux
    port map (
            O => \N__33372\,
            I => n12943
        );

    \I__5718\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33366\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33363\
        );

    \I__5716\ : Span4Mux_h
    port map (
            O => \N__33363\,
            I => \N__33359\
        );

    \I__5715\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33356\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__33359\,
            I => n15852
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__33356\,
            I => n15852
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__33351\,
            I => \N__33346\
        );

    \I__5711\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33336\
        );

    \I__5710\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33331\
        );

    \I__5709\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33325\
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__33345\,
            I => \N__33322\
        );

    \I__5707\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33318\
        );

    \I__5706\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33315\
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__33342\,
            I => \N__33311\
        );

    \I__5704\ : CascadeMux
    port map (
            O => \N__33341\,
            I => \N__33307\
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__33340\,
            I => \N__33304\
        );

    \I__5702\ : CascadeMux
    port map (
            O => \N__33339\,
            I => \N__33298\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__33336\,
            I => \N__33293\
        );

    \I__5700\ : InMux
    port map (
            O => \N__33335\,
            I => \N__33288\
        );

    \I__5699\ : InMux
    port map (
            O => \N__33334\,
            I => \N__33288\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__33331\,
            I => \N__33285\
        );

    \I__5697\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33282\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__33329\,
            I => \N__33279\
        );

    \I__5695\ : CascadeMux
    port map (
            O => \N__33328\,
            I => \N__33275\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__33325\,
            I => \N__33270\
        );

    \I__5693\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33265\
        );

    \I__5692\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33265\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__33318\,
            I => \N__33260\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__33315\,
            I => \N__33260\
        );

    \I__5689\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33253\
        );

    \I__5688\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33253\
        );

    \I__5687\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33253\
        );

    \I__5686\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33244\
        );

    \I__5685\ : InMux
    port map (
            O => \N__33304\,
            I => \N__33244\
        );

    \I__5684\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33244\
        );

    \I__5683\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33244\
        );

    \I__5682\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33235\
        );

    \I__5681\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33235\
        );

    \I__5680\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33235\
        );

    \I__5679\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33235\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__33293\,
            I => \N__33226\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__33288\,
            I => \N__33226\
        );

    \I__5676\ : Span4Mux_s3_h
    port map (
            O => \N__33285\,
            I => \N__33226\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33226\
        );

    \I__5674\ : InMux
    port map (
            O => \N__33279\,
            I => \N__33215\
        );

    \I__5673\ : InMux
    port map (
            O => \N__33278\,
            I => \N__33215\
        );

    \I__5672\ : InMux
    port map (
            O => \N__33275\,
            I => \N__33215\
        );

    \I__5671\ : InMux
    port map (
            O => \N__33274\,
            I => \N__33215\
        );

    \I__5670\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33215\
        );

    \I__5669\ : Odrv4
    port map (
            O => \N__33270\,
            I => n2643
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__33265\,
            I => n2643
        );

    \I__5667\ : Odrv4
    port map (
            O => \N__33260\,
            I => n2643
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__33253\,
            I => n2643
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__33244\,
            I => n2643
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__33235\,
            I => n2643
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__33226\,
            I => n2643
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__33215\,
            I => n2643
        );

    \I__5661\ : InMux
    port map (
            O => \N__33198\,
            I => n12944
        );

    \I__5660\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33192\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__5658\ : Span4Mux_h
    port map (
            O => \N__33189\,
            I => \N__33185\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__33188\,
            I => \N__33182\
        );

    \I__5656\ : Span4Mux_h
    port map (
            O => \N__33185\,
            I => \N__33179\
        );

    \I__5655\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33176\
        );

    \I__5654\ : Odrv4
    port map (
            O => \N__33179\,
            I => n15821
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__33176\,
            I => n15821
        );

    \I__5652\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33167\
        );

    \I__5651\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33160\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__33167\,
            I => \N__33152\
        );

    \I__5649\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33149\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__33165\,
            I => \N__33145\
        );

    \I__5647\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33140\
        );

    \I__5646\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33140\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__33160\,
            I => \N__33137\
        );

    \I__5644\ : CascadeMux
    port map (
            O => \N__33159\,
            I => \N__33132\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__33158\,
            I => \N__33128\
        );

    \I__5642\ : CascadeMux
    port map (
            O => \N__33157\,
            I => \N__33122\
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__33156\,
            I => \N__33115\
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__33155\,
            I => \N__33111\
        );

    \I__5639\ : Span4Mux_h
    port map (
            O => \N__33152\,
            I => \N__33105\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__33149\,
            I => \N__33105\
        );

    \I__5637\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33102\
        );

    \I__5636\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33099\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__33140\,
            I => \N__33096\
        );

    \I__5634\ : Span4Mux_s2_h
    port map (
            O => \N__33137\,
            I => \N__33092\
        );

    \I__5633\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33083\
        );

    \I__5632\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33083\
        );

    \I__5631\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33083\
        );

    \I__5630\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33083\
        );

    \I__5629\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33070\
        );

    \I__5628\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33070\
        );

    \I__5627\ : InMux
    port map (
            O => \N__33126\,
            I => \N__33070\
        );

    \I__5626\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33070\
        );

    \I__5625\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33070\
        );

    \I__5624\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33070\
        );

    \I__5623\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33065\
        );

    \I__5622\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33065\
        );

    \I__5621\ : InMux
    port map (
            O => \N__33118\,
            I => \N__33054\
        );

    \I__5620\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33054\
        );

    \I__5619\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33054\
        );

    \I__5618\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33054\
        );

    \I__5617\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33054\
        );

    \I__5616\ : Span4Mux_h
    port map (
            O => \N__33105\,
            I => \N__33045\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__33102\,
            I => \N__33045\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33045\
        );

    \I__5613\ : Span4Mux_h
    port map (
            O => \N__33096\,
            I => \N__33045\
        );

    \I__5612\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33042\
        );

    \I__5611\ : Odrv4
    port map (
            O => \N__33092\,
            I => n2544
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__33083\,
            I => n2544
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__33070\,
            I => n2544
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__33065\,
            I => n2544
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__33054\,
            I => n2544
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__33045\,
            I => n2544
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__33042\,
            I => n2544
        );

    \I__5604\ : InMux
    port map (
            O => \N__33027\,
            I => \bfn_7_24_0_\
        );

    \I__5603\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__33021\,
            I => \N__33017\
        );

    \I__5601\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33014\
        );

    \I__5600\ : Span4Mux_v
    port map (
            O => \N__33017\,
            I => \N__33011\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__33014\,
            I => \N__33008\
        );

    \I__5598\ : Span4Mux_h
    port map (
            O => \N__33011\,
            I => \N__33005\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__33008\,
            I => n15791
        );

    \I__5596\ : Odrv4
    port map (
            O => \N__33005\,
            I => n15791
        );

    \I__5595\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32994\
        );

    \I__5594\ : InMux
    port map (
            O => \N__32999\,
            I => \N__32991\
        );

    \I__5593\ : CascadeMux
    port map (
            O => \N__32998\,
            I => \N__32988\
        );

    \I__5592\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32981\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__32994\,
            I => \N__32978\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32973\
        );

    \I__5589\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32970\
        );

    \I__5588\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32967\
        );

    \I__5587\ : CascadeMux
    port map (
            O => \N__32986\,
            I => \N__32962\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__32985\,
            I => \N__32959\
        );

    \I__5585\ : CascadeMux
    port map (
            O => \N__32984\,
            I => \N__32955\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__32981\,
            I => \N__32947\
        );

    \I__5583\ : Span4Mux_s2_h
    port map (
            O => \N__32978\,
            I => \N__32947\
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__32977\,
            I => \N__32942\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__32976\,
            I => \N__32937\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__32973\,
            I => \N__32930\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__32970\,
            I => \N__32930\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__32967\,
            I => \N__32930\
        );

    \I__5577\ : InMux
    port map (
            O => \N__32966\,
            I => \N__32927\
        );

    \I__5576\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32914\
        );

    \I__5575\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32914\
        );

    \I__5574\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32914\
        );

    \I__5573\ : InMux
    port map (
            O => \N__32958\,
            I => \N__32914\
        );

    \I__5572\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32914\
        );

    \I__5571\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32914\
        );

    \I__5570\ : CascadeMux
    port map (
            O => \N__32953\,
            I => \N__32911\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__32952\,
            I => \N__32908\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__32947\,
            I => \N__32901\
        );

    \I__5567\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32898\
        );

    \I__5566\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32887\
        );

    \I__5565\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32887\
        );

    \I__5564\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32887\
        );

    \I__5563\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32887\
        );

    \I__5562\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32887\
        );

    \I__5561\ : Span4Mux_v
    port map (
            O => \N__32930\,
            I => \N__32882\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__32927\,
            I => \N__32882\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32879\
        );

    \I__5558\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32866\
        );

    \I__5557\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32866\
        );

    \I__5556\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32866\
        );

    \I__5555\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32866\
        );

    \I__5554\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32866\
        );

    \I__5553\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32866\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__32901\,
            I => n2445
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__32898\,
            I => n2445
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__32887\,
            I => n2445
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__32882\,
            I => n2445
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__32879\,
            I => n2445
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__32866\,
            I => n2445
        );

    \I__5546\ : InMux
    port map (
            O => \N__32853\,
            I => n12946
        );

    \I__5545\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32847\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__32847\,
            I => \N__32843\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__32846\,
            I => \N__32840\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__32843\,
            I => \N__32837\
        );

    \I__5541\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32834\
        );

    \I__5540\ : Odrv4
    port map (
            O => \N__32837\,
            I => n15765
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__32834\,
            I => n15765
        );

    \I__5538\ : InMux
    port map (
            O => \N__32829\,
            I => \N__32825\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__32828\,
            I => \N__32814\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__32825\,
            I => \N__32809\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__32824\,
            I => \N__32802\
        );

    \I__5534\ : CascadeMux
    port map (
            O => \N__32823\,
            I => \N__32799\
        );

    \I__5533\ : CascadeMux
    port map (
            O => \N__32822\,
            I => \N__32795\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__32821\,
            I => \N__32789\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__32820\,
            I => \N__32786\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__32819\,
            I => \N__32783\
        );

    \I__5529\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32779\
        );

    \I__5528\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32772\
        );

    \I__5527\ : InMux
    port map (
            O => \N__32814\,
            I => \N__32772\
        );

    \I__5526\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32772\
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__32812\,
            I => \N__32769\
        );

    \I__5524\ : Span12Mux_h
    port map (
            O => \N__32809\,
            I => \N__32765\
        );

    \I__5523\ : InMux
    port map (
            O => \N__32808\,
            I => \N__32762\
        );

    \I__5522\ : InMux
    port map (
            O => \N__32807\,
            I => \N__32753\
        );

    \I__5521\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32753\
        );

    \I__5520\ : InMux
    port map (
            O => \N__32805\,
            I => \N__32753\
        );

    \I__5519\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32753\
        );

    \I__5518\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32742\
        );

    \I__5517\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32742\
        );

    \I__5516\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32742\
        );

    \I__5515\ : InMux
    port map (
            O => \N__32794\,
            I => \N__32742\
        );

    \I__5514\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32742\
        );

    \I__5513\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32731\
        );

    \I__5512\ : InMux
    port map (
            O => \N__32789\,
            I => \N__32731\
        );

    \I__5511\ : InMux
    port map (
            O => \N__32786\,
            I => \N__32731\
        );

    \I__5510\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32731\
        );

    \I__5509\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32731\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__32779\,
            I => \N__32726\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32726\
        );

    \I__5506\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32721\
        );

    \I__5505\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32721\
        );

    \I__5504\ : Odrv12
    port map (
            O => \N__32765\,
            I => n2346
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__32762\,
            I => n2346
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__32753\,
            I => n2346
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__32742\,
            I => n2346
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__32731\,
            I => n2346
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__32726\,
            I => n2346
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__32721\,
            I => n2346
        );

    \I__5497\ : InMux
    port map (
            O => \N__32706\,
            I => n12947
        );

    \I__5496\ : InMux
    port map (
            O => \N__32703\,
            I => \N__32699\
        );

    \I__5495\ : CascadeMux
    port map (
            O => \N__32702\,
            I => \N__32696\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__32699\,
            I => \N__32693\
        );

    \I__5493\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32690\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__32693\,
            I => n15739
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__32690\,
            I => n15739
        );

    \I__5490\ : CascadeMux
    port map (
            O => \N__32685\,
            I => \N__32677\
        );

    \I__5489\ : CascadeMux
    port map (
            O => \N__32684\,
            I => \N__32673\
        );

    \I__5488\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32668\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__32682\,
            I => \N__32665\
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__32681\,
            I => \N__32661\
        );

    \I__5485\ : CascadeMux
    port map (
            O => \N__32680\,
            I => \N__32657\
        );

    \I__5484\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32647\
        );

    \I__5483\ : InMux
    port map (
            O => \N__32676\,
            I => \N__32647\
        );

    \I__5482\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32644\
        );

    \I__5481\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32641\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__32671\,
            I => \N__32638\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__32668\,
            I => \N__32632\
        );

    \I__5478\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32627\
        );

    \I__5477\ : InMux
    port map (
            O => \N__32664\,
            I => \N__32627\
        );

    \I__5476\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32618\
        );

    \I__5475\ : InMux
    port map (
            O => \N__32660\,
            I => \N__32618\
        );

    \I__5474\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32618\
        );

    \I__5473\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32618\
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__32655\,
            I => \N__32615\
        );

    \I__5471\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32608\
        );

    \I__5470\ : InMux
    port map (
            O => \N__32653\,
            I => \N__32608\
        );

    \I__5469\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32605\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32602\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__32644\,
            I => \N__32597\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32597\
        );

    \I__5465\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32594\
        );

    \I__5464\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32589\
        );

    \I__5463\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32589\
        );

    \I__5462\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32586\
        );

    \I__5461\ : Span4Mux_v
    port map (
            O => \N__32632\,
            I => \N__32581\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__32627\,
            I => \N__32581\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__32618\,
            I => \N__32578\
        );

    \I__5458\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32573\
        );

    \I__5457\ : InMux
    port map (
            O => \N__32614\,
            I => \N__32573\
        );

    \I__5456\ : InMux
    port map (
            O => \N__32613\,
            I => \N__32570\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__32608\,
            I => \N__32567\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__32605\,
            I => \N__32562\
        );

    \I__5453\ : Span4Mux_h
    port map (
            O => \N__32602\,
            I => \N__32562\
        );

    \I__5452\ : Span4Mux_v
    port map (
            O => \N__32597\,
            I => \N__32555\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__32594\,
            I => \N__32555\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32555\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__32586\,
            I => n2247
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__32581\,
            I => n2247
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__32578\,
            I => n2247
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__32573\,
            I => n2247
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__32570\,
            I => n2247
        );

    \I__5444\ : Odrv4
    port map (
            O => \N__32567\,
            I => n2247
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__32562\,
            I => n2247
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__32555\,
            I => n2247
        );

    \I__5441\ : InMux
    port map (
            O => \N__32538\,
            I => n12948
        );

    \I__5440\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32532\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32529\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__32529\,
            I => n2284
        );

    \I__5437\ : CascadeMux
    port map (
            O => \N__32526\,
            I => \N__32523\
        );

    \I__5436\ : InMux
    port map (
            O => \N__32523\,
            I => \N__32519\
        );

    \I__5435\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32516\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__32519\,
            I => n2217
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__32516\,
            I => n2217
        );

    \I__5432\ : CascadeMux
    port map (
            O => \N__32511\,
            I => \N__32508\
        );

    \I__5431\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32504\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__32507\,
            I => \N__32501\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32497\
        );

    \I__5428\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32494\
        );

    \I__5427\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32491\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__32497\,
            I => \N__32488\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N__32485\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__32491\,
            I => \N__32482\
        );

    \I__5423\ : Span4Mux_h
    port map (
            O => \N__32488\,
            I => \N__32479\
        );

    \I__5422\ : Span4Mux_v
    port map (
            O => \N__32485\,
            I => \N__32474\
        );

    \I__5421\ : Span4Mux_v
    port map (
            O => \N__32482\,
            I => \N__32474\
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__32479\,
            I => n2316
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__32474\,
            I => n2316
        );

    \I__5418\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32466\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__32466\,
            I => \N__32463\
        );

    \I__5416\ : Odrv12
    port map (
            O => \N__32463\,
            I => n2100
        );

    \I__5415\ : CascadeMux
    port map (
            O => \N__32460\,
            I => \N__32457\
        );

    \I__5414\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32454\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__32454\,
            I => \N__32450\
        );

    \I__5412\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32446\
        );

    \I__5411\ : Span12Mux_v
    port map (
            O => \N__32450\,
            I => \N__32443\
        );

    \I__5410\ : InMux
    port map (
            O => \N__32449\,
            I => \N__32440\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__32446\,
            I => n2132
        );

    \I__5408\ : Odrv12
    port map (
            O => \N__32443\,
            I => n2132
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__32440\,
            I => n2132
        );

    \I__5406\ : InMux
    port map (
            O => \N__32433\,
            I => \N__32429\
        );

    \I__5405\ : InMux
    port map (
            O => \N__32432\,
            I => \N__32426\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__32429\,
            I => \N__32420\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__32426\,
            I => \N__32420\
        );

    \I__5402\ : InMux
    port map (
            O => \N__32425\,
            I => \N__32417\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__32420\,
            I => \N__32414\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__32417\,
            I => \N__32411\
        );

    \I__5399\ : Span4Mux_h
    port map (
            O => \N__32414\,
            I => \N__32408\
        );

    \I__5398\ : Span12Mux_s6_h
    port map (
            O => \N__32411\,
            I => \N__32405\
        );

    \I__5397\ : Span4Mux_v
    port map (
            O => \N__32408\,
            I => \N__32402\
        );

    \I__5396\ : Odrv12
    port map (
            O => \N__32405\,
            I => n315
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__32402\,
            I => n315
        );

    \I__5394\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32394\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__32394\,
            I => n15484
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__32391\,
            I => \N__32387\
        );

    \I__5391\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32384\
        );

    \I__5390\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32381\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__32384\,
            I => n12034
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__32381\,
            I => n12034
        );

    \I__5387\ : InMux
    port map (
            O => \N__32376\,
            I => \bfn_7_23_0_\
        );

    \I__5386\ : InMux
    port map (
            O => \N__32373\,
            I => n12938
        );

    \I__5385\ : InMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__32367\,
            I => \N__32363\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__32366\,
            I => \N__32360\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__32363\,
            I => \N__32357\
        );

    \I__5381\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32354\
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__32357\,
            I => n15445
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__32354\,
            I => n15445
        );

    \I__5378\ : InMux
    port map (
            O => \N__32349\,
            I => n12939
        );

    \I__5377\ : InMux
    port map (
            O => \N__32346\,
            I => \N__32343\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32340\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__32340\,
            I => \N__32337\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__32337\,
            I => \N__32333\
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__32336\,
            I => \N__32330\
        );

    \I__5372\ : Span4Mux_h
    port map (
            O => \N__32333\,
            I => \N__32327\
        );

    \I__5371\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32324\
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__32327\,
            I => n15412
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__32324\,
            I => n15412
        );

    \I__5368\ : InMux
    port map (
            O => \N__32319\,
            I => n12940
        );

    \I__5367\ : InMux
    port map (
            O => \N__32316\,
            I => \N__32313\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__32313\,
            I => \N__32310\
        );

    \I__5365\ : Span4Mux_v
    port map (
            O => \N__32310\,
            I => \N__32307\
        );

    \I__5364\ : Span4Mux_v
    port map (
            O => \N__32307\,
            I => \N__32303\
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__32306\,
            I => \N__32300\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__32303\,
            I => \N__32297\
        );

    \I__5361\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32294\
        );

    \I__5360\ : Odrv4
    port map (
            O => \N__32297\,
            I => n15378
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__32294\,
            I => n15378
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__32289\,
            I => \N__32286\
        );

    \I__5357\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32282\
        );

    \I__5356\ : InMux
    port map (
            O => \N__32285\,
            I => \N__32279\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__32282\,
            I => \N__32276\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__32279\,
            I => \N__32273\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__32276\,
            I => \N__32270\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__32273\,
            I => n2127
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__32270\,
            I => n2127
        );

    \I__5350\ : CascadeMux
    port map (
            O => \N__32265\,
            I => \N__32262\
        );

    \I__5349\ : InMux
    port map (
            O => \N__32262\,
            I => \N__32259\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__32259\,
            I => \N__32256\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__32256\,
            I => \N__32253\
        );

    \I__5346\ : Odrv4
    port map (
            O => \N__32253\,
            I => n2194
        );

    \I__5345\ : InMux
    port map (
            O => \N__32250\,
            I => \N__32246\
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__32249\,
            I => \N__32243\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__32246\,
            I => \N__32240\
        );

    \I__5342\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32237\
        );

    \I__5341\ : Span4Mux_v
    port map (
            O => \N__32240\,
            I => \N__32231\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__32237\,
            I => \N__32231\
        );

    \I__5339\ : InMux
    port map (
            O => \N__32236\,
            I => \N__32228\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__32231\,
            I => n2226
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__32228\,
            I => n2226
        );

    \I__5336\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32220\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__32220\,
            I => \N__32217\
        );

    \I__5334\ : Odrv12
    port map (
            O => \N__32217\,
            I => n2101
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__32214\,
            I => \N__32211\
        );

    \I__5332\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32208\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32204\
        );

    \I__5330\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32201\
        );

    \I__5329\ : Span4Mux_h
    port map (
            O => \N__32204\,
            I => \N__32198\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__32201\,
            I => n2133
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__32198\,
            I => n2133
        );

    \I__5326\ : CascadeMux
    port map (
            O => \N__32193\,
            I => \n2133_cascade_\
        );

    \I__5325\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32187\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__32187\,
            I => n11892
        );

    \I__5323\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32179\
        );

    \I__5322\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32174\
        );

    \I__5321\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32174\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__32179\,
            I => \N__32171\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__32174\,
            I => \N__32168\
        );

    \I__5318\ : Span4Mux_v
    port map (
            O => \N__32171\,
            I => \N__32165\
        );

    \I__5317\ : Span4Mux_h
    port map (
            O => \N__32168\,
            I => \N__32162\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__32165\,
            I => n307
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__32162\,
            I => n307
        );

    \I__5314\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32154\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__32154\,
            I => \N__32151\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__5311\ : Odrv4
    port map (
            O => \N__32148\,
            I => n2201
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__32145\,
            I => \N__32142\
        );

    \I__5309\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__32139\,
            I => \N__32135\
        );

    \I__5307\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32132\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__32135\,
            I => \N__32129\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__32132\,
            I => n2233
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__32129\,
            I => n2233
        );

    \I__5303\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32120\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__32123\,
            I => \N__32117\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__32120\,
            I => \N__32113\
        );

    \I__5300\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32110\
        );

    \I__5299\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32107\
        );

    \I__5298\ : Odrv12
    port map (
            O => \N__32113\,
            I => n2231
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__32110\,
            I => n2231
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__32107\,
            I => n2231
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__32100\,
            I => \n2233_cascade_\
        );

    \I__5294\ : CascadeMux
    port map (
            O => \N__32097\,
            I => \N__32093\
        );

    \I__5293\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32089\
        );

    \I__5292\ : InMux
    port map (
            O => \N__32093\,
            I => \N__32086\
        );

    \I__5291\ : InMux
    port map (
            O => \N__32092\,
            I => \N__32083\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__32089\,
            I => n2232
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__32086\,
            I => n2232
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__32083\,
            I => n2232
        );

    \I__5287\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32073\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__32073\,
            I => n11950
        );

    \I__5285\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32067\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__32067\,
            I => \N__32064\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__32064\,
            I => n2086
        );

    \I__5282\ : InMux
    port map (
            O => \N__32061\,
            I => \N__32058\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__32058\,
            I => \N__32054\
        );

    \I__5280\ : InMux
    port map (
            O => \N__32057\,
            I => \N__32050\
        );

    \I__5279\ : Span4Mux_h
    port map (
            O => \N__32054\,
            I => \N__32047\
        );

    \I__5278\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32044\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__32050\,
            I => n2118
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__32047\,
            I => n2118
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__32044\,
            I => n2118
        );

    \I__5274\ : InMux
    port map (
            O => \N__32037\,
            I => \N__32033\
        );

    \I__5273\ : InMux
    port map (
            O => \N__32036\,
            I => \N__32030\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__32033\,
            I => \N__32027\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__32024\
        );

    \I__5270\ : Span4Mux_v
    port map (
            O => \N__32027\,
            I => \N__32020\
        );

    \I__5269\ : Span12Mux_s6_h
    port map (
            O => \N__32024\,
            I => \N__32017\
        );

    \I__5268\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32014\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__32020\,
            I => n308
        );

    \I__5266\ : Odrv12
    port map (
            O => \N__32017\,
            I => n308
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__32014\,
            I => n308
        );

    \I__5264\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__32004\,
            I => \N__32001\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__32001\,
            I => n2098
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__31998\,
            I => \N__31995\
        );

    \I__5260\ : InMux
    port map (
            O => \N__31995\,
            I => \N__31992\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__31992\,
            I => \N__31988\
        );

    \I__5258\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31985\
        );

    \I__5257\ : Span4Mux_h
    port map (
            O => \N__31988\,
            I => \N__31982\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__31985\,
            I => n2130
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__31982\,
            I => n2130
        );

    \I__5254\ : CascadeMux
    port map (
            O => \N__31977\,
            I => \N__31974\
        );

    \I__5253\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31971\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__31971\,
            I => \N__31966\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__31970\,
            I => \N__31963\
        );

    \I__5250\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31960\
        );

    \I__5249\ : Span4Mux_v
    port map (
            O => \N__31966\,
            I => \N__31957\
        );

    \I__5248\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31954\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__31960\,
            I => \N__31951\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__31957\,
            I => n2131
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__31954\,
            I => n2131
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__31951\,
            I => n2131
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__31944\,
            I => \N__31941\
        );

    \I__5242\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31937\
        );

    \I__5241\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31933\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__31937\,
            I => \N__31930\
        );

    \I__5239\ : CascadeMux
    port map (
            O => \N__31936\,
            I => \N__31927\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__31933\,
            I => \N__31924\
        );

    \I__5237\ : Span4Mux_v
    port map (
            O => \N__31930\,
            I => \N__31921\
        );

    \I__5236\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31918\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__31924\,
            I => \N__31915\
        );

    \I__5234\ : Odrv4
    port map (
            O => \N__31921\,
            I => n2129
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__31918\,
            I => n2129
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__31915\,
            I => n2129
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__31908\,
            I => \n2130_cascade_\
        );

    \I__5230\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31900\
        );

    \I__5229\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31897\
        );

    \I__5228\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31894\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__31900\,
            I => n2119
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__31897\,
            I => n2119
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__31894\,
            I => n2119
        );

    \I__5224\ : CascadeMux
    port map (
            O => \N__31887\,
            I => \n13775_cascade_\
        );

    \I__5223\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31881\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__31881\,
            I => n14398
        );

    \I__5221\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31875\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__31875\,
            I => \N__31872\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__31872\,
            I => n2090
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__31869\,
            I => \N__31866\
        );

    \I__5217\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31863\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31859\
        );

    \I__5215\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31856\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__31859\,
            I => \N__31853\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__31856\,
            I => n2122
        );

    \I__5212\ : Odrv4
    port map (
            O => \N__31853\,
            I => n2122
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__31848\,
            I => \N__31844\
        );

    \I__5210\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31840\
        );

    \I__5209\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31837\
        );

    \I__5208\ : InMux
    port map (
            O => \N__31843\,
            I => \N__31834\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__31840\,
            I => n2125
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__31837\,
            I => n2125
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__31834\,
            I => n2125
        );

    \I__5204\ : CascadeMux
    port map (
            O => \N__31827\,
            I => \n2122_cascade_\
        );

    \I__5203\ : CascadeMux
    port map (
            O => \N__31824\,
            I => \N__31819\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__31823\,
            I => \N__31816\
        );

    \I__5201\ : InMux
    port map (
            O => \N__31822\,
            I => \N__31813\
        );

    \I__5200\ : InMux
    port map (
            O => \N__31819\,
            I => \N__31810\
        );

    \I__5199\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31807\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__31813\,
            I => \N__31804\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__31810\,
            I => n2128
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__31807\,
            I => n2128
        );

    \I__5195\ : Odrv4
    port map (
            O => \N__31804\,
            I => n2128
        );

    \I__5194\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31794\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__31794\,
            I => \N__31789\
        );

    \I__5192\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31786\
        );

    \I__5191\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31783\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__31789\,
            I => n2120
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__31786\,
            I => n2120
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__31783\,
            I => n2120
        );

    \I__5187\ : CascadeMux
    port map (
            O => \N__31776\,
            I => \n14386_cascade_\
        );

    \I__5186\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31770\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__31770\,
            I => n14384
        );

    \I__5184\ : InMux
    port map (
            O => \N__31767\,
            I => \N__31764\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__31764\,
            I => n14392
        );

    \I__5182\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__31758\,
            I => \N__31755\
        );

    \I__5180\ : Odrv4
    port map (
            O => \N__31755\,
            I => n2089
        );

    \I__5179\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31748\
        );

    \I__5178\ : CascadeMux
    port map (
            O => \N__31751\,
            I => \N__31745\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__31748\,
            I => \N__31742\
        );

    \I__5176\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31738\
        );

    \I__5175\ : Span4Mux_h
    port map (
            O => \N__31742\,
            I => \N__31735\
        );

    \I__5174\ : InMux
    port map (
            O => \N__31741\,
            I => \N__31732\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__31738\,
            I => n2121
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__31735\,
            I => n2121
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__31732\,
            I => n2121
        );

    \I__5170\ : InMux
    port map (
            O => \N__31725\,
            I => n12639
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__31722\,
            I => \N__31719\
        );

    \I__5168\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__31716\,
            I => n2085
        );

    \I__5166\ : InMux
    port map (
            O => \N__31713\,
            I => \bfn_7_19_0_\
        );

    \I__5165\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__31707\,
            I => n2084
        );

    \I__5163\ : InMux
    port map (
            O => \N__31704\,
            I => n12641
        );

    \I__5162\ : InMux
    port map (
            O => \N__31701\,
            I => n12642
        );

    \I__5161\ : CascadeMux
    port map (
            O => \N__31698\,
            I => \N__31695\
        );

    \I__5160\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__31692\,
            I => \N__31688\
        );

    \I__5158\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31685\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__31688\,
            I => n2115
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__31685\,
            I => n2115
        );

    \I__5155\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31677\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__31677\,
            I => \N__31674\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__31674\,
            I => n2095
        );

    \I__5152\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31667\
        );

    \I__5151\ : CascadeMux
    port map (
            O => \N__31670\,
            I => \N__31664\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__31667\,
            I => \N__31660\
        );

    \I__5149\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31657\
        );

    \I__5148\ : InMux
    port map (
            O => \N__31663\,
            I => \N__31654\
        );

    \I__5147\ : Odrv4
    port map (
            O => \N__31660\,
            I => n2123
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__31657\,
            I => n2123
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__31654\,
            I => n2123
        );

    \I__5144\ : CascadeMux
    port map (
            O => \N__31647\,
            I => \n2127_cascade_\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__31644\,
            I => \N__31641\
        );

    \I__5142\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31637\
        );

    \I__5141\ : InMux
    port map (
            O => \N__31640\,
            I => \N__31634\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__31637\,
            I => n2126
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__31634\,
            I => n2126
        );

    \I__5138\ : CascadeMux
    port map (
            O => \N__31629\,
            I => \N__31624\
        );

    \I__5137\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31621\
        );

    \I__5136\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31618\
        );

    \I__5135\ : InMux
    port map (
            O => \N__31624\,
            I => \N__31615\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__31621\,
            I => n2018
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__31618\,
            I => n2018
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__31615\,
            I => n2018
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__31608\,
            I => \N__31605\
        );

    \I__5130\ : InMux
    port map (
            O => \N__31605\,
            I => \N__31602\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__31602\,
            I => n2092
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__31599\,
            I => \N__31596\
        );

    \I__5127\ : InMux
    port map (
            O => \N__31596\,
            I => \N__31592\
        );

    \I__5126\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31589\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__31592\,
            I => \N__31586\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__31589\,
            I => \N__31580\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__31586\,
            I => \N__31580\
        );

    \I__5122\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31577\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__31580\,
            I => n2124
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__31577\,
            I => n2124
        );

    \I__5119\ : InMux
    port map (
            O => \N__31572\,
            I => n12630
        );

    \I__5118\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31566\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__31566\,
            I => n2094
        );

    \I__5116\ : InMux
    port map (
            O => \N__31563\,
            I => n12631
        );

    \I__5115\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31557\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__31557\,
            I => n2093
        );

    \I__5113\ : InMux
    port map (
            O => \N__31554\,
            I => \bfn_7_18_0_\
        );

    \I__5112\ : InMux
    port map (
            O => \N__31551\,
            I => n12633
        );

    \I__5111\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31545\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__31545\,
            I => n2091
        );

    \I__5109\ : InMux
    port map (
            O => \N__31542\,
            I => n12634
        );

    \I__5108\ : InMux
    port map (
            O => \N__31539\,
            I => n12635
        );

    \I__5107\ : InMux
    port map (
            O => \N__31536\,
            I => n12636
        );

    \I__5106\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31530\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__31530\,
            I => n2088
        );

    \I__5104\ : InMux
    port map (
            O => \N__31527\,
            I => n12637
        );

    \I__5103\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31521\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__31521\,
            I => n2087
        );

    \I__5101\ : InMux
    port map (
            O => \N__31518\,
            I => n12638
        );

    \I__5100\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__31512\,
            I => n14258
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__31509\,
            I => \n14260_cascade_\
        );

    \I__5097\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31503\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__31503\,
            I => n14262
        );

    \I__5095\ : InMux
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__31497\,
            I => \N__31493\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__31496\,
            I => \N__31490\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__31493\,
            I => \N__31486\
        );

    \I__5091\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31483\
        );

    \I__5090\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31480\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__31486\,
            I => n3021
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__31483\,
            I => n3021
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__31480\,
            I => n3021
        );

    \I__5086\ : CascadeMux
    port map (
            O => \N__31473\,
            I => \N__31470\
        );

    \I__5085\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31467\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__31467\,
            I => \N__31464\
        );

    \I__5083\ : Span4Mux_s2_v
    port map (
            O => \N__31464\,
            I => \N__31461\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__31461\,
            I => n3088
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__31458\,
            I => \N__31454\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__31457\,
            I => \N__31451\
        );

    \I__5079\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31448\
        );

    \I__5078\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31445\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__31448\,
            I => \N__31442\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__31445\,
            I => \N__31436\
        );

    \I__5075\ : Span12Mux_s5_h
    port map (
            O => \N__31442\,
            I => \N__31436\
        );

    \I__5074\ : InMux
    port map (
            O => \N__31441\,
            I => \N__31433\
        );

    \I__5073\ : Odrv12
    port map (
            O => \N__31436\,
            I => n3120
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__31433\,
            I => n3120
        );

    \I__5071\ : InMux
    port map (
            O => \N__31428\,
            I => \bfn_7_17_0_\
        );

    \I__5070\ : InMux
    port map (
            O => \N__31425\,
            I => n12625
        );

    \I__5069\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31419\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__31419\,
            I => n2099
        );

    \I__5067\ : InMux
    port map (
            O => \N__31416\,
            I => n12626
        );

    \I__5066\ : InMux
    port map (
            O => \N__31413\,
            I => n12627
        );

    \I__5065\ : InMux
    port map (
            O => \N__31410\,
            I => \N__31407\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__31407\,
            I => n2097
        );

    \I__5063\ : InMux
    port map (
            O => \N__31404\,
            I => n12628
        );

    \I__5062\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__31398\,
            I => n2096
        );

    \I__5060\ : InMux
    port map (
            O => \N__31395\,
            I => n12629
        );

    \I__5059\ : CascadeMux
    port map (
            O => \N__31392\,
            I => \n14250_cascade_\
        );

    \I__5058\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31386\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31381\
        );

    \I__5056\ : InMux
    port map (
            O => \N__31385\,
            I => \N__31378\
        );

    \I__5055\ : InMux
    port map (
            O => \N__31384\,
            I => \N__31375\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__31381\,
            I => \N__31370\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__31378\,
            I => \N__31370\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31367\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__31370\,
            I => n3026
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__31367\,
            I => n3026
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__31362\,
            I => \N__31359\
        );

    \I__5048\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31356\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__31356\,
            I => \N__31353\
        );

    \I__5046\ : Span4Mux_s2_v
    port map (
            O => \N__31353\,
            I => \N__31350\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__31350\,
            I => n3093
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__31347\,
            I => \N__31344\
        );

    \I__5043\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31341\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__31338\,
            I => \N__31335\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__31335\,
            I => n59
        );

    \I__5039\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31329\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__31329\,
            I => n14252
        );

    \I__5037\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__31323\,
            I => n5_adj_703
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__31320\,
            I => \n14254_cascade_\
        );

    \I__5034\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31314\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__5032\ : Odrv4
    port map (
            O => \N__31311\,
            I => n11926
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__31308\,
            I => \n14256_cascade_\
        );

    \I__5030\ : InMux
    port map (
            O => \N__31305\,
            I => \N__31302\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__31302\,
            I => n7_adj_708
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__31299\,
            I => \n14264_cascade_\
        );

    \I__5027\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31293\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__31293\,
            I => \N__31290\
        );

    \I__5025\ : Span4Mux_v
    port map (
            O => \N__31290\,
            I => \N__31287\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__31287\,
            I => n14266
        );

    \I__5023\ : InMux
    port map (
            O => \N__31284\,
            I => \N__31281\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31278\
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__31278\,
            I => n3101
        );

    \I__5020\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31272\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__31269\,
            I => \N__31266\
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__31266\,
            I => n3200
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__31263\,
            I => \n3133_cascade_\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__31260\,
            I => \n3232_cascade_\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__31257\,
            I => \n25_adj_712_cascade_\
        );

    \I__5013\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31251\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__31251\,
            I => n37_adj_715
        );

    \I__5011\ : InMux
    port map (
            O => \N__31248\,
            I => \N__31245\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__31245\,
            I => n14234
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__31242\,
            I => \n14238_cascade_\
        );

    \I__5008\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31236\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__5006\ : Odrv12
    port map (
            O => \N__31233\,
            I => n14248
        );

    \I__5005\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31224\
        );

    \I__5003\ : Span4Mux_v
    port map (
            O => \N__31224\,
            I => \N__31221\
        );

    \I__5002\ : Span4Mux_h
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__31218\,
            I => n3201
        );

    \I__5000\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31212\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__4998\ : Odrv4
    port map (
            O => \N__31209\,
            I => n11861
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__31206\,
            I => \n3233_cascade_\
        );

    \I__4996\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31196\
        );

    \I__4995\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31196\
        );

    \I__4994\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31193\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__31196\,
            I => \N__31190\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__31193\,
            I => \N__31187\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__31190\,
            I => \N__31184\
        );

    \I__4990\ : Odrv12
    port map (
            O => \N__31187\,
            I => n3111
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__31184\,
            I => n3111
        );

    \I__4988\ : CascadeMux
    port map (
            O => \N__31179\,
            I => \N__31176\
        );

    \I__4987\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31173\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__31173\,
            I => n3178
        );

    \I__4985\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31166\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__31169\,
            I => \N__31163\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__31166\,
            I => \N__31160\
        );

    \I__4982\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31157\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__31160\,
            I => n3023
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__31157\,
            I => n3023
        );

    \I__4979\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__31149\,
            I => \N__31146\
        );

    \I__4977\ : Span4Mux_h
    port map (
            O => \N__31146\,
            I => \N__31143\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__31143\,
            I => n3090
        );

    \I__4975\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31135\
        );

    \I__4974\ : InMux
    port map (
            O => \N__31139\,
            I => \N__31132\
        );

    \I__4973\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31129\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__31135\,
            I => \N__31126\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__31132\,
            I => \N__31121\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__31129\,
            I => \N__31121\
        );

    \I__4969\ : Span4Mux_s1_v
    port map (
            O => \N__31126\,
            I => \N__31118\
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__31121\,
            I => n3122
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__31118\,
            I => n3122
        );

    \I__4966\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__31110\,
            I => \N__31107\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__31107\,
            I => n3181
        );

    \I__4963\ : CascadeMux
    port map (
            O => \N__31104\,
            I => \N__31101\
        );

    \I__4962\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__31098\,
            I => \N__31095\
        );

    \I__4960\ : Span4Mux_v
    port map (
            O => \N__31095\,
            I => \N__31092\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__31092\,
            I => n3199
        );

    \I__4958\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__31086\,
            I => \N__31083\
        );

    \I__4956\ : Span4Mux_v
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__31080\,
            I => n3198
        );

    \I__4954\ : InMux
    port map (
            O => \N__31077\,
            I => \N__31073\
        );

    \I__4953\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31069\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31066\
        );

    \I__4951\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31063\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__31069\,
            I => \N__31060\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__31066\,
            I => \N__31055\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__31063\,
            I => \N__31055\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__31060\,
            I => n3115
        );

    \I__4946\ : Odrv4
    port map (
            O => \N__31055\,
            I => n3115
        );

    \I__4945\ : InMux
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__31047\,
            I => \N__31043\
        );

    \I__4943\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31039\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__31043\,
            I => \N__31036\
        );

    \I__4941\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31033\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__31039\,
            I => n3114
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__31036\,
            I => n3114
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__31033\,
            I => n3114
        );

    \I__4937\ : InMux
    port map (
            O => \N__31026\,
            I => \N__31023\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__31023\,
            I => \N__31020\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__31020\,
            I => n14204
        );

    \I__4934\ : InMux
    port map (
            O => \N__31017\,
            I => \N__31014\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__31014\,
            I => n14210
        );

    \I__4932\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__31008\,
            I => n3175
        );

    \I__4930\ : CascadeMux
    port map (
            O => \N__31005\,
            I => \N__31001\
        );

    \I__4929\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30998\
        );

    \I__4928\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30995\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__30998\,
            I => \N__30992\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__30995\,
            I => \N__30989\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__30992\,
            I => \N__30985\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__30989\,
            I => \N__30982\
        );

    \I__4923\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30979\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__30985\,
            I => n3121
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__30982\,
            I => n3121
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__30979\,
            I => n3121
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__4918\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__30966\,
            I => n3188
        );

    \I__4916\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30960\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__30960\,
            I => n3191
        );

    \I__4914\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30954\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__30954\,
            I => \N__30950\
        );

    \I__4912\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30947\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__30950\,
            I => \N__30943\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__30947\,
            I => \N__30940\
        );

    \I__4909\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30937\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__30943\,
            I => n3124
        );

    \I__4907\ : Odrv12
    port map (
            O => \N__30940\,
            I => n3124
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__30937\,
            I => n3124
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__30930\,
            I => \N__30927\
        );

    \I__4904\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30924\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__30924\,
            I => n3179
        );

    \I__4902\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30916\
        );

    \I__4901\ : CascadeMux
    port map (
            O => \N__30920\,
            I => \N__30913\
        );

    \I__4900\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30910\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__30916\,
            I => \N__30907\
        );

    \I__4898\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30904\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__30910\,
            I => n3113
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__30907\,
            I => n3113
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__30904\,
            I => n3113
        );

    \I__4894\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__30894\,
            I => \N__30889\
        );

    \I__4892\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30886\
        );

    \I__4891\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30883\
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__30889\,
            I => n3108
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__30886\,
            I => n3108
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__30883\,
            I => n3108
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__30876\,
            I => \n14216_cascade_\
        );

    \I__4886\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30869\
        );

    \I__4885\ : InMux
    port map (
            O => \N__30872\,
            I => \N__30866\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__30869\,
            I => \N__30861\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30861\
        );

    \I__4882\ : Span4Mux_h
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__30858\,
            I => n3105
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__30855\,
            I => \n14222_cascade_\
        );

    \I__4879\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30849\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__30849\,
            I => \N__30844\
        );

    \I__4877\ : InMux
    port map (
            O => \N__30848\,
            I => \N__30841\
        );

    \I__4876\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30838\
        );

    \I__4875\ : Span4Mux_v
    port map (
            O => \N__30844\,
            I => \N__30835\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__30841\,
            I => \N__30830\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30830\
        );

    \I__4872\ : Span4Mux_v
    port map (
            O => \N__30835\,
            I => \N__30827\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__30830\,
            I => \N__30824\
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__30827\,
            I => n3106
        );

    \I__4869\ : Odrv4
    port map (
            O => \N__30824\,
            I => n3106
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__30819\,
            I => \n3138_cascade_\
        );

    \I__4867\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30811\
        );

    \I__4866\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30806\
        );

    \I__4865\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30806\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__30811\,
            I => \N__30801\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__30806\,
            I => \N__30801\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__30798\,
            I => n3107
        );

    \I__4860\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30792\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__30792\,
            I => n3174
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__30789\,
            I => \n3214_cascade_\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__30786\,
            I => \N__30783\
        );

    \I__4856\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30780\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__30780\,
            I => n3190
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__30777\,
            I => \n3222_cascade_\
        );

    \I__4853\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30771\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__30771\,
            I => n27_adj_713
        );

    \I__4851\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30765\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__30765\,
            I => n3183
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__30762\,
            I => \N__30759\
        );

    \I__4848\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30756\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30752\
        );

    \I__4846\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30749\
        );

    \I__4845\ : Span4Mux_v
    port map (
            O => \N__30752\,
            I => \N__30745\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__30749\,
            I => \N__30742\
        );

    \I__4843\ : InMux
    port map (
            O => \N__30748\,
            I => \N__30739\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__30745\,
            I => n3116
        );

    \I__4841\ : Odrv12
    port map (
            O => \N__30742\,
            I => n3116
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__30739\,
            I => n3116
        );

    \I__4839\ : InMux
    port map (
            O => \N__30732\,
            I => \N__30729\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__30729\,
            I => n14794
        );

    \I__4837\ : InMux
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__30723\,
            I => n14800
        );

    \I__4835\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30717\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__30717\,
            I => \N__30714\
        );

    \I__4833\ : Odrv12
    port map (
            O => \N__30714\,
            I => n2891
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__30711\,
            I => \N__30707\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__30710\,
            I => \N__30704\
        );

    \I__4830\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30701\
        );

    \I__4829\ : InMux
    port map (
            O => \N__30704\,
            I => \N__30698\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__30701\,
            I => \N__30694\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__30698\,
            I => \N__30691\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__30697\,
            I => \N__30688\
        );

    \I__4825\ : Span4Mux_v
    port map (
            O => \N__30694\,
            I => \N__30685\
        );

    \I__4824\ : Span4Mux_v
    port map (
            O => \N__30691\,
            I => \N__30682\
        );

    \I__4823\ : InMux
    port map (
            O => \N__30688\,
            I => \N__30679\
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__30685\,
            I => n2824
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__30682\,
            I => n2824
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__30679\,
            I => n2824
        );

    \I__4819\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30668\
        );

    \I__4818\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__30668\,
            I => \N__30661\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30658\
        );

    \I__4815\ : InMux
    port map (
            O => \N__30664\,
            I => \N__30655\
        );

    \I__4814\ : Span4Mux_s3_v
    port map (
            O => \N__30661\,
            I => \N__30652\
        );

    \I__4813\ : Span12Mux_s5_v
    port map (
            O => \N__30658\,
            I => \N__30649\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30646\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__30652\,
            I => n2923
        );

    \I__4810\ : Odrv12
    port map (
            O => \N__30649\,
            I => n2923
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__30646\,
            I => n2923
        );

    \I__4808\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__30636\,
            I => n3187
        );

    \I__4806\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__30630\,
            I => n3189
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__30627\,
            I => \n3221_cascade_\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__30624\,
            I => \n14268_cascade_\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__30621\,
            I => \n14806_cascade_\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__30618\,
            I => \n3237_cascade_\
        );

    \I__4800\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30612\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__30612\,
            I => n14228
        );

    \I__4798\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30606\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__30606\,
            I => n14270
        );

    \I__4796\ : InMux
    port map (
            O => \N__30603\,
            I => \N__30600\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__30600\,
            I => n14272
        );

    \I__4794\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30594\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__30591\,
            I => n3173
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__30588\,
            I => \N__30585\
        );

    \I__4790\ : InMux
    port map (
            O => \N__30585\,
            I => \N__30582\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__30582\,
            I => n3182
        );

    \I__4788\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30575\
        );

    \I__4787\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30572\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__30575\,
            I => \N__30569\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__30572\,
            I => \N__30566\
        );

    \I__4784\ : Span4Mux_h
    port map (
            O => \N__30569\,
            I => \N__30562\
        );

    \I__4783\ : Span4Mux_v
    port map (
            O => \N__30566\,
            I => \N__30559\
        );

    \I__4782\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30556\
        );

    \I__4781\ : Span4Mux_v
    port map (
            O => \N__30562\,
            I => \N__30553\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__30559\,
            I => \N__30548\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__30556\,
            I => \N__30548\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__30553\,
            I => n309
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__30548\,
            I => n309
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__30543\,
            I => \n17_adj_710_cascade_\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__30540\,
            I => \n19_adj_711_cascade_\
        );

    \I__4774\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__30534\,
            I => n14236
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__30531\,
            I => \n14230_cascade_\
        );

    \I__4771\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__30525\,
            I => n61
        );

    \I__4769\ : CascadeMux
    port map (
            O => \N__30522\,
            I => \N__30519\
        );

    \I__4768\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30513\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__30513\,
            I => \N__30510\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__30510\,
            I => n2190
        );

    \I__4764\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30503\
        );

    \I__4763\ : CascadeMux
    port map (
            O => \N__30506\,
            I => \N__30500\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__30503\,
            I => \N__30496\
        );

    \I__4761\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30493\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__30499\,
            I => \N__30490\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__30496\,
            I => \N__30487\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__30493\,
            I => \N__30484\
        );

    \I__4757\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30481\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__30487\,
            I => n2228
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__30484\,
            I => n2228
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__30481\,
            I => n2228
        );

    \I__4753\ : CascadeMux
    port map (
            O => \N__30474\,
            I => \N__30471\
        );

    \I__4752\ : InMux
    port map (
            O => \N__30471\,
            I => \N__30468\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__30468\,
            I => \N__30464\
        );

    \I__4750\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30461\
        );

    \I__4749\ : Sp12to4
    port map (
            O => \N__30464\,
            I => \N__30456\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__30461\,
            I => \N__30456\
        );

    \I__4747\ : Odrv12
    port map (
            O => \N__30456\,
            I => n2224
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__30453\,
            I => \N__30448\
        );

    \I__4745\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30445\
        );

    \I__4744\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30442\
        );

    \I__4743\ : InMux
    port map (
            O => \N__30448\,
            I => \N__30439\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__30445\,
            I => \N__30436\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__30442\,
            I => n2227
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__30439\,
            I => n2227
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__30436\,
            I => n2227
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__30429\,
            I => \n14578_cascade_\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__30426\,
            I => \N__30423\
        );

    \I__4736\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30419\
        );

    \I__4735\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30416\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__30419\,
            I => \N__30413\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__30416\,
            I => \N__30410\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__30413\,
            I => n2225
        );

    \I__4731\ : Odrv12
    port map (
            O => \N__30410\,
            I => n2225
        );

    \I__4730\ : CascadeMux
    port map (
            O => \N__30405\,
            I => \N__30400\
        );

    \I__4729\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30397\
        );

    \I__4728\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30394\
        );

    \I__4727\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30391\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30388\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__30394\,
            I => n2223
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__30391\,
            I => n2223
        );

    \I__4723\ : Odrv4
    port map (
            O => \N__30388\,
            I => n2223
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__30381\,
            I => \N__30377\
        );

    \I__4721\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30373\
        );

    \I__4720\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30370\
        );

    \I__4719\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30367\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__30373\,
            I => n2222
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__30370\,
            I => n2222
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__30367\,
            I => n2222
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__30360\,
            I => \n14582_cascade_\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__30357\,
            I => \N__30354\
        );

    \I__4713\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30349\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__30353\,
            I => \N__30346\
        );

    \I__4711\ : InMux
    port map (
            O => \N__30352\,
            I => \N__30343\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__30349\,
            I => \N__30340\
        );

    \I__4709\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30337\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__30343\,
            I => \N__30334\
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__30340\,
            I => n2221
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__30337\,
            I => n2221
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__30334\,
            I => n2221
        );

    \I__4704\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30324\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__30324\,
            I => \N__30321\
        );

    \I__4702\ : Span4Mux_h
    port map (
            O => \N__30321\,
            I => \N__30316\
        );

    \I__4701\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30313\
        );

    \I__4700\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30310\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__30316\,
            I => n2220
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__30313\,
            I => n2220
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__30310\,
            I => n2220
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__30303\,
            I => \n14588_cascade_\
        );

    \I__4695\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__30297\,
            I => \N__30294\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__30294\,
            I => n14812
        );

    \I__4692\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__30288\,
            I => n14592
        );

    \I__4690\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30282\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__30282\,
            I => \N__30279\
        );

    \I__4688\ : Odrv4
    port map (
            O => \N__30279\,
            I => n2187
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__30276\,
            I => \N__30273\
        );

    \I__4686\ : InMux
    port map (
            O => \N__30273\,
            I => \N__30270\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__30270\,
            I => \N__30267\
        );

    \I__4684\ : Span4Mux_v
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__30264\,
            I => n2199
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__30261\,
            I => \N__30258\
        );

    \I__4681\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30255\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__30255\,
            I => n2285
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__30252\,
            I => \N__30248\
        );

    \I__4678\ : CascadeMux
    port map (
            O => \N__30251\,
            I => \N__30244\
        );

    \I__4677\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30241\
        );

    \I__4676\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30238\
        );

    \I__4675\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30235\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__30241\,
            I => \N__30232\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__30238\,
            I => \N__30227\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__30235\,
            I => \N__30227\
        );

    \I__4671\ : Span4Mux_v
    port map (
            O => \N__30232\,
            I => \N__30224\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__30227\,
            I => \N__30221\
        );

    \I__4669\ : Odrv4
    port map (
            O => \N__30224\,
            I => n2317
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__30221\,
            I => n2317
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__30216\,
            I => \N__30213\
        );

    \I__4666\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30210\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__4664\ : Span4Mux_v
    port map (
            O => \N__30207\,
            I => \N__30204\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__30204\,
            I => n2200
        );

    \I__4662\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30198\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__30195\,
            I => n2191
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__30192\,
            I => \N__30189\
        );

    \I__4658\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30186\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__30186\,
            I => \N__30183\
        );

    \I__4656\ : Span4Mux_v
    port map (
            O => \N__30183\,
            I => \N__30180\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__30180\,
            I => n2185
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__30177\,
            I => \N__30174\
        );

    \I__4653\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30169\
        );

    \I__4652\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30164\
        );

    \I__4651\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30164\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30161\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__30164\,
            I => \N__30158\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__30161\,
            I => n2218
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__30158\,
            I => n2218
        );

    \I__4646\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__30147\,
            I => \N__30142\
        );

    \I__4643\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30139\
        );

    \I__4642\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30136\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__30142\,
            I => n2219
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__30139\,
            I => n2219
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__30136\,
            I => n2219
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__30129\,
            I => \n2217_cascade_\
        );

    \I__4637\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30123\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__30123\,
            I => n14598
        );

    \I__4635\ : InMux
    port map (
            O => \N__30120\,
            I => \N__30117\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__4633\ : Odrv4
    port map (
            O => \N__30114\,
            I => n2188
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__30111\,
            I => \N__30108\
        );

    \I__4631\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30105\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__30105\,
            I => \N__30102\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__30102\,
            I => n2300
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__30099\,
            I => \N__30095\
        );

    \I__4627\ : InMux
    port map (
            O => \N__30098\,
            I => \N__30092\
        );

    \I__4626\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30089\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__30092\,
            I => \N__30086\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__30089\,
            I => \N__30083\
        );

    \I__4623\ : Span4Mux_h
    port map (
            O => \N__30086\,
            I => \N__30078\
        );

    \I__4622\ : Span4Mux_v
    port map (
            O => \N__30083\,
            I => \N__30078\
        );

    \I__4621\ : Span4Mux_v
    port map (
            O => \N__30078\,
            I => \N__30074\
        );

    \I__4620\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30071\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__30074\,
            I => n2332
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__30071\,
            I => n2332
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__30066\,
            I => \N__30063\
        );

    \I__4616\ : InMux
    port map (
            O => \N__30063\,
            I => \N__30060\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__30060\,
            I => n2290
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__30057\,
            I => \N__30053\
        );

    \I__4613\ : InMux
    port map (
            O => \N__30056\,
            I => \N__30050\
        );

    \I__4612\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30047\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__30050\,
            I => \N__30041\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__30047\,
            I => \N__30041\
        );

    \I__4609\ : InMux
    port map (
            O => \N__30046\,
            I => \N__30038\
        );

    \I__4608\ : Span4Mux_v
    port map (
            O => \N__30041\,
            I => \N__30033\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__30038\,
            I => \N__30033\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__30033\,
            I => n2322
        );

    \I__4605\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30026\
        );

    \I__4604\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30023\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__30026\,
            I => n2116
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__30023\,
            I => n2116
        );

    \I__4601\ : CascadeMux
    port map (
            O => \N__30018\,
            I => \n2117_cascade_\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__30015\,
            I => \n2148_cascade_\
        );

    \I__4599\ : InMux
    port map (
            O => \N__30012\,
            I => \N__30009\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__30009\,
            I => \N__30006\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__30006\,
            I => n2197
        );

    \I__4596\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29998\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__30002\,
            I => \N__29995\
        );

    \I__4594\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29992\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__29998\,
            I => \N__29989\
        );

    \I__4592\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29986\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__29992\,
            I => \N__29983\
        );

    \I__4590\ : Odrv12
    port map (
            O => \N__29989\,
            I => n2229
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__29986\,
            I => n2229
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__29983\,
            I => n2229
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__4586\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29970\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29967\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__29967\,
            I => n2189
        );

    \I__4583\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29961\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__29961\,
            I => n2184
        );

    \I__4581\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29954\
        );

    \I__4580\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29951\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__29954\,
            I => \N__29948\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__29951\,
            I => \N__29945\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__29948\,
            I => n2117
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__29945\,
            I => n2117
        );

    \I__4575\ : InMux
    port map (
            O => \N__29940\,
            I => \N__29936\
        );

    \I__4574\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29933\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__29936\,
            I => \N__29930\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__29933\,
            I => n2216
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__29930\,
            I => n2216
        );

    \I__4570\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29920\
        );

    \I__4569\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29917\
        );

    \I__4568\ : InMux
    port map (
            O => \N__29923\,
            I => \N__29914\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__29920\,
            I => \N__29911\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__29917\,
            I => \N__29906\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__29914\,
            I => \N__29906\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__29911\,
            I => n2215
        );

    \I__4563\ : Odrv4
    port map (
            O => \N__29906\,
            I => n2215
        );

    \I__4562\ : InMux
    port map (
            O => \N__29901\,
            I => \N__29898\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__29898\,
            I => \N__29894\
        );

    \I__4560\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29891\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__29894\,
            I => n2214
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__29891\,
            I => n2214
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__29886\,
            I => \n2216_cascade_\
        );

    \I__4556\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29880\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__29880\,
            I => n2298
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__29877\,
            I => \n2247_cascade_\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__29874\,
            I => \N__29869\
        );

    \I__4552\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29866\
        );

    \I__4551\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29863\
        );

    \I__4550\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29860\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29857\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29854\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__29860\,
            I => \N__29851\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__29857\,
            I => \N__29848\
        );

    \I__4545\ : Span4Mux_h
    port map (
            O => \N__29854\,
            I => \N__29843\
        );

    \I__4544\ : Span4Mux_v
    port map (
            O => \N__29851\,
            I => \N__29843\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__29848\,
            I => n2330
        );

    \I__4542\ : Odrv4
    port map (
            O => \N__29843\,
            I => n2330
        );

    \I__4541\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__29835\,
            I => n2193
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__29832\,
            I => \n2126_cascade_\
        );

    \I__4538\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29826\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__29826\,
            I => \N__29823\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__29823\,
            I => n2292
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__29820\,
            I => \n2225_cascade_\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__29817\,
            I => \N__29812\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__29816\,
            I => \N__29809\
        );

    \I__4532\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29806\
        );

    \I__4531\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29803\
        );

    \I__4530\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29800\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29797\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__29803\,
            I => \N__29794\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__29800\,
            I => \N__29791\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__29797\,
            I => \N__29788\
        );

    \I__4525\ : Odrv4
    port map (
            O => \N__29794\,
            I => n2324
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__29791\,
            I => n2324
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__29788\,
            I => n2324
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__29781\,
            I => \n2116_cascade_\
        );

    \I__4521\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29772\
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__29772\,
            I => n2183
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__29769\,
            I => \n2049_cascade_\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__29766\,
            I => \N__29763\
        );

    \I__4516\ : InMux
    port map (
            O => \N__29763\,
            I => \N__29760\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__29760\,
            I => n2186
        );

    \I__4514\ : InMux
    port map (
            O => \N__29757\,
            I => \N__29754\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__29754\,
            I => \N__29749\
        );

    \I__4512\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29746\
        );

    \I__4511\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29743\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__29749\,
            I => n3010
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__29746\,
            I => n3010
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__29743\,
            I => n3010
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__29736\,
            I => \N__29733\
        );

    \I__4506\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29730\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__29730\,
            I => \N__29727\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__29727\,
            I => n3077
        );

    \I__4503\ : CascadeMux
    port map (
            O => \N__29724\,
            I => \N__29721\
        );

    \I__4502\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29718\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__29718\,
            I => n2192
        );

    \I__4500\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29712\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__29712\,
            I => \N__29709\
        );

    \I__4498\ : Odrv4
    port map (
            O => \N__29709\,
            I => n2291
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__29706\,
            I => \n2224_cascade_\
        );

    \I__4496\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29698\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__29702\,
            I => \N__29695\
        );

    \I__4494\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29692\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__29698\,
            I => \N__29689\
        );

    \I__4492\ : InMux
    port map (
            O => \N__29695\,
            I => \N__29686\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__29692\,
            I => \N__29683\
        );

    \I__4490\ : Span4Mux_s2_h
    port map (
            O => \N__29689\,
            I => \N__29676\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__29686\,
            I => \N__29676\
        );

    \I__4488\ : Span4Mux_v
    port map (
            O => \N__29683\,
            I => \N__29676\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__29676\,
            I => n2323
        );

    \I__4486\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29670\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__29667\,
            I => \N__29662\
        );

    \I__4483\ : InMux
    port map (
            O => \N__29666\,
            I => \N__29659\
        );

    \I__4482\ : InMux
    port map (
            O => \N__29665\,
            I => \N__29656\
        );

    \I__4481\ : Odrv4
    port map (
            O => \N__29662\,
            I => n3009
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__29659\,
            I => n3009
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__29656\,
            I => n3009
        );

    \I__4478\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29645\
        );

    \I__4477\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29642\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__29645\,
            I => n3007
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__29642\,
            I => n3007
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__4473\ : InMux
    port map (
            O => \N__29634\,
            I => \N__29630\
        );

    \I__4472\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29627\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__29630\,
            I => \N__29624\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__29627\,
            I => \N__29620\
        );

    \I__4469\ : Span4Mux_h
    port map (
            O => \N__29624\,
            I => \N__29617\
        );

    \I__4468\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29614\
        );

    \I__4467\ : Span4Mux_h
    port map (
            O => \N__29620\,
            I => \N__29611\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__29617\,
            I => n3008
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__29614\,
            I => n3008
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__29611\,
            I => n3008
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__29604\,
            I => \n14754_cascade_\
        );

    \I__4462\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29598\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__29598\,
            I => \N__29594\
        );

    \I__4460\ : InMux
    port map (
            O => \N__29597\,
            I => \N__29591\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__29594\,
            I => \N__29588\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__29591\,
            I => n3006
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__29588\,
            I => n3006
        );

    \I__4456\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29580\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__29580\,
            I => \N__29577\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__29577\,
            I => n3079
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__29574\,
            I => \n3039_cascade_\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__29571\,
            I => \N__29566\
        );

    \I__4451\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29563\
        );

    \I__4450\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29558\
        );

    \I__4449\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29558\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__29563\,
            I => n3012
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__29558\,
            I => n3012
        );

    \I__4446\ : CascadeMux
    port map (
            O => \N__29553\,
            I => \n14194_cascade_\
        );

    \I__4445\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29547\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__29547\,
            I => n14196
        );

    \I__4443\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29537\
        );

    \I__4441\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29534\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__29537\,
            I => n3018
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__29534\,
            I => n3018
        );

    \I__4438\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__4436\ : Span4Mux_s1_v
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__4435\ : Odrv4
    port map (
            O => \N__29520\,
            I => n3085
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__29517\,
            I => \n3117_cascade_\
        );

    \I__4433\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29511\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__29511\,
            I => n14198
        );

    \I__4431\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29505\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__29505\,
            I => \N__29500\
        );

    \I__4429\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29497\
        );

    \I__4428\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29494\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__29500\,
            I => n3017
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__29497\,
            I => n3017
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__29494\,
            I => n3017
        );

    \I__4424\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__4422\ : Span4Mux_s1_v
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__29478\,
            I => n3084
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__29475\,
            I => \N__29471\
        );

    \I__4419\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29468\
        );

    \I__4418\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29465\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__29468\,
            I => \N__29462\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29459\
        );

    \I__4415\ : Span4Mux_s2_v
    port map (
            O => \N__29462\,
            I => \N__29454\
        );

    \I__4414\ : Span4Mux_h
    port map (
            O => \N__29459\,
            I => \N__29454\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__29454\,
            I => n3025
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__29451\,
            I => \N__29448\
        );

    \I__4411\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29445\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__4409\ : Span4Mux_s2_v
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__29439\,
            I => n3092
        );

    \I__4407\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29433\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__4405\ : Span4Mux_h
    port map (
            O => \N__29430\,
            I => \N__29427\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__29427\,
            I => n2999
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__29424\,
            I => \N__29421\
        );

    \I__4402\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29418\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__29418\,
            I => \N__29414\
        );

    \I__4400\ : CascadeMux
    port map (
            O => \N__29417\,
            I => \N__29411\
        );

    \I__4399\ : Span4Mux_h
    port map (
            O => \N__29414\,
            I => \N__29408\
        );

    \I__4398\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29405\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__29408\,
            I => n2932
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__29405\,
            I => n2932
        );

    \I__4395\ : CascadeMux
    port map (
            O => \N__29400\,
            I => \N__29397\
        );

    \I__4394\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29393\
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__29396\,
            I => \N__29390\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__29393\,
            I => \N__29387\
        );

    \I__4391\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29384\
        );

    \I__4390\ : Span4Mux_v
    port map (
            O => \N__29387\,
            I => \N__29381\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__29384\,
            I => n3031
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__29381\,
            I => n3031
        );

    \I__4387\ : InMux
    port map (
            O => \N__29376\,
            I => \N__29373\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__29373\,
            I => \N__29370\
        );

    \I__4385\ : Span4Mux_s3_v
    port map (
            O => \N__29370\,
            I => \N__29367\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__29367\,
            I => n3098
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__29364\,
            I => \n3031_cascade_\
        );

    \I__4382\ : InMux
    port map (
            O => \N__29361\,
            I => \N__29357\
        );

    \I__4381\ : InMux
    port map (
            O => \N__29360\,
            I => \N__29353\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__29357\,
            I => \N__29350\
        );

    \I__4379\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29347\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__29353\,
            I => \N__29344\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__29350\,
            I => \N__29341\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__29347\,
            I => \N__29338\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__29344\,
            I => \N__29335\
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__29341\,
            I => n2916
        );

    \I__4373\ : Odrv12
    port map (
            O => \N__29338\,
            I => n2916
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__29335\,
            I => n2916
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__29328\,
            I => \N__29325\
        );

    \I__4370\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29322\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__29322\,
            I => \N__29319\
        );

    \I__4368\ : Span4Mux_h
    port map (
            O => \N__29319\,
            I => \N__29316\
        );

    \I__4367\ : Odrv4
    port map (
            O => \N__29316\,
            I => n2983
        );

    \I__4366\ : InMux
    port map (
            O => \N__29313\,
            I => \N__29310\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__4364\ : Span4Mux_s2_v
    port map (
            O => \N__29307\,
            I => \N__29303\
        );

    \I__4363\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29300\
        );

    \I__4362\ : Odrv4
    port map (
            O => \N__29303\,
            I => n3015
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__29300\,
            I => n3015
        );

    \I__4360\ : InMux
    port map (
            O => \N__29295\,
            I => \N__29292\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__29292\,
            I => \N__29289\
        );

    \I__4358\ : Span4Mux_h
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__29286\,
            I => n3082
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__29283\,
            I => \n3015_cascade_\
        );

    \I__4355\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29277\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__29277\,
            I => \N__29274\
        );

    \I__4353\ : Span4Mux_s2_v
    port map (
            O => \N__29274\,
            I => \N__29271\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__29271\,
            I => n3089
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__29268\,
            I => \N__29265\
        );

    \I__4350\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29261\
        );

    \I__4349\ : InMux
    port map (
            O => \N__29264\,
            I => \N__29258\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__29261\,
            I => \N__29255\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__29258\,
            I => \N__29252\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__29255\,
            I => n3022
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__29252\,
            I => n3022
        );

    \I__4344\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29244\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__29241\,
            I => \N__29238\
        );

    \I__4341\ : Odrv4
    port map (
            O => \N__29238\,
            I => n3095
        );

    \I__4340\ : CascadeMux
    port map (
            O => \N__29235\,
            I => \N__29230\
        );

    \I__4339\ : InMux
    port map (
            O => \N__29234\,
            I => \N__29227\
        );

    \I__4338\ : InMux
    port map (
            O => \N__29233\,
            I => \N__29224\
        );

    \I__4337\ : InMux
    port map (
            O => \N__29230\,
            I => \N__29221\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__29227\,
            I => \N__29216\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__29224\,
            I => \N__29216\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__29221\,
            I => n3028
        );

    \I__4333\ : Odrv4
    port map (
            O => \N__29216\,
            I => n3028
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__29211\,
            I => \n3127_cascade_\
        );

    \I__4331\ : InMux
    port map (
            O => \N__29208\,
            I => \N__29203\
        );

    \I__4330\ : InMux
    port map (
            O => \N__29207\,
            I => \N__29200\
        );

    \I__4329\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29197\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__29203\,
            I => n3011
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__29200\,
            I => n3011
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__29197\,
            I => n3011
        );

    \I__4325\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29187\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__29187\,
            I => n14744
        );

    \I__4323\ : InMux
    port map (
            O => \N__29184\,
            I => \N__29181\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__29181\,
            I => n14816
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__29178\,
            I => \n14750_cascade_\
        );

    \I__4320\ : InMux
    port map (
            O => \N__29175\,
            I => \N__29172\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__29172\,
            I => \N__29167\
        );

    \I__4318\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29164\
        );

    \I__4317\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29161\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__29167\,
            I => n3014
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__29164\,
            I => n3014
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__29161\,
            I => n3014
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__4312\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__4310\ : Span4Mux_v
    port map (
            O => \N__29145\,
            I => \N__29142\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__29142\,
            I => n3081
        );

    \I__4308\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29136\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__29133\,
            I => n3100
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__4304\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29124\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__29124\,
            I => \N__29121\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__29121\,
            I => n3001
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__29118\,
            I => \N__29115\
        );

    \I__4300\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29111\
        );

    \I__4299\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29108\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__29111\,
            I => \N__29105\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__29108\,
            I => n3033
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__29105\,
            I => n3033
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__29100\,
            I => \n3033_cascade_\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__29097\,
            I => \N__29094\
        );

    \I__4293\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29089\
        );

    \I__4292\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29084\
        );

    \I__4291\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29084\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29079\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29079\
        );

    \I__4288\ : Span4Mux_h
    port map (
            O => \N__29079\,
            I => \N__29076\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__29076\,
            I => n3032
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__29073\,
            I => \N__29070\
        );

    \I__4285\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29067\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__29067\,
            I => \N__29064\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__29064\,
            I => n2990
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__29061\,
            I => \n3022_cascade_\
        );

    \I__4281\ : InMux
    port map (
            O => \N__29058\,
            I => \N__29055\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__29055\,
            I => n14732
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__29052\,
            I => \N__29049\
        );

    \I__4278\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29045\
        );

    \I__4277\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29042\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__29045\,
            I => n3030
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__29042\,
            I => n3030
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__29037\,
            I => \N__29034\
        );

    \I__4273\ : InMux
    port map (
            O => \N__29034\,
            I => \N__29030\
        );

    \I__4272\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29027\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__29030\,
            I => n3029
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__29027\,
            I => n3029
        );

    \I__4269\ : InMux
    port map (
            O => \N__29022\,
            I => \N__29019\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__29019\,
            I => n11932
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__29016\,
            I => \n13859_cascade_\
        );

    \I__4266\ : InMux
    port map (
            O => \N__29013\,
            I => \N__29010\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__29010\,
            I => n14738
        );

    \I__4264\ : InMux
    port map (
            O => \N__29007\,
            I => n12904
        );

    \I__4263\ : InMux
    port map (
            O => \N__29004\,
            I => n12905
        );

    \I__4262\ : InMux
    port map (
            O => \N__29001\,
            I => n12906
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__28998\,
            I => \N__28995\
        );

    \I__4260\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28992\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__28992\,
            I => \N__28989\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__28989\,
            I => n3180
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__28986\,
            I => \N__28982\
        );

    \I__4256\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28979\
        );

    \I__4255\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28976\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__28979\,
            I => \N__28972\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__28976\,
            I => \N__28969\
        );

    \I__4252\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28966\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__28972\,
            I => n2925
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__28969\,
            I => n2925
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__28966\,
            I => n2925
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__28959\,
            I => \N__28956\
        );

    \I__4247\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28953\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__28953\,
            I => \N__28950\
        );

    \I__4245\ : Span4Mux_h
    port map (
            O => \N__28950\,
            I => \N__28947\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__28947\,
            I => n2992
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__4242\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28938\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__28938\,
            I => \N__28935\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__28935\,
            I => n3099
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__28932\,
            I => \N__28929\
        );

    \I__4238\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28926\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__28926\,
            I => \N__28923\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__28923\,
            I => \N__28920\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__28920\,
            I => n3076
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__28917\,
            I => \N__28914\
        );

    \I__4233\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28910\
        );

    \I__4232\ : InMux
    port map (
            O => \N__28913\,
            I => \N__28907\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__28910\,
            I => \N__28904\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__28907\,
            I => \N__28901\
        );

    \I__4229\ : Span4Mux_s3_h
    port map (
            O => \N__28904\,
            I => \N__28898\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__28901\,
            I => n2926
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__28898\,
            I => n2926
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__28893\,
            I => \N__28890\
        );

    \I__4225\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28887\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__4223\ : Span4Mux_v
    port map (
            O => \N__28884\,
            I => \N__28881\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__28881\,
            I => n2993
        );

    \I__4221\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28874\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__28877\,
            I => \N__28871\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__28874\,
            I => \N__28867\
        );

    \I__4218\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28864\
        );

    \I__4217\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28861\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__28867\,
            I => n3027
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__28864\,
            I => n3027
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__28861\,
            I => n3027
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__28854\,
            I => \n3025_cascade_\
        );

    \I__4212\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28848\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__28848\,
            I => n14736
        );

    \I__4210\ : InMux
    port map (
            O => \N__28845\,
            I => n12895
        );

    \I__4209\ : InMux
    port map (
            O => \N__28842\,
            I => n12896
        );

    \I__4208\ : InMux
    port map (
            O => \N__28839\,
            I => n12897
        );

    \I__4207\ : InMux
    port map (
            O => \N__28836\,
            I => n12898
        );

    \I__4206\ : InMux
    port map (
            O => \N__28833\,
            I => n12899
        );

    \I__4205\ : InMux
    port map (
            O => \N__28830\,
            I => n12900
        );

    \I__4204\ : InMux
    port map (
            O => \N__28827\,
            I => \bfn_5_28_0_\
        );

    \I__4203\ : InMux
    port map (
            O => \N__28824\,
            I => n12902
        );

    \I__4202\ : InMux
    port map (
            O => \N__28821\,
            I => n12903
        );

    \I__4201\ : InMux
    port map (
            O => \N__28818\,
            I => n12886
        );

    \I__4200\ : InMux
    port map (
            O => \N__28815\,
            I => n12887
        );

    \I__4199\ : InMux
    port map (
            O => \N__28812\,
            I => n12888
        );

    \I__4198\ : InMux
    port map (
            O => \N__28809\,
            I => n12889
        );

    \I__4197\ : InMux
    port map (
            O => \N__28806\,
            I => n12890
        );

    \I__4196\ : InMux
    port map (
            O => \N__28803\,
            I => n12891
        );

    \I__4195\ : InMux
    port map (
            O => \N__28800\,
            I => n12892
        );

    \I__4194\ : InMux
    port map (
            O => \N__28797\,
            I => \bfn_5_27_0_\
        );

    \I__4193\ : InMux
    port map (
            O => \N__28794\,
            I => n12894
        );

    \I__4192\ : InMux
    port map (
            O => \N__28791\,
            I => \bfn_5_25_0_\
        );

    \I__4191\ : InMux
    port map (
            O => \N__28788\,
            I => n12878
        );

    \I__4190\ : InMux
    port map (
            O => \N__28785\,
            I => n12879
        );

    \I__4189\ : InMux
    port map (
            O => \N__28782\,
            I => n12880
        );

    \I__4188\ : InMux
    port map (
            O => \N__28779\,
            I => n12881
        );

    \I__4187\ : InMux
    port map (
            O => \N__28776\,
            I => n12882
        );

    \I__4186\ : InMux
    port map (
            O => \N__28773\,
            I => n12883
        );

    \I__4185\ : InMux
    port map (
            O => \N__28770\,
            I => n12884
        );

    \I__4184\ : InMux
    port map (
            O => \N__28767\,
            I => \bfn_5_26_0_\
        );

    \I__4183\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28761\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__28761\,
            I => \N__28758\
        );

    \I__4181\ : Odrv4
    port map (
            O => \N__28758\,
            I => n2289
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__28755\,
            I => \N__28751\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__28754\,
            I => \N__28748\
        );

    \I__4178\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28745\
        );

    \I__4177\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28741\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__28745\,
            I => \N__28738\
        );

    \I__4175\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28735\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__28741\,
            I => \N__28732\
        );

    \I__4173\ : Span4Mux_v
    port map (
            O => \N__28738\,
            I => \N__28729\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__28735\,
            I => \N__28726\
        );

    \I__4171\ : Span4Mux_v
    port map (
            O => \N__28732\,
            I => \N__28723\
        );

    \I__4170\ : Span4Mux_v
    port map (
            O => \N__28729\,
            I => \N__28718\
        );

    \I__4169\ : Span4Mux_v
    port map (
            O => \N__28726\,
            I => \N__28718\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__28723\,
            I => n2321
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__28718\,
            I => n2321
        );

    \I__4166\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28709\
        );

    \I__4165\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28706\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__28709\,
            I => \N__28702\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__28706\,
            I => \N__28699\
        );

    \I__4162\ : CascadeMux
    port map (
            O => \N__28705\,
            I => \N__28696\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__28702\,
            I => \N__28691\
        );

    \I__4160\ : Span4Mux_v
    port map (
            O => \N__28699\,
            I => \N__28691\
        );

    \I__4159\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28688\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__28691\,
            I => n2331
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__28688\,
            I => n2331
        );

    \I__4156\ : InMux
    port map (
            O => \N__28683\,
            I => \N__28680\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__28680\,
            I => \N__28677\
        );

    \I__4154\ : Span4Mux_h
    port map (
            O => \N__28677\,
            I => \N__28674\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__28674\,
            I => n11954
        );

    \I__4152\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28666\
        );

    \I__4151\ : InMux
    port map (
            O => \N__28670\,
            I => \N__28663\
        );

    \I__4150\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28660\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28655\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28655\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__28660\,
            I => \N__28652\
        );

    \I__4146\ : Span4Mux_v
    port map (
            O => \N__28655\,
            I => \N__28649\
        );

    \I__4145\ : Span4Mux_h
    port map (
            O => \N__28652\,
            I => \N__28646\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__28649\,
            I => \N__28643\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__28646\,
            I => n311
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__28643\,
            I => n311
        );

    \I__4141\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28634\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__28637\,
            I => \N__28631\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__28634\,
            I => \N__28628\
        );

    \I__4138\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28625\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__28628\,
            I => \N__28622\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__28625\,
            I => \N__28619\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__28622\,
            I => \N__28613\
        );

    \I__4134\ : Span4Mux_v
    port map (
            O => \N__28619\,
            I => \N__28613\
        );

    \I__4133\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28610\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__28613\,
            I => n2533
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__28610\,
            I => n2533
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__28605\,
            I => \N__28602\
        );

    \I__4129\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__4127\ : Span4Mux_v
    port map (
            O => \N__28596\,
            I => \N__28593\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__28593\,
            I => n2600
        );

    \I__4125\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28587\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__28587\,
            I => \N__28583\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__28586\,
            I => \N__28580\
        );

    \I__4122\ : Span4Mux_h
    port map (
            O => \N__28583\,
            I => \N__28577\
        );

    \I__4121\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28574\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__28577\,
            I => \N__28569\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__28574\,
            I => \N__28569\
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__28569\,
            I => n2532
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__28566\,
            I => \N__28563\
        );

    \I__4116\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28560\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__28557\,
            I => \N__28554\
        );

    \I__4113\ : Odrv4
    port map (
            O => \N__28554\,
            I => n2599
        );

    \I__4112\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28547\
        );

    \I__4111\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28544\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__28547\,
            I => \N__28541\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__28544\,
            I => n2631
        );

    \I__4108\ : Odrv4
    port map (
            O => \N__28541\,
            I => n2631
        );

    \I__4107\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28531\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__28535\,
            I => \N__28528\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__28534\,
            I => \N__28525\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__28531\,
            I => \N__28522\
        );

    \I__4103\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28519\
        );

    \I__4102\ : InMux
    port map (
            O => \N__28525\,
            I => \N__28516\
        );

    \I__4101\ : Span4Mux_v
    port map (
            O => \N__28522\,
            I => \N__28513\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__28519\,
            I => n2633
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__28516\,
            I => n2633
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__28513\,
            I => n2633
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__28506\,
            I => \n2631_cascade_\
        );

    \I__4096\ : InMux
    port map (
            O => \N__28503\,
            I => \N__28499\
        );

    \I__4095\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28495\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__28499\,
            I => \N__28492\
        );

    \I__4093\ : InMux
    port map (
            O => \N__28498\,
            I => \N__28489\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__28495\,
            I => n2632
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__28492\,
            I => n2632
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__28489\,
            I => n2632
        );

    \I__4089\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28479\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__28476\,
            I => \N__28473\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__28473\,
            I => n12044
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__28470\,
            I => \N__28467\
        );

    \I__4084\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28464\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__28464\,
            I => \N__28461\
        );

    \I__4082\ : Odrv12
    port map (
            O => \N__28461\,
            I => n2301
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__4080\ : InMux
    port map (
            O => \N__28455\,
            I => \N__28451\
        );

    \I__4079\ : InMux
    port map (
            O => \N__28454\,
            I => \N__28448\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__28451\,
            I => \N__28445\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__28448\,
            I => \N__28442\
        );

    \I__4076\ : Span12Mux_v
    port map (
            O => \N__28445\,
            I => \N__28438\
        );

    \I__4075\ : Sp12to4
    port map (
            O => \N__28442\,
            I => \N__28435\
        );

    \I__4074\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28432\
        );

    \I__4073\ : Odrv12
    port map (
            O => \N__28438\,
            I => n2333
        );

    \I__4072\ : Odrv12
    port map (
            O => \N__28435\,
            I => n2333
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__28432\,
            I => n2333
        );

    \I__4070\ : InMux
    port map (
            O => \N__28425\,
            I => \bfn_5_22_0_\
        );

    \I__4069\ : InMux
    port map (
            O => \N__28422\,
            I => n12678
        );

    \I__4068\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28416\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__28416\,
            I => \N__28413\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__28413\,
            I => n2283
        );

    \I__4065\ : InMux
    port map (
            O => \N__28410\,
            I => n12679
        );

    \I__4064\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__28404\,
            I => \N__28401\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__28401\,
            I => \N__28398\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__28398\,
            I => n2282
        );

    \I__4060\ : InMux
    port map (
            O => \N__28395\,
            I => n12680
        );

    \I__4059\ : InMux
    port map (
            O => \N__28392\,
            I => n12681
        );

    \I__4058\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28385\
        );

    \I__4057\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28382\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28379\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__28382\,
            I => \N__28376\
        );

    \I__4054\ : Span4Mux_v
    port map (
            O => \N__28379\,
            I => \N__28373\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__28376\,
            I => n2313
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__28373\,
            I => n2313
        );

    \I__4051\ : InMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__28365\,
            I => \N__28362\
        );

    \I__4049\ : Odrv4
    port map (
            O => \N__28362\,
            I => n2299
        );

    \I__4048\ : InMux
    port map (
            O => \N__28359\,
            I => \N__28356\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__28350\,
            I => n2196
        );

    \I__4044\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__4042\ : Odrv12
    port map (
            O => \N__28341\,
            I => n2198
        );

    \I__4041\ : InMux
    port map (
            O => \N__28338\,
            I => \N__28335\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__28335\,
            I => \N__28331\
        );

    \I__4039\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28328\
        );

    \I__4038\ : Span4Mux_h
    port map (
            O => \N__28331\,
            I => \N__28325\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__28328\,
            I => \N__28322\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__28325\,
            I => n2230
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__28322\,
            I => n2230
        );

    \I__4034\ : CascadeMux
    port map (
            O => \N__28317\,
            I => \n2230_cascade_\
        );

    \I__4033\ : InMux
    port map (
            O => \N__28314\,
            I => n12668
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__4031\ : InMux
    port map (
            O => \N__28308\,
            I => \N__28305\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__28305\,
            I => \N__28302\
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__28302\,
            I => n2293
        );

    \I__4028\ : InMux
    port map (
            O => \N__28299\,
            I => \bfn_5_21_0_\
        );

    \I__4027\ : InMux
    port map (
            O => \N__28296\,
            I => n12670
        );

    \I__4026\ : InMux
    port map (
            O => \N__28293\,
            I => n12671
        );

    \I__4025\ : InMux
    port map (
            O => \N__28290\,
            I => n12672
        );

    \I__4024\ : InMux
    port map (
            O => \N__28287\,
            I => n12673
        );

    \I__4023\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28281\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__28281\,
            I => n2288
        );

    \I__4021\ : InMux
    port map (
            O => \N__28278\,
            I => n12674
        );

    \I__4020\ : InMux
    port map (
            O => \N__28275\,
            I => \N__28272\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__28272\,
            I => n2287
        );

    \I__4018\ : InMux
    port map (
            O => \N__28269\,
            I => n12675
        );

    \I__4017\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28263\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__28263\,
            I => n2286
        );

    \I__4015\ : InMux
    port map (
            O => \N__28260\,
            I => n12676
        );

    \I__4014\ : InMux
    port map (
            O => \N__28257\,
            I => \N__28254\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__28254\,
            I => \N__28251\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__28251\,
            I => n2195
        );

    \I__4011\ : InMux
    port map (
            O => \N__28248\,
            I => \bfn_5_20_0_\
        );

    \I__4010\ : InMux
    port map (
            O => \N__28245\,
            I => n12662
        );

    \I__4009\ : InMux
    port map (
            O => \N__28242\,
            I => n12663
        );

    \I__4008\ : InMux
    port map (
            O => \N__28239\,
            I => n12664
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__4006\ : InMux
    port map (
            O => \N__28233\,
            I => \N__28230\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__28230\,
            I => \N__28227\
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__28227\,
            I => n2297
        );

    \I__4003\ : InMux
    port map (
            O => \N__28224\,
            I => n12665
        );

    \I__4002\ : InMux
    port map (
            O => \N__28221\,
            I => \N__28218\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__28218\,
            I => \N__28215\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__28215\,
            I => n2296
        );

    \I__3999\ : InMux
    port map (
            O => \N__28212\,
            I => n12666
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__28209\,
            I => \N__28206\
        );

    \I__3997\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28203\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__28203\,
            I => n2295
        );

    \I__3995\ : InMux
    port map (
            O => \N__28200\,
            I => n12667
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__28197\,
            I => \N__28194\
        );

    \I__3993\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28191\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__28191\,
            I => n2294
        );

    \I__3991\ : InMux
    port map (
            O => \N__28188\,
            I => n12655
        );

    \I__3990\ : InMux
    port map (
            O => \N__28185\,
            I => n12656
        );

    \I__3989\ : InMux
    port map (
            O => \N__28182\,
            I => n12657
        );

    \I__3988\ : InMux
    port map (
            O => \N__28179\,
            I => \bfn_5_19_0_\
        );

    \I__3987\ : InMux
    port map (
            O => \N__28176\,
            I => n12659
        );

    \I__3986\ : InMux
    port map (
            O => \N__28173\,
            I => n12660
        );

    \I__3985\ : InMux
    port map (
            O => \N__28170\,
            I => n12661
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__28167\,
            I => \N__28163\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__28166\,
            I => \N__28159\
        );

    \I__3982\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28154\
        );

    \I__3981\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28154\
        );

    \I__3980\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28151\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__28154\,
            I => \N__28148\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__28151\,
            I => n2315
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__28148\,
            I => n2315
        );

    \I__3976\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__28140\,
            I => \N__28136\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__28139\,
            I => \N__28133\
        );

    \I__3973\ : Span4Mux_h
    port map (
            O => \N__28136\,
            I => \N__28129\
        );

    \I__3972\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28126\
        );

    \I__3971\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28123\
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__28129\,
            I => n2325
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__28126\,
            I => n2325
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__28123\,
            I => n2325
        );

    \I__3967\ : InMux
    port map (
            O => \N__28116\,
            I => n12645
        );

    \I__3966\ : InMux
    port map (
            O => \N__28113\,
            I => n12646
        );

    \I__3965\ : InMux
    port map (
            O => \N__28110\,
            I => n12647
        );

    \I__3964\ : InMux
    port map (
            O => \N__28107\,
            I => n12648
        );

    \I__3963\ : InMux
    port map (
            O => \N__28104\,
            I => n12649
        );

    \I__3962\ : InMux
    port map (
            O => \N__28101\,
            I => \bfn_5_18_0_\
        );

    \I__3961\ : InMux
    port map (
            O => \N__28098\,
            I => n12651
        );

    \I__3960\ : InMux
    port map (
            O => \N__28095\,
            I => n12652
        );

    \I__3959\ : InMux
    port map (
            O => \N__28092\,
            I => n12653
        );

    \I__3958\ : InMux
    port map (
            O => \N__28089\,
            I => n12654
        );

    \I__3957\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28082\
        );

    \I__3956\ : InMux
    port map (
            O => \N__28085\,
            I => \N__28079\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__28082\,
            I => \N__28076\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28070\
        );

    \I__3953\ : Span4Mux_s3_h
    port map (
            O => \N__28076\,
            I => \N__28070\
        );

    \I__3952\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28067\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__28070\,
            I => \N__28062\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__28067\,
            I => \N__28062\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__28059\,
            I => n2908
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__28056\,
            I => \N__28053\
        );

    \I__3946\ : InMux
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__28050\,
            I => \N__28047\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__28047\,
            I => n2975
        );

    \I__3943\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28041\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__28041\,
            I => n3074
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__28038\,
            I => \n3007_cascade_\
        );

    \I__3940\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28032\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__28032\,
            I => \N__28028\
        );

    \I__3938\ : InMux
    port map (
            O => \N__28031\,
            I => \N__28025\
        );

    \I__3937\ : Span12Mux_s4_v
    port map (
            O => \N__28028\,
            I => \N__28021\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__28025\,
            I => \N__28018\
        );

    \I__3935\ : InMux
    port map (
            O => \N__28024\,
            I => \N__28015\
        );

    \I__3934\ : Odrv12
    port map (
            O => \N__28021\,
            I => n2910
        );

    \I__3933\ : Odrv12
    port map (
            O => \N__28018\,
            I => n2910
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__28015\,
            I => n2910
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__28008\,
            I => \N__28005\
        );

    \I__3930\ : InMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__28002\,
            I => \N__27999\
        );

    \I__3928\ : Odrv12
    port map (
            O => \N__27999\,
            I => n2977
        );

    \I__3927\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27992\
        );

    \I__3926\ : InMux
    port map (
            O => \N__27995\,
            I => \N__27989\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__27992\,
            I => \N__27984\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__27989\,
            I => \N__27984\
        );

    \I__3923\ : Span4Mux_s2_v
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__27981\,
            I => \debounce.reg_A_2\
        );

    \I__3921\ : SRMux
    port map (
            O => \N__27978\,
            I => \N__27975\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__27975\,
            I => \N__27971\
        );

    \I__3919\ : SRMux
    port map (
            O => \N__27974\,
            I => \N__27968\
        );

    \I__3918\ : Span4Mux_v
    port map (
            O => \N__27971\,
            I => \N__27965\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27962\
        );

    \I__3916\ : Span4Mux_s1_h
    port map (
            O => \N__27965\,
            I => \N__27957\
        );

    \I__3915\ : Span4Mux_s1_h
    port map (
            O => \N__27962\,
            I => \N__27957\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__27957\,
            I => \debounce.cnt_next_9__N_424\
        );

    \I__3913\ : InMux
    port map (
            O => \N__27954\,
            I => \bfn_5_17_0_\
        );

    \I__3912\ : InMux
    port map (
            O => \N__27951\,
            I => n12643
        );

    \I__3911\ : InMux
    port map (
            O => \N__27948\,
            I => n12644
        );

    \I__3910\ : InMux
    port map (
            O => \N__27945\,
            I => \N__27942\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__27942\,
            I => \N__27939\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__27939\,
            I => \N__27936\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__27936\,
            I => n2985
        );

    \I__3906\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27929\
        );

    \I__3905\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27926\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27923\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27920\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__27923\,
            I => \N__27917\
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__27920\,
            I => n2918
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__27917\,
            I => n2918
        );

    \I__3899\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27908\
        );

    \I__3898\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27905\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__27908\,
            I => \N__27902\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__27905\,
            I => \N__27899\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__27902\,
            I => n2911
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__27899\,
            I => n2911
        );

    \I__3893\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27891\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__27891\,
            I => \N__27888\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__27888\,
            I => n2978
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__27885\,
            I => \N__27881\
        );

    \I__3889\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27878\
        );

    \I__3888\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27875\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__27878\,
            I => \N__27872\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__27875\,
            I => \N__27869\
        );

    \I__3885\ : Span4Mux_s3_v
    port map (
            O => \N__27872\,
            I => \N__27865\
        );

    \I__3884\ : Span4Mux_s2_h
    port map (
            O => \N__27869\,
            I => \N__27862\
        );

    \I__3883\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27859\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__27865\,
            I => n2825
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__27862\,
            I => n2825
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__27859\,
            I => n2825
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__27852\,
            I => \N__27849\
        );

    \I__3878\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27846\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__27846\,
            I => \N__27843\
        );

    \I__3876\ : Span4Mux_v
    port map (
            O => \N__27843\,
            I => \N__27840\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__27840\,
            I => n2892
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__27837\,
            I => \N__27834\
        );

    \I__3873\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27830\
        );

    \I__3872\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27826\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__27830\,
            I => \N__27823\
        );

    \I__3870\ : InMux
    port map (
            O => \N__27829\,
            I => \N__27820\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__27826\,
            I => \N__27817\
        );

    \I__3868\ : Span4Mux_v
    port map (
            O => \N__27823\,
            I => \N__27814\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__27820\,
            I => \N__27809\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__27817\,
            I => \N__27809\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__27814\,
            I => n2924
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__27809\,
            I => n2924
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__27804\,
            I => \N__27801\
        );

    \I__3862\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27797\
        );

    \I__3861\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27794\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__27797\,
            I => \N__27791\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__27794\,
            I => \N__27787\
        );

    \I__3858\ : Span4Mux_v
    port map (
            O => \N__27791\,
            I => \N__27784\
        );

    \I__3857\ : InMux
    port map (
            O => \N__27790\,
            I => \N__27781\
        );

    \I__3856\ : Odrv12
    port map (
            O => \N__27787\,
            I => n2913
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__27784\,
            I => n2913
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__27781\,
            I => n2913
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__27774\,
            I => \N__27771\
        );

    \I__3852\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27768\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__3850\ : Odrv12
    port map (
            O => \N__27765\,
            I => n2980
        );

    \I__3849\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27758\
        );

    \I__3848\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27755\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__27758\,
            I => \N__27752\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27746\
        );

    \I__3845\ : Span4Mux_s3_h
    port map (
            O => \N__27752\,
            I => \N__27746\
        );

    \I__3844\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27743\
        );

    \I__3843\ : Span4Mux_v
    port map (
            O => \N__27746\,
            I => \N__27740\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__27743\,
            I => \N__27737\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__27740\,
            I => n2915
        );

    \I__3840\ : Odrv12
    port map (
            O => \N__27737\,
            I => n2915
        );

    \I__3839\ : CascadeMux
    port map (
            O => \N__27732\,
            I => \N__27729\
        );

    \I__3838\ : InMux
    port map (
            O => \N__27729\,
            I => \N__27726\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27723\
        );

    \I__3836\ : Odrv4
    port map (
            O => \N__27723\,
            I => n2982
        );

    \I__3835\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27717\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__27717\,
            I => \N__27713\
        );

    \I__3833\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27710\
        );

    \I__3832\ : Span4Mux_h
    port map (
            O => \N__27713\,
            I => \N__27704\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27704\
        );

    \I__3830\ : InMux
    port map (
            O => \N__27709\,
            I => \N__27701\
        );

    \I__3829\ : Odrv4
    port map (
            O => \N__27704\,
            I => n2912
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__27701\,
            I => n2912
        );

    \I__3827\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27693\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__27693\,
            I => \N__27690\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__27690\,
            I => n2979
        );

    \I__3824\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27683\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__27686\,
            I => \N__27680\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__27683\,
            I => \N__27677\
        );

    \I__3821\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27674\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__27677\,
            I => \N__27670\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__27674\,
            I => \N__27667\
        );

    \I__3818\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27664\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__27670\,
            I => n2919
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__27667\,
            I => n2919
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__27664\,
            I => n2919
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__27657\,
            I => \N__27654\
        );

    \I__3813\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27651\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__27651\,
            I => \N__27648\
        );

    \I__3811\ : Span4Mux_s2_v
    port map (
            O => \N__27648\,
            I => \N__27645\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__27645\,
            I => n2986
        );

    \I__3809\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27637\
        );

    \I__3808\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27634\
        );

    \I__3807\ : InMux
    port map (
            O => \N__27640\,
            I => \N__27631\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__27637\,
            I => n3016
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__27634\,
            I => n3016
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__27631\,
            I => n3016
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__27624\,
            I => \n3018_cascade_\
        );

    \I__3802\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__27618\,
            I => \N__27614\
        );

    \I__3800\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27611\
        );

    \I__3799\ : Span4Mux_s1_v
    port map (
            O => \N__27614\,
            I => \N__27607\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__27611\,
            I => \N__27604\
        );

    \I__3797\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27601\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__27607\,
            I => n2914
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__27604\,
            I => n2914
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__27601\,
            I => n2914
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__27594\,
            I => \N__27591\
        );

    \I__3792\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27588\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27585\
        );

    \I__3790\ : Span4Mux_s1_v
    port map (
            O => \N__27585\,
            I => \N__27582\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__27582\,
            I => n2981
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__27579\,
            I => \N__27576\
        );

    \I__3787\ : InMux
    port map (
            O => \N__27576\,
            I => \N__27572\
        );

    \I__3786\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27568\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__27572\,
            I => \N__27565\
        );

    \I__3784\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27562\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__27568\,
            I => n3019
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__27565\,
            I => n3019
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__27562\,
            I => n3019
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__27555\,
            I => \n3023_cascade_\
        );

    \I__3779\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27548\
        );

    \I__3778\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27545\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__27548\,
            I => \N__27541\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27538\
        );

    \I__3775\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27535\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__27541\,
            I => n2922
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__27538\,
            I => n2922
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__27535\,
            I => n2922
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__3770\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27522\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__27522\,
            I => \N__27519\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__27519\,
            I => \N__27516\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__27516\,
            I => n2989
        );

    \I__3766\ : CascadeMux
    port map (
            O => \N__27513\,
            I => \N__27510\
        );

    \I__3765\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27507\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__27507\,
            I => n3078
        );

    \I__3763\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__27501\,
            I => \N__27498\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__27498\,
            I => n3075
        );

    \I__3760\ : InMux
    port map (
            O => \N__27495\,
            I => \N__27492\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__27492\,
            I => \N__27489\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__27486\,
            I => n2984
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__27483\,
            I => \N__27479\
        );

    \I__3755\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27476\
        );

    \I__3754\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27473\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27470\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__27473\,
            I => \N__27466\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__27470\,
            I => \N__27463\
        );

    \I__3750\ : InMux
    port map (
            O => \N__27469\,
            I => \N__27460\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__27466\,
            I => n2917
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__27463\,
            I => n2917
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__27460\,
            I => n2917
        );

    \I__3746\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27449\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__27452\,
            I => \N__27446\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__27449\,
            I => \N__27442\
        );

    \I__3743\ : InMux
    port map (
            O => \N__27446\,
            I => \N__27439\
        );

    \I__3742\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27436\
        );

    \I__3741\ : Odrv12
    port map (
            O => \N__27442\,
            I => n2931
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__27439\,
            I => n2931
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__27436\,
            I => n2931
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__27429\,
            I => \N__27426\
        );

    \I__3737\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27423\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27420\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__27420\,
            I => \N__27417\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__27417\,
            I => n2998
        );

    \I__3733\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__27411\,
            I => n3097
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__27408\,
            I => \n3030_cascade_\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__27405\,
            I => \N__27401\
        );

    \I__3729\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27397\
        );

    \I__3728\ : InMux
    port map (
            O => \N__27401\,
            I => \N__27394\
        );

    \I__3727\ : InMux
    port map (
            O => \N__27400\,
            I => \N__27391\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__27397\,
            I => n3020
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__27394\,
            I => n3020
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__27391\,
            I => n3020
        );

    \I__3723\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27381\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__27381\,
            I => n3087
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__27378\,
            I => \N__27375\
        );

    \I__3720\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27372\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__27372\,
            I => \N__27368\
        );

    \I__3718\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27364\
        );

    \I__3717\ : Span4Mux_s3_h
    port map (
            O => \N__27368\,
            I => \N__27361\
        );

    \I__3716\ : InMux
    port map (
            O => \N__27367\,
            I => \N__27358\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__27364\,
            I => n2927
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__27361\,
            I => n2927
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__27358\,
            I => n2927
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__27351\,
            I => \N__27348\
        );

    \I__3711\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__3709\ : Span4Mux_h
    port map (
            O => \N__27342\,
            I => \N__27339\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__27339\,
            I => n2994
        );

    \I__3707\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27329\
        );

    \I__3706\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27329\
        );

    \I__3705\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27326\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27323\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27320\
        );

    \I__3702\ : Odrv12
    port map (
            O => \N__27323\,
            I => n2909
        );

    \I__3701\ : Odrv4
    port map (
            O => \N__27320\,
            I => n2909
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__27315\,
            I => \N__27312\
        );

    \I__3699\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27308\
        );

    \I__3698\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27305\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27302\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__27305\,
            I => \N__27299\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__27302\,
            I => \N__27296\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__27299\,
            I => n2907
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__27296\,
            I => n2907
        );

    \I__3692\ : InMux
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__27288\,
            I => n14372
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__27285\,
            I => \N__27280\
        );

    \I__3689\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27275\
        );

    \I__3688\ : InMux
    port map (
            O => \N__27283\,
            I => \N__27275\
        );

    \I__3687\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27272\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__27275\,
            I => \N__27269\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__27272\,
            I => n2929
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__27269\,
            I => n2929
        );

    \I__3683\ : CascadeMux
    port map (
            O => \N__27264\,
            I => \n2940_cascade_\
        );

    \I__3682\ : InMux
    port map (
            O => \N__27261\,
            I => \N__27258\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__27258\,
            I => \N__27255\
        );

    \I__3680\ : Span4Mux_h
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__27252\,
            I => n2996
        );

    \I__3678\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27245\
        );

    \I__3677\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27242\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__27245\,
            I => \N__27239\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27236\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__27239\,
            I => \N__27233\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__27236\,
            I => n2921
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__27233\,
            I => n2921
        );

    \I__3671\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__27225\,
            I => \N__27222\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__27222\,
            I => \N__27219\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__27219\,
            I => n2988
        );

    \I__3667\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__27210\,
            I => n3083
        );

    \I__3664\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__27201\,
            I => n2995
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__27198\,
            I => \N__27194\
        );

    \I__3660\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27190\
        );

    \I__3659\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27187\
        );

    \I__3658\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27184\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__27190\,
            I => n2928
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__27187\,
            I => n2928
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__27184\,
            I => n2928
        );

    \I__3654\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__27171\,
            I => n2997
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__27168\,
            I => \N__27164\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__27167\,
            I => \N__27161\
        );

    \I__3649\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27157\
        );

    \I__3648\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27154\
        );

    \I__3647\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27151\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__27157\,
            I => n2930
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__27154\,
            I => n2930
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__27151\,
            I => n2930
        );

    \I__3643\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__27141\,
            I => n3096
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__27138\,
            I => \n3029_cascade_\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__3639\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27129\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__27126\,
            I => \N__27123\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__27123\,
            I => n2991
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__27120\,
            I => \n2926_cascade_\
        );

    \I__3634\ : InMux
    port map (
            O => \N__27117\,
            I => \N__27114\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__27114\,
            I => n14346
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__27111\,
            I => \n14336_cascade_\
        );

    \I__3631\ : CascadeMux
    port map (
            O => \N__27108\,
            I => \n14352_cascade_\
        );

    \I__3630\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27102\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__27102\,
            I => n14350
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__3627\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27092\
        );

    \I__3626\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27088\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__27092\,
            I => \N__27085\
        );

    \I__3624\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27082\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__27088\,
            I => n2828
        );

    \I__3622\ : Odrv4
    port map (
            O => \N__27085\,
            I => n2828
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__27082\,
            I => n2828
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__27075\,
            I => \N__27072\
        );

    \I__3619\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27069\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__27069\,
            I => \N__27066\
        );

    \I__3617\ : Span4Mux_h
    port map (
            O => \N__27066\,
            I => \N__27063\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__27063\,
            I => n2895
        );

    \I__3615\ : InMux
    port map (
            O => \N__27060\,
            I => \N__27057\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__27057\,
            I => \N__27054\
        );

    \I__3613\ : Span4Mux_v
    port map (
            O => \N__27054\,
            I => \N__27051\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__27051\,
            I => n2885
        );

    \I__3611\ : InMux
    port map (
            O => \N__27048\,
            I => \N__27045\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__27045\,
            I => \N__27041\
        );

    \I__3609\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27038\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__27041\,
            I => \N__27034\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27031\
        );

    \I__3606\ : InMux
    port map (
            O => \N__27037\,
            I => \N__27028\
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__27034\,
            I => n2818
        );

    \I__3604\ : Odrv12
    port map (
            O => \N__27031\,
            I => n2818
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__27028\,
            I => n2818
        );

    \I__3602\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__27015\,
            I => n2881
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__27012\,
            I => \N__27009\
        );

    \I__3598\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27006\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__27006\,
            I => \N__27002\
        );

    \I__3596\ : InMux
    port map (
            O => \N__27005\,
            I => \N__26999\
        );

    \I__3595\ : Span4Mux_h
    port map (
            O => \N__27002\,
            I => \N__26993\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__26999\,
            I => \N__26993\
        );

    \I__3593\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26990\
        );

    \I__3592\ : Odrv4
    port map (
            O => \N__26993\,
            I => n2814
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__26990\,
            I => n2814
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__26985\,
            I => \N__26982\
        );

    \I__3589\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26979\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__26979\,
            I => \N__26976\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__26976\,
            I => \N__26973\
        );

    \I__3586\ : Odrv4
    port map (
            O => \N__26973\,
            I => n12038
        );

    \I__3585\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26967\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__26967\,
            I => n14358
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__26964\,
            I => \n14360_cascade_\
        );

    \I__3582\ : InMux
    port map (
            O => \N__26961\,
            I => \N__26958\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__26958\,
            I => n14366
        );

    \I__3580\ : CascadeMux
    port map (
            O => \N__26955\,
            I => \N__26952\
        );

    \I__3579\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26949\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__26949\,
            I => \N__26946\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__26946\,
            I => \N__26943\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__26943\,
            I => n3094
        );

    \I__3575\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__3573\ : Span4Mux_v
    port map (
            O => \N__26934\,
            I => \N__26931\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__26931\,
            I => n2701
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__26928\,
            I => \N__26924\
        );

    \I__3570\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26921\
        );

    \I__3569\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26918\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__26921\,
            I => \N__26915\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__26918\,
            I => \N__26912\
        );

    \I__3566\ : Span4Mux_s3_h
    port map (
            O => \N__26915\,
            I => \N__26907\
        );

    \I__3565\ : Span4Mux_s3_h
    port map (
            O => \N__26912\,
            I => \N__26907\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__26907\,
            I => n2733
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__26904\,
            I => \n2733_cascade_\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__26901\,
            I => \N__26898\
        );

    \I__3561\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__26895\,
            I => \N__26890\
        );

    \I__3559\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26887\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__26893\,
            I => \N__26884\
        );

    \I__3557\ : Span4Mux_s3_h
    port map (
            O => \N__26890\,
            I => \N__26879\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__26887\,
            I => \N__26879\
        );

    \I__3555\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26876\
        );

    \I__3554\ : Span4Mux_v
    port map (
            O => \N__26879\,
            I => \N__26873\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__26876\,
            I => n2732
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__26873\,
            I => n2732
        );

    \I__3551\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__26865\,
            I => n11936
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__3548\ : InMux
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__26856\,
            I => \N__26852\
        );

    \I__3546\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26849\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__26852\,
            I => \N__26846\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__26849\,
            I => n2729
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__26846\,
            I => n2729
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__26841\,
            I => \N__26838\
        );

    \I__3541\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__26835\,
            I => \N__26832\
        );

    \I__3539\ : Span4Mux_h
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__3538\ : Odrv4
    port map (
            O => \N__26829\,
            I => n2796
        );

    \I__3537\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26823\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__26823\,
            I => \N__26819\
        );

    \I__3535\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26815\
        );

    \I__3534\ : Span4Mux_s2_h
    port map (
            O => \N__26819\,
            I => \N__26812\
        );

    \I__3533\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26809\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__26815\,
            I => n2819
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__26812\,
            I => n2819
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__26809\,
            I => n2819
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__3528\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26796\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__3526\ : Odrv12
    port map (
            O => \N__26793\,
            I => n2886
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__26790\,
            I => \n2918_cascade_\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__26787\,
            I => \N__26784\
        );

    \I__3523\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26780\
        );

    \I__3522\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26776\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__26780\,
            I => \N__26773\
        );

    \I__3520\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26770\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__26776\,
            I => n2827
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__26773\,
            I => n2827
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__26770\,
            I => n2827
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__3515\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26757\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__26757\,
            I => \N__26754\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__26751\,
            I => n2894
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__26748\,
            I => \N__26745\
        );

    \I__3510\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26739\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__26739\,
            I => n2688
        );

    \I__3507\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26732\
        );

    \I__3506\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26729\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26726\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__26729\,
            I => \N__26723\
        );

    \I__3503\ : Odrv4
    port map (
            O => \N__26726\,
            I => n2720
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__26723\,
            I => n2720
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__26718\,
            I => \N__26714\
        );

    \I__3500\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26710\
        );

    \I__3499\ : InMux
    port map (
            O => \N__26714\,
            I => \N__26707\
        );

    \I__3498\ : InMux
    port map (
            O => \N__26713\,
            I => \N__26704\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__26710\,
            I => n2726
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__26707\,
            I => n2726
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__26704\,
            I => n2726
        );

    \I__3494\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26693\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__26696\,
            I => \N__26690\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__26693\,
            I => \N__26686\
        );

    \I__3491\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26683\
        );

    \I__3490\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26680\
        );

    \I__3489\ : Odrv12
    port map (
            O => \N__26686\,
            I => n2724
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__26683\,
            I => n2724
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__26680\,
            I => n2724
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__26673\,
            I => \n2720_cascade_\
        );

    \I__3485\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26666\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__26669\,
            I => \N__26663\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__26666\,
            I => \N__26659\
        );

    \I__3482\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26656\
        );

    \I__3481\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26653\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__26659\,
            I => n2723
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__26656\,
            I => n2723
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__26653\,
            I => n2723
        );

    \I__3477\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__26643\,
            I => n14136
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__26640\,
            I => \N__26637\
        );

    \I__3474\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26634\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__26634\,
            I => \N__26631\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__26631\,
            I => \N__26628\
        );

    \I__3471\ : Odrv4
    port map (
            O => \N__26628\,
            I => n2699
        );

    \I__3470\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26622\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__3468\ : Odrv12
    port map (
            O => \N__26619\,
            I => n2698
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__26616\,
            I => \N__26613\
        );

    \I__3466\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__26610\,
            I => \N__26606\
        );

    \I__3464\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26602\
        );

    \I__3463\ : Span4Mux_s2_h
    port map (
            O => \N__26606\,
            I => \N__26599\
        );

    \I__3462\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26596\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__26602\,
            I => n2820
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__26599\,
            I => n2820
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__26596\,
            I => n2820
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__26589\,
            I => \n14688_cascade_\
        );

    \I__3457\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26583\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__3455\ : Odrv4
    port map (
            O => \N__26580\,
            I => n14690
        );

    \I__3454\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__26574\,
            I => \N__26571\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__26571\,
            I => n14696
        );

    \I__3451\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26565\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__26565\,
            I => \N__26562\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__26562\,
            I => \N__26559\
        );

    \I__3448\ : Span4Mux_h
    port map (
            O => \N__26559\,
            I => \N__26556\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__26556\,
            I => \N__26553\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__26553\,
            I => \ENCODER0_B_N\
        );

    \I__3445\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26547\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__26547\,
            I => \N__26544\
        );

    \I__3443\ : Odrv12
    port map (
            O => \N__26544\,
            I => n2697
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__26541\,
            I => \N__26538\
        );

    \I__3441\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26534\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__26537\,
            I => \N__26531\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__26534\,
            I => \N__26527\
        );

    \I__3438\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26524\
        );

    \I__3437\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26521\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__26527\,
            I => n2630
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__26524\,
            I => n2630
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__26521\,
            I => n2630
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__26514\,
            I => \N__26510\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__26513\,
            I => \N__26507\
        );

    \I__3431\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26504\
        );

    \I__3430\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26501\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__26504\,
            I => \N__26498\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26494\
        );

    \I__3427\ : Span4Mux_s1_h
    port map (
            O => \N__26498\,
            I => \N__26491\
        );

    \I__3426\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26488\
        );

    \I__3425\ : Span4Mux_s3_h
    port map (
            O => \N__26494\,
            I => \N__26485\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__26491\,
            I => n2731
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__26488\,
            I => n2731
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__26485\,
            I => n2731
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__26478\,
            I => \N__26475\
        );

    \I__3420\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26471\
        );

    \I__3419\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26468\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__26471\,
            I => \N__26464\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26461\
        );

    \I__3416\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26458\
        );

    \I__3415\ : Span4Mux_s3_h
    port map (
            O => \N__26464\,
            I => \N__26455\
        );

    \I__3414\ : Odrv12
    port map (
            O => \N__26461\,
            I => n2730
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__26458\,
            I => n2730
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__26455\,
            I => n2730
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__26448\,
            I => \n2729_cascade_\
        );

    \I__3410\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26442\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__26442\,
            I => n13796
        );

    \I__3408\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26436\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__26436\,
            I => \N__26432\
        );

    \I__3406\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26429\
        );

    \I__3405\ : Odrv12
    port map (
            O => \N__26432\,
            I => n2613
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__26429\,
            I => n2613
        );

    \I__3403\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26421\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__26421\,
            I => \N__26418\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__26418\,
            I => n2680
        );

    \I__3400\ : InMux
    port map (
            O => \N__26415\,
            I => n12768
        );

    \I__3399\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26409\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__26409\,
            I => \N__26405\
        );

    \I__3397\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26402\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__26405\,
            I => \N__26399\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__26402\,
            I => \N__26396\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__26399\,
            I => n2612
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__26396\,
            I => n2612
        );

    \I__3392\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26388\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26385\
        );

    \I__3390\ : Span4Mux_s3_h
    port map (
            O => \N__26385\,
            I => \N__26382\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__26382\,
            I => n2679
        );

    \I__3388\ : InMux
    port map (
            O => \N__26379\,
            I => n12769
        );

    \I__3387\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26372\
        );

    \I__3386\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26369\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26365\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__26369\,
            I => \N__26362\
        );

    \I__3383\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26359\
        );

    \I__3382\ : Span4Mux_h
    port map (
            O => \N__26365\,
            I => \N__26356\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__26362\,
            I => \N__26351\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26351\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__26356\,
            I => n2611
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__26351\,
            I => n2611
        );

    \I__3377\ : CascadeMux
    port map (
            O => \N__26346\,
            I => \N__26343\
        );

    \I__3376\ : InMux
    port map (
            O => \N__26343\,
            I => \N__26340\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__26340\,
            I => \N__26337\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__26337\,
            I => \N__26334\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__26334\,
            I => n2678
        );

    \I__3372\ : InMux
    port map (
            O => \N__26331\,
            I => n12770
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__26328\,
            I => \N__26325\
        );

    \I__3370\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26322\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__26322\,
            I => \N__26318\
        );

    \I__3368\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26315\
        );

    \I__3367\ : Span4Mux_h
    port map (
            O => \N__26318\,
            I => \N__26312\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__26315\,
            I => \N__26309\
        );

    \I__3365\ : Span4Mux_s0_h
    port map (
            O => \N__26312\,
            I => \N__26304\
        );

    \I__3364\ : Span4Mux_h
    port map (
            O => \N__26309\,
            I => \N__26304\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__26304\,
            I => n2610
        );

    \I__3362\ : InMux
    port map (
            O => \N__26301\,
            I => \bfn_4_24_0_\
        );

    \I__3361\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26292\
        );

    \I__3360\ : InMux
    port map (
            O => \N__26297\,
            I => \N__26292\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__26292\,
            I => \N__26289\
        );

    \I__3358\ : Span4Mux_s3_h
    port map (
            O => \N__26289\,
            I => \N__26286\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__26286\,
            I => n2709
        );

    \I__3356\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26279\
        );

    \I__3355\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26276\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__26279\,
            I => \N__26273\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__26276\,
            I => \N__26270\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__26273\,
            I => n2816
        );

    \I__3351\ : Odrv12
    port map (
            O => \N__26270\,
            I => n2816
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__26265\,
            I => \N__26262\
        );

    \I__3349\ : InMux
    port map (
            O => \N__26262\,
            I => \N__26259\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__26259\,
            I => \N__26256\
        );

    \I__3347\ : Span4Mux_h
    port map (
            O => \N__26256\,
            I => \N__26253\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__26253\,
            I => n2883
        );

    \I__3345\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26246\
        );

    \I__3344\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26243\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__26246\,
            I => \N__26237\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__26243\,
            I => \N__26237\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__26242\,
            I => \N__26234\
        );

    \I__3340\ : Span4Mux_v
    port map (
            O => \N__26237\,
            I => \N__26231\
        );

    \I__3339\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26228\
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__26231\,
            I => n2621
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__26228\,
            I => n2621
        );

    \I__3336\ : InMux
    port map (
            O => \N__26223\,
            I => n12760
        );

    \I__3335\ : InMux
    port map (
            O => \N__26220\,
            I => \N__26216\
        );

    \I__3334\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26212\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__26216\,
            I => \N__26209\
        );

    \I__3332\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26206\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__26212\,
            I => n2620
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__26209\,
            I => n2620
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__26206\,
            I => n2620
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__26199\,
            I => \N__26196\
        );

    \I__3327\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26193\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__26193\,
            I => \N__26190\
        );

    \I__3325\ : Span4Mux_s3_h
    port map (
            O => \N__26190\,
            I => \N__26187\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__26187\,
            I => n2687
        );

    \I__3323\ : InMux
    port map (
            O => \N__26184\,
            I => n12761
        );

    \I__3322\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26178\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__26178\,
            I => \N__26174\
        );

    \I__3320\ : InMux
    port map (
            O => \N__26177\,
            I => \N__26170\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__26174\,
            I => \N__26167\
        );

    \I__3318\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26164\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__26170\,
            I => n2619
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__26167\,
            I => n2619
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__26164\,
            I => n2619
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__26157\,
            I => \N__26154\
        );

    \I__3313\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26151\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__26151\,
            I => n2686
        );

    \I__3311\ : InMux
    port map (
            O => \N__26148\,
            I => n12762
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__26145\,
            I => \N__26142\
        );

    \I__3309\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26139\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__26139\,
            I => \N__26135\
        );

    \I__3307\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26132\
        );

    \I__3306\ : Span4Mux_v
    port map (
            O => \N__26135\,
            I => \N__26129\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26126\
        );

    \I__3304\ : Span4Mux_s2_h
    port map (
            O => \N__26129\,
            I => \N__26122\
        );

    \I__3303\ : Span4Mux_v
    port map (
            O => \N__26126\,
            I => \N__26119\
        );

    \I__3302\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26116\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__26122\,
            I => n2618
        );

    \I__3300\ : Odrv4
    port map (
            O => \N__26119\,
            I => n2618
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__26116\,
            I => n2618
        );

    \I__3298\ : InMux
    port map (
            O => \N__26109\,
            I => \N__26106\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__26106\,
            I => n2685
        );

    \I__3296\ : InMux
    port map (
            O => \N__26103\,
            I => \bfn_4_23_0_\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__26100\,
            I => \N__26096\
        );

    \I__3294\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26093\
        );

    \I__3293\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26090\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__26093\,
            I => n2617
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__26090\,
            I => n2617
        );

    \I__3290\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26082\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__26082\,
            I => n2684
        );

    \I__3288\ : InMux
    port map (
            O => \N__26079\,
            I => n12764
        );

    \I__3287\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26071\
        );

    \I__3286\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26068\
        );

    \I__3285\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26065\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__26071\,
            I => \N__26060\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__26068\,
            I => \N__26060\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__26065\,
            I => n2616
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__26060\,
            I => n2616
        );

    \I__3280\ : InMux
    port map (
            O => \N__26055\,
            I => \N__26052\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__26052\,
            I => \N__26049\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__26049\,
            I => n2683
        );

    \I__3277\ : InMux
    port map (
            O => \N__26046\,
            I => n12765
        );

    \I__3276\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26040\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__26040\,
            I => \N__26036\
        );

    \I__3274\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26033\
        );

    \I__3273\ : Span4Mux_s3_h
    port map (
            O => \N__26036\,
            I => \N__26027\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__26033\,
            I => \N__26027\
        );

    \I__3271\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26024\
        );

    \I__3270\ : Span4Mux_v
    port map (
            O => \N__26027\,
            I => \N__26021\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__26024\,
            I => \N__26018\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__26021\,
            I => n2615
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__26018\,
            I => n2615
        );

    \I__3266\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26010\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__26010\,
            I => \N__26007\
        );

    \I__3264\ : Span4Mux_s3_h
    port map (
            O => \N__26007\,
            I => \N__26004\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__26004\,
            I => n2682
        );

    \I__3262\ : InMux
    port map (
            O => \N__26001\,
            I => n12766
        );

    \I__3261\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25991\
        );

    \I__3260\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25991\
        );

    \I__3259\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25988\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25985\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__25988\,
            I => n2614
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__25985\,
            I => n2614
        );

    \I__3255\ : InMux
    port map (
            O => \N__25980\,
            I => \N__25977\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__25977\,
            I => n2681
        );

    \I__3253\ : InMux
    port map (
            O => \N__25974\,
            I => n12767
        );

    \I__3252\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25967\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__25970\,
            I => \N__25964\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__25967\,
            I => \N__25961\
        );

    \I__3249\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25958\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__25961\,
            I => n2629
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__25958\,
            I => n2629
        );

    \I__3246\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25950\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25947\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__25947\,
            I => n2696
        );

    \I__3243\ : InMux
    port map (
            O => \N__25944\,
            I => n12752
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__25941\,
            I => \N__25937\
        );

    \I__3241\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25934\
        );

    \I__3240\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25931\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__25934\,
            I => \N__25928\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__25931\,
            I => \N__25925\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__25928\,
            I => n2628
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__25925\,
            I => n2628
        );

    \I__3235\ : InMux
    port map (
            O => \N__25920\,
            I => \N__25917\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__25917\,
            I => \N__25914\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__25914\,
            I => n2695
        );

    \I__3232\ : InMux
    port map (
            O => \N__25911\,
            I => n12753
        );

    \I__3231\ : InMux
    port map (
            O => \N__25908\,
            I => \N__25905\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__25905\,
            I => \N__25901\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__25904\,
            I => \N__25898\
        );

    \I__3228\ : Span4Mux_h
    port map (
            O => \N__25901\,
            I => \N__25895\
        );

    \I__3227\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25892\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__25895\,
            I => \N__25887\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__25892\,
            I => \N__25887\
        );

    \I__3224\ : Odrv4
    port map (
            O => \N__25887\,
            I => n2627
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__25884\,
            I => \N__25881\
        );

    \I__3222\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25878\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__25878\,
            I => \N__25875\
        );

    \I__3220\ : Span4Mux_v
    port map (
            O => \N__25875\,
            I => \N__25872\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__25872\,
            I => n2694
        );

    \I__3218\ : InMux
    port map (
            O => \N__25869\,
            I => n12754
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__25866\,
            I => \N__25862\
        );

    \I__3216\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25859\
        );

    \I__3215\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25855\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__25859\,
            I => \N__25852\
        );

    \I__3213\ : InMux
    port map (
            O => \N__25858\,
            I => \N__25849\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__25855\,
            I => n2626
        );

    \I__3211\ : Odrv12
    port map (
            O => \N__25852\,
            I => n2626
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__25849\,
            I => n2626
        );

    \I__3209\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25839\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__25839\,
            I => n2693
        );

    \I__3207\ : InMux
    port map (
            O => \N__25836\,
            I => \bfn_4_22_0_\
        );

    \I__3206\ : InMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__25830\,
            I => \N__25825\
        );

    \I__3204\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25822\
        );

    \I__3203\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25819\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__25825\,
            I => n2625
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__25822\,
            I => n2625
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__25819\,
            I => n2625
        );

    \I__3199\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__25809\,
            I => n2692
        );

    \I__3197\ : InMux
    port map (
            O => \N__25806\,
            I => n12756
        );

    \I__3196\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__25800\,
            I => \N__25797\
        );

    \I__3194\ : Span4Mux_h
    port map (
            O => \N__25797\,
            I => \N__25793\
        );

    \I__3193\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25790\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__25793\,
            I => n2624
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__25790\,
            I => n2624
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__25785\,
            I => \N__25782\
        );

    \I__3189\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__25779\,
            I => \N__25776\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__25776\,
            I => n2691
        );

    \I__3186\ : InMux
    port map (
            O => \N__25773\,
            I => n12757
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__25770\,
            I => \N__25767\
        );

    \I__3184\ : InMux
    port map (
            O => \N__25767\,
            I => \N__25764\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__25764\,
            I => \N__25759\
        );

    \I__3182\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25756\
        );

    \I__3181\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25753\
        );

    \I__3180\ : Odrv12
    port map (
            O => \N__25759\,
            I => n2623
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__25756\,
            I => n2623
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__25753\,
            I => n2623
        );

    \I__3177\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25743\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__25743\,
            I => \N__25740\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__25740\,
            I => n2690
        );

    \I__3174\ : InMux
    port map (
            O => \N__25737\,
            I => n12758
        );

    \I__3173\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25731\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__25731\,
            I => \N__25726\
        );

    \I__3171\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25723\
        );

    \I__3170\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25720\
        );

    \I__3169\ : Odrv12
    port map (
            O => \N__25726\,
            I => n2622
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__25723\,
            I => n2622
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__25720\,
            I => n2622
        );

    \I__3166\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25710\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__25710\,
            I => \N__25707\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__25707\,
            I => n2689
        );

    \I__3163\ : InMux
    port map (
            O => \N__25704\,
            I => n12759
        );

    \I__3162\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__25698\,
            I => \N__25695\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__25695\,
            I => \N__25692\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__25692\,
            I => n2492
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__25689\,
            I => \N__25686\
        );

    \I__3157\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25682\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__25685\,
            I => \N__25679\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__25682\,
            I => \N__25676\
        );

    \I__3154\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25673\
        );

    \I__3153\ : Span4Mux_v
    port map (
            O => \N__25676\,
            I => \N__25670\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__25673\,
            I => n2425
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__25670\,
            I => n2425
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__25665\,
            I => \N__25662\
        );

    \I__3149\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25659\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__25659\,
            I => \N__25656\
        );

    \I__3147\ : Span4Mux_v
    port map (
            O => \N__25656\,
            I => \N__25651\
        );

    \I__3146\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25646\
        );

    \I__3145\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25646\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__25651\,
            I => n2524
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__25646\,
            I => n2524
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__3141\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25633\
        );

    \I__3140\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25628\
        );

    \I__3139\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25628\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__25633\,
            I => n2318
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__25628\,
            I => n2318
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__25623\,
            I => \N__25620\
        );

    \I__3135\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25616\
        );

    \I__3134\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25612\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__25616\,
            I => \N__25609\
        );

    \I__3132\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25606\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__25612\,
            I => n2320
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__25609\,
            I => n2320
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__25606\,
            I => n2320
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__3127\ : InMux
    port map (
            O => \N__25596\,
            I => \N__25593\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__25593\,
            I => \N__25589\
        );

    \I__3125\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25586\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__25589\,
            I => \N__25582\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__25586\,
            I => \N__25579\
        );

    \I__3122\ : InMux
    port map (
            O => \N__25585\,
            I => \N__25576\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__25582\,
            I => n2319
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__25579\,
            I => n2319
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__25576\,
            I => n2319
        );

    \I__3118\ : InMux
    port map (
            O => \N__25569\,
            I => \bfn_4_21_0_\
        );

    \I__3117\ : InMux
    port map (
            O => \N__25566\,
            I => \N__25563\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__25563\,
            I => \N__25560\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__25560\,
            I => n2700
        );

    \I__3114\ : InMux
    port map (
            O => \N__25557\,
            I => n12748
        );

    \I__3113\ : InMux
    port map (
            O => \N__25554\,
            I => n12749
        );

    \I__3112\ : InMux
    port map (
            O => \N__25551\,
            I => n12750
        );

    \I__3111\ : InMux
    port map (
            O => \N__25548\,
            I => n12751
        );

    \I__3110\ : InMux
    port map (
            O => \N__25545\,
            I => n12699
        );

    \I__3109\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25539\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__25539\,
            I => n2382
        );

    \I__3107\ : InMux
    port map (
            O => \N__25536\,
            I => n12700
        );

    \I__3106\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__25530\,
            I => n2381
        );

    \I__3104\ : InMux
    port map (
            O => \N__25527\,
            I => n12701
        );

    \I__3103\ : InMux
    port map (
            O => \N__25524\,
            I => n12702
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__25521\,
            I => \N__25518\
        );

    \I__3101\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__25515\,
            I => \N__25511\
        );

    \I__3099\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25508\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__25511\,
            I => n2412
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__25508\,
            I => n2412
        );

    \I__3096\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25498\
        );

    \I__3095\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25495\
        );

    \I__3094\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25492\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__25498\,
            I => n2314_adj_622
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__25495\,
            I => n2314_adj_622
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__25492\,
            I => n2314_adj_622
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__25485\,
            I => \N__25481\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__25484\,
            I => \N__25478\
        );

    \I__3088\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25475\
        );

    \I__3087\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25472\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__25475\,
            I => \N__25467\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__25472\,
            I => \N__25467\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__25467\,
            I => n2327
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__25464\,
            I => \n2327_cascade_\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__25461\,
            I => \N__25457\
        );

    \I__3081\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25453\
        );

    \I__3080\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25450\
        );

    \I__3079\ : InMux
    port map (
            O => \N__25456\,
            I => \N__25447\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__25453\,
            I => n2326
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__25450\,
            I => n2326
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__25447\,
            I => n2326
        );

    \I__3075\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__25437\,
            I => n14440
        );

    \I__3073\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__25431\,
            I => n2391
        );

    \I__3071\ : InMux
    port map (
            O => \N__25428\,
            I => n12691
        );

    \I__3070\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__25419\,
            I => n2390
        );

    \I__3067\ : InMux
    port map (
            O => \N__25416\,
            I => n12692
        );

    \I__3066\ : InMux
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__25410\,
            I => n2389
        );

    \I__3064\ : InMux
    port map (
            O => \N__25407\,
            I => n12693
        );

    \I__3063\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__25401\,
            I => n2388
        );

    \I__3061\ : InMux
    port map (
            O => \N__25398\,
            I => n12694
        );

    \I__3060\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__25392\,
            I => n2387
        );

    \I__3058\ : InMux
    port map (
            O => \N__25389\,
            I => n12695
        );

    \I__3057\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__25383\,
            I => \N__25380\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__25380\,
            I => n2386
        );

    \I__3054\ : InMux
    port map (
            O => \N__25377\,
            I => n12696
        );

    \I__3053\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__25371\,
            I => n2385
        );

    \I__3051\ : InMux
    port map (
            O => \N__25368\,
            I => \bfn_4_19_0_\
        );

    \I__3050\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__25359\,
            I => n2384
        );

    \I__3047\ : InMux
    port map (
            O => \N__25356\,
            I => n12698
        );

    \I__3046\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25350\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__25350\,
            I => n2383
        );

    \I__3044\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25344\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__25344\,
            I => \N__25341\
        );

    \I__3042\ : Span4Mux_s3_h
    port map (
            O => \N__25341\,
            I => \N__25338\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__25338\,
            I => n2399
        );

    \I__3040\ : InMux
    port map (
            O => \N__25335\,
            I => n12683
        );

    \I__3039\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25329\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__25329\,
            I => \N__25326\
        );

    \I__3037\ : Span4Mux_s3_h
    port map (
            O => \N__25326\,
            I => \N__25323\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__25323\,
            I => n2398
        );

    \I__3035\ : InMux
    port map (
            O => \N__25320\,
            I => n12684
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__25317\,
            I => \N__25314\
        );

    \I__3033\ : InMux
    port map (
            O => \N__25314\,
            I => \N__25311\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__25311\,
            I => n2397
        );

    \I__3031\ : InMux
    port map (
            O => \N__25308\,
            I => n12685
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__25305\,
            I => \N__25301\
        );

    \I__3029\ : CascadeMux
    port map (
            O => \N__25304\,
            I => \N__25298\
        );

    \I__3028\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25294\
        );

    \I__3027\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25291\
        );

    \I__3026\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25288\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__25294\,
            I => \N__25285\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__25291\,
            I => n2329
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__25288\,
            I => n2329
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__25285\,
            I => n2329
        );

    \I__3021\ : InMux
    port map (
            O => \N__25278\,
            I => \N__25275\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__25275\,
            I => \N__25272\
        );

    \I__3019\ : Span4Mux_s3_h
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__25269\,
            I => n2396
        );

    \I__3017\ : InMux
    port map (
            O => \N__25266\,
            I => n12686
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__25263\,
            I => \N__25259\
        );

    \I__3015\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25256\
        );

    \I__3014\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25253\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__25256\,
            I => \N__25248\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25248\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__25248\,
            I => n2328
        );

    \I__3010\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__25242\,
            I => n2395
        );

    \I__3008\ : InMux
    port map (
            O => \N__25239\,
            I => n12687
        );

    \I__3007\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25233\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__25233\,
            I => n2394
        );

    \I__3005\ : InMux
    port map (
            O => \N__25230\,
            I => n12688
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__25227\,
            I => \N__25224\
        );

    \I__3003\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__25221\,
            I => n2393
        );

    \I__3001\ : InMux
    port map (
            O => \N__25218\,
            I => \bfn_4_18_0_\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__25215\,
            I => \N__25212\
        );

    \I__2999\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25209\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__25209\,
            I => \N__25206\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__25206\,
            I => n2392
        );

    \I__2996\ : InMux
    port map (
            O => \N__25203\,
            I => n12690
        );

    \I__2995\ : InMux
    port map (
            O => \N__25200\,
            I => \bfn_3_32_0_\
        );

    \I__2994\ : InMux
    port map (
            O => \N__25197\,
            I => n12874
        );

    \I__2993\ : InMux
    port map (
            O => \N__25194\,
            I => n12875
        );

    \I__2992\ : InMux
    port map (
            O => \N__25191\,
            I => n12876
        );

    \I__2991\ : InMux
    port map (
            O => \N__25188\,
            I => n12877
        );

    \I__2990\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__25182\,
            I => \N__25178\
        );

    \I__2988\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25175\
        );

    \I__2987\ : Span4Mux_s1_v
    port map (
            O => \N__25178\,
            I => \N__25172\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__25175\,
            I => \debounce.cnt_reg_6\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__25172\,
            I => \debounce.cnt_reg_6\
        );

    \I__2984\ : InMux
    port map (
            O => \N__25167\,
            I => \N__25164\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__25164\,
            I => \debounce.n16\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__2981\ : InMux
    port map (
            O => \N__25158\,
            I => \N__25155\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__25155\,
            I => \N__25151\
        );

    \I__2979\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25148\
        );

    \I__2978\ : Span4Mux_s1_v
    port map (
            O => \N__25151\,
            I => \N__25145\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__25148\,
            I => \debounce.cnt_reg_3\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__25145\,
            I => \debounce.cnt_reg_3\
        );

    \I__2975\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25137\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__25137\,
            I => \debounce.n17\
        );

    \I__2973\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25131\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__2971\ : Odrv4
    port map (
            O => \N__25128\,
            I => n2401
        );

    \I__2970\ : InMux
    port map (
            O => \N__25125\,
            I => \bfn_4_17_0_\
        );

    \I__2969\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25119\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__25119\,
            I => \N__25116\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__25116\,
            I => n2400
        );

    \I__2966\ : InMux
    port map (
            O => \N__25113\,
            I => n12682
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__25110\,
            I => \N__25107\
        );

    \I__2964\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__25104\,
            I => \N__25101\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__25101\,
            I => n3086
        );

    \I__2961\ : InMux
    port map (
            O => \N__25098\,
            I => n12864
        );

    \I__2960\ : InMux
    port map (
            O => \N__25095\,
            I => \bfn_3_31_0_\
        );

    \I__2959\ : InMux
    port map (
            O => \N__25092\,
            I => n12866
        );

    \I__2958\ : InMux
    port map (
            O => \N__25089\,
            I => n12867
        );

    \I__2957\ : InMux
    port map (
            O => \N__25086\,
            I => n12868
        );

    \I__2956\ : InMux
    port map (
            O => \N__25083\,
            I => n12869
        );

    \I__2955\ : InMux
    port map (
            O => \N__25080\,
            I => n12870
        );

    \I__2954\ : InMux
    port map (
            O => \N__25077\,
            I => n12871
        );

    \I__2953\ : InMux
    port map (
            O => \N__25074\,
            I => n12872
        );

    \I__2952\ : InMux
    port map (
            O => \N__25071\,
            I => n12855
        );

    \I__2951\ : InMux
    port map (
            O => \N__25068\,
            I => n12856
        );

    \I__2950\ : InMux
    port map (
            O => \N__25065\,
            I => \bfn_3_30_0_\
        );

    \I__2949\ : InMux
    port map (
            O => \N__25062\,
            I => n12858
        );

    \I__2948\ : InMux
    port map (
            O => \N__25059\,
            I => n12859
        );

    \I__2947\ : InMux
    port map (
            O => \N__25056\,
            I => n12860
        );

    \I__2946\ : InMux
    port map (
            O => \N__25053\,
            I => n12861
        );

    \I__2945\ : InMux
    port map (
            O => \N__25050\,
            I => n12862
        );

    \I__2944\ : InMux
    port map (
            O => \N__25047\,
            I => n12863
        );

    \I__2943\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__2941\ : Span4Mux_h
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__2940\ : Odrv4
    port map (
            O => \N__25035\,
            I => n2893
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__25032\,
            I => \N__25028\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__25031\,
            I => \N__25025\
        );

    \I__2937\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25021\
        );

    \I__2936\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25018\
        );

    \I__2935\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25015\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__25021\,
            I => n2826
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__25018\,
            I => n2826
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__25015\,
            I => n2826
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__2930\ : InMux
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__24999\,
            I => n2882
        );

    \I__2927\ : InMux
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__24993\,
            I => \N__24989\
        );

    \I__2925\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24986\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__24989\,
            I => \N__24980\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__24986\,
            I => \N__24980\
        );

    \I__2922\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24977\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__24980\,
            I => n2815
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__24977\,
            I => n2815
        );

    \I__2919\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24967\
        );

    \I__2918\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24964\
        );

    \I__2917\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24961\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__24967\,
            I => n2813
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__24964\,
            I => n2813
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__24961\,
            I => n2813
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__24954\,
            I => \N__24951\
        );

    \I__2912\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__2910\ : Span4Mux_h
    port map (
            O => \N__24945\,
            I => \N__24942\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__24942\,
            I => n2880
        );

    \I__2908\ : InMux
    port map (
            O => \N__24939\,
            I => \bfn_3_29_0_\
        );

    \I__2907\ : InMux
    port map (
            O => \N__24936\,
            I => n12850
        );

    \I__2906\ : InMux
    port map (
            O => \N__24933\,
            I => n12851
        );

    \I__2905\ : InMux
    port map (
            O => \N__24930\,
            I => n12852
        );

    \I__2904\ : InMux
    port map (
            O => \N__24927\,
            I => n12853
        );

    \I__2903\ : InMux
    port map (
            O => \N__24924\,
            I => n12854
        );

    \I__2902\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24918\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__24918\,
            I => n2777
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__24915\,
            I => \N__24912\
        );

    \I__2899\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24907\
        );

    \I__2898\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24902\
        );

    \I__2897\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24902\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__24907\,
            I => n2710
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__24902\,
            I => n2710
        );

    \I__2894\ : InMux
    port map (
            O => \N__24897\,
            I => \N__24893\
        );

    \I__2893\ : InMux
    port map (
            O => \N__24896\,
            I => \N__24890\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__24893\,
            I => \N__24887\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__24890\,
            I => \N__24884\
        );

    \I__2890\ : Span4Mux_v
    port map (
            O => \N__24887\,
            I => \N__24881\
        );

    \I__2889\ : Span4Mux_s2_h
    port map (
            O => \N__24884\,
            I => \N__24878\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__24881\,
            I => n2809
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__24878\,
            I => n2809
        );

    \I__2886\ : InMux
    port map (
            O => \N__24873\,
            I => \N__24868\
        );

    \I__2885\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24865\
        );

    \I__2884\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24862\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__24868\,
            I => \N__24857\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__24865\,
            I => \N__24857\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__24862\,
            I => \N__24854\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__24857\,
            I => n2810
        );

    \I__2879\ : Odrv4
    port map (
            O => \N__24854\,
            I => n2810
        );

    \I__2878\ : InMux
    port map (
            O => \N__24849\,
            I => \N__24846\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__2876\ : Span4Mux_v
    port map (
            O => \N__24843\,
            I => \N__24839\
        );

    \I__2875\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24836\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__24839\,
            I => n2808
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__24836\,
            I => n2808
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__24831\,
            I => \n2809_cascade_\
        );

    \I__2871\ : InMux
    port map (
            O => \N__24828\,
            I => \N__24825\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__24825\,
            I => n14714
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__24822\,
            I => \N__24819\
        );

    \I__2868\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24815\
        );

    \I__2867\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24812\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24809\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__24812\,
            I => n2823
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__24809\,
            I => n2823
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__24804\,
            I => \n2841_cascade_\
        );

    \I__2862\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__24798\,
            I => \N__24795\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__24795\,
            I => n2890
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__2858\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24785\
        );

    \I__2857\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24781\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__24785\,
            I => \N__24778\
        );

    \I__2855\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24775\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__24781\,
            I => n2920
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__24778\,
            I => n2920
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__24775\,
            I => n2920
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__24768\,
            I => \N__24765\
        );

    \I__2850\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24762\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24759\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__24759\,
            I => n2987
        );

    \I__2847\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24753\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__2845\ : Span4Mux_v
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__24747\,
            I => n2898
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__24744\,
            I => \N__24741\
        );

    \I__2842\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24738\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__24738\,
            I => \N__24734\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__24737\,
            I => \N__24731\
        );

    \I__2839\ : Span4Mux_h
    port map (
            O => \N__24734\,
            I => \N__24727\
        );

    \I__2838\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24724\
        );

    \I__2837\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24721\
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__24727\,
            I => n2831
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__24724\,
            I => n2831
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__24721\,
            I => n2831
        );

    \I__2833\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24711\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__24708\,
            I => n2879
        );

    \I__2830\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24700\
        );

    \I__2829\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24697\
        );

    \I__2828\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24694\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__24700\,
            I => n2812
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__24697\,
            I => n2812
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__24694\,
            I => n2812
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__24687\,
            I => \n2911_cascade_\
        );

    \I__2823\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24681\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__24681\,
            I => \N__24677\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__24677\,
            I => \N__24671\
        );

    \I__2819\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24668\
        );

    \I__2818\ : Odrv4
    port map (
            O => \N__24671\,
            I => n2829
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__24668\,
            I => n2829
        );

    \I__2816\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24660\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__24660\,
            I => \N__24657\
        );

    \I__2814\ : Span4Mux_h
    port map (
            O => \N__24657\,
            I => \N__24654\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__24654\,
            I => n2896
        );

    \I__2812\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24646\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__24650\,
            I => \N__24643\
        );

    \I__2810\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24640\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24637\
        );

    \I__2808\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24634\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24631\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__24637\,
            I => n2725
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__24634\,
            I => n2725
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__24631\,
            I => n2725
        );

    \I__2803\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24621\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__24621\,
            I => \N__24618\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__24618\,
            I => \N__24615\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__24615\,
            I => n2792
        );

    \I__2799\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24608\
        );

    \I__2798\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24605\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__24608\,
            I => n2721
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__24605\,
            I => n2721
        );

    \I__2795\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24597\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__24597\,
            I => \N__24594\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__24594\,
            I => n2788
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__24591\,
            I => \N__24588\
        );

    \I__2791\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24585\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24582\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__24582\,
            I => n2793
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__24579\,
            I => \N__24576\
        );

    \I__2787\ : InMux
    port map (
            O => \N__24576\,
            I => \N__24573\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__24573\,
            I => \N__24570\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__24570\,
            I => n2889
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__24567\,
            I => \n2921_cascade_\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__24564\,
            I => \N__24561\
        );

    \I__2782\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24558\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__24555\,
            I => n2888
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__24552\,
            I => \N__24549\
        );

    \I__2778\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24546\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__24546\,
            I => \N__24543\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__24543\,
            I => n2791
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__2774\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24532\
        );

    \I__2773\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24527\
        );

    \I__2772\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24527\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__24532\,
            I => n2822
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__24527\,
            I => n2822
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__24522\,
            I => \n2823_cascade_\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__24519\,
            I => \N__24516\
        );

    \I__2767\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24511\
        );

    \I__2766\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24506\
        );

    \I__2765\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24506\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__24511\,
            I => n2821
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__24506\,
            I => n2821
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__24501\,
            I => \n2721_cascade_\
        );

    \I__2761\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__24495\,
            I => \N__24490\
        );

    \I__2759\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24487\
        );

    \I__2758\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24484\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__24490\,
            I => n2717
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__24487\,
            I => n2717
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__24484\,
            I => n2717
        );

    \I__2754\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24473\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__24476\,
            I => \N__24470\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__24473\,
            I => \N__24466\
        );

    \I__2751\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24463\
        );

    \I__2750\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24460\
        );

    \I__2749\ : Span4Mux_s2_h
    port map (
            O => \N__24466\,
            I => \N__24453\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__24463\,
            I => \N__24453\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__24460\,
            I => \N__24453\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__24453\,
            I => n2718
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__24450\,
            I => \n14140_cascade_\
        );

    \I__2744\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24444\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24441\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__24441\,
            I => \N__24438\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__24438\,
            I => n14138
        );

    \I__2740\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24431\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__24434\,
            I => \N__24428\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__24431\,
            I => \N__24424\
        );

    \I__2737\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24421\
        );

    \I__2736\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24418\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__24424\,
            I => \N__24415\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__24421\,
            I => \N__24410\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__24418\,
            I => \N__24410\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__24415\,
            I => n2716
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__24410\,
            I => n2716
        );

    \I__2730\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__24402\,
            I => \N__24397\
        );

    \I__2728\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24394\
        );

    \I__2727\ : InMux
    port map (
            O => \N__24400\,
            I => \N__24391\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__24397\,
            I => n2715
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__24394\,
            I => n2715
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__24391\,
            I => n2715
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__24384\,
            I => \n14146_cascade_\
        );

    \I__2722\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24378\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__24378\,
            I => n14152
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__24375\,
            I => \N__24371\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__24374\,
            I => \N__24368\
        );

    \I__2718\ : InMux
    port map (
            O => \N__24371\,
            I => \N__24364\
        );

    \I__2717\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24361\
        );

    \I__2716\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24358\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__24364\,
            I => n2722
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__24361\,
            I => n2722
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__24358\,
            I => n2722
        );

    \I__2712\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24348\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__24345\,
            I => n2787
        );

    \I__2709\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24339\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__24339\,
            I => \N__24336\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__24336\,
            I => n2795
        );

    \I__2706\ : InMux
    port map (
            O => \N__24333\,
            I => \N__24330\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__24330\,
            I => \N__24325\
        );

    \I__2704\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24322\
        );

    \I__2703\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24319\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__24325\,
            I => n2728
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__24322\,
            I => n2728
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__24319\,
            I => n2728
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__24312\,
            I => \N__24307\
        );

    \I__2698\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24304\
        );

    \I__2697\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24301\
        );

    \I__2696\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24298\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__24304\,
            I => n2712
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__24301\,
            I => n2712
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__24298\,
            I => n2712
        );

    \I__2692\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24288\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__24288\,
            I => \N__24284\
        );

    \I__2690\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24281\
        );

    \I__2689\ : Span4Mux_v
    port map (
            O => \N__24284\,
            I => \N__24277\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__24281\,
            I => \N__24274\
        );

    \I__2687\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24271\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__24277\,
            I => n2514
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__24274\,
            I => n2514
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__24271\,
            I => n2514
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__24264\,
            I => \N__24261\
        );

    \I__2682\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24258\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__24258\,
            I => \N__24255\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__24255\,
            I => \N__24252\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__24252\,
            I => n2581
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__24249\,
            I => \n2613_cascade_\
        );

    \I__2677\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__24243\,
            I => n14664
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__24240\,
            I => \n14670_cascade_\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__24237\,
            I => \n2643_cascade_\
        );

    \I__2673\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24229\
        );

    \I__2672\ : InMux
    port map (
            O => \N__24233\,
            I => \N__24226\
        );

    \I__2671\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24223\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24218\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__24226\,
            I => \N__24218\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__24223\,
            I => n2713
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__24218\,
            I => n2713
        );

    \I__2666\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24210\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__24210\,
            I => \N__24206\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__24209\,
            I => \N__24203\
        );

    \I__2663\ : Span4Mux_v
    port map (
            O => \N__24206\,
            I => \N__24200\
        );

    \I__2662\ : InMux
    port map (
            O => \N__24203\,
            I => \N__24197\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__24200\,
            I => n2592
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__24197\,
            I => n2592
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__24192\,
            I => \n14889_cascade_\
        );

    \I__2658\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24185\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__24188\,
            I => \N__24182\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24179\
        );

    \I__2655\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24175\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__24179\,
            I => \N__24171\
        );

    \I__2653\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24168\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__24175\,
            I => \N__24165\
        );

    \I__2651\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24162\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__24171\,
            I => n2525
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__24168\,
            I => n2525
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__24165\,
            I => n2525
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__24162\,
            I => n2525
        );

    \I__2646\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24150\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__24150\,
            I => \N__24147\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__24147\,
            I => n2582
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__24144\,
            I => \N__24140\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__24143\,
            I => \N__24137\
        );

    \I__2641\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24134\
        );

    \I__2640\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24131\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__24134\,
            I => \N__24127\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__24131\,
            I => \N__24124\
        );

    \I__2637\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24121\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__24127\,
            I => n2515
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__24124\,
            I => n2515
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__24121\,
            I => n2515
        );

    \I__2633\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24110\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__24113\,
            I => \N__24107\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__24110\,
            I => \N__24103\
        );

    \I__2630\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24100\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__24106\,
            I => \N__24097\
        );

    \I__2628\ : Span4Mux_v
    port map (
            O => \N__24103\,
            I => \N__24094\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__24100\,
            I => \N__24091\
        );

    \I__2626\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24088\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__24094\,
            I => n2531
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__24091\,
            I => n2531
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__24088\,
            I => n2531
        );

    \I__2622\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24075\
        );

    \I__2620\ : Span4Mux_v
    port map (
            O => \N__24075\,
            I => \N__24072\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__24072\,
            I => n2598
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__24069\,
            I => \N__24066\
        );

    \I__2617\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24063\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24058\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__24062\,
            I => \N__24055\
        );

    \I__2614\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24052\
        );

    \I__2613\ : Span4Mux_v
    port map (
            O => \N__24058\,
            I => \N__24049\
        );

    \I__2612\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24046\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__24052\,
            I => \N__24043\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__24049\,
            I => n2727
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__24046\,
            I => n2727
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__24043\,
            I => n2727
        );

    \I__2607\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24033\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__24033\,
            I => \N__24030\
        );

    \I__2605\ : Span4Mux_h
    port map (
            O => \N__24030\,
            I => \N__24027\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__24027\,
            I => n2585
        );

    \I__2603\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24020\
        );

    \I__2602\ : InMux
    port map (
            O => \N__24023\,
            I => \N__24017\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__24013\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__24017\,
            I => \N__24010\
        );

    \I__2599\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24007\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__24013\,
            I => \N__24004\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__24010\,
            I => n2518
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__24007\,
            I => n2518
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__24004\,
            I => n2518
        );

    \I__2594\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23994\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__23994\,
            I => n14658
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__23991\,
            I => \n2617_cascade_\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__23988\,
            I => \N__23985\
        );

    \I__2590\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23982\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__23982\,
            I => n14324
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__23979\,
            I => \N__23976\
        );

    \I__2587\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23972\
        );

    \I__2586\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23969\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__23972\,
            I => n2516
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__23969\,
            I => n2516
        );

    \I__2583\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23959\
        );

    \I__2582\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23956\
        );

    \I__2581\ : InMux
    port map (
            O => \N__23962\,
            I => \N__23953\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23950\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__23956\,
            I => \N__23945\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__23953\,
            I => \N__23945\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__23950\,
            I => \N__23942\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__23945\,
            I => n2512
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__23942\,
            I => n2512
        );

    \I__2574\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23933\
        );

    \I__2573\ : InMux
    port map (
            O => \N__23936\,
            I => \N__23930\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__23933\,
            I => \N__23924\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23924\
        );

    \I__2570\ : InMux
    port map (
            O => \N__23929\,
            I => \N__23921\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__23924\,
            I => n2513
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__23921\,
            I => n2513
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__23916\,
            I => \n14330_cascade_\
        );

    \I__2566\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23909\
        );

    \I__2565\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23906\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23903\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__23906\,
            I => \N__23900\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__23903\,
            I => \N__23897\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__23900\,
            I => n2511
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__23897\,
            I => n2511
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__23892\,
            I => \N__23889\
        );

    \I__2558\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23884\
        );

    \I__2557\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23879\
        );

    \I__2556\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23879\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__23884\,
            I => n2523
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__23879\,
            I => n2523
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__23874\,
            I => \n2544_cascade_\
        );

    \I__2552\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__23868\,
            I => \N__23865\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__23865\,
            I => n2590
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__23862\,
            I => \N__23859\
        );

    \I__2548\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__23856\,
            I => \N__23853\
        );

    \I__2546\ : Odrv12
    port map (
            O => \N__23853\,
            I => n2591
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__23850\,
            I => \N__23846\
        );

    \I__2544\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23843\
        );

    \I__2543\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23840\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__23843\,
            I => \N__23837\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__23840\,
            I => \N__23834\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__23837\,
            I => \N__23830\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__23834\,
            I => \N__23827\
        );

    \I__2538\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23824\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__23830\,
            I => n2530
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__23827\,
            I => n2530
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__23824\,
            I => n2530
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__23817\,
            I => \N__23814\
        );

    \I__2533\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23811\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__23811\,
            I => \N__23808\
        );

    \I__2531\ : Span4Mux_h
    port map (
            O => \N__23808\,
            I => \N__23805\
        );

    \I__2530\ : Span4Mux_s0_h
    port map (
            O => \N__23805\,
            I => \N__23802\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__23802\,
            I => n2597
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__23799\,
            I => \n2629_cascade_\
        );

    \I__2527\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23793\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__23793\,
            I => n14656
        );

    \I__2525\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23787\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__23784\,
            I => \N__23781\
        );

    \I__2522\ : Sp12to4
    port map (
            O => \N__23781\,
            I => \N__23778\
        );

    \I__2521\ : Odrv12
    port map (
            O => \N__23778\,
            I => n2601
        );

    \I__2520\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23772\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23769\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__23769\,
            I => n2584
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__23766\,
            I => \N__23762\
        );

    \I__2516\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23759\
        );

    \I__2515\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23756\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__23759\,
            I => \N__23752\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__23756\,
            I => \N__23749\
        );

    \I__2512\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23746\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__23752\,
            I => n2517
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__23749\,
            I => n2517
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__23746\,
            I => n2517
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__23739\,
            I => \n2328_cascade_\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__23736\,
            I => \n14442_cascade_\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__23733\,
            I => \n14448_cascade_\
        );

    \I__2505\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__23727\,
            I => n14450
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__23724\,
            I => \N__23721\
        );

    \I__2502\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23718\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__23718\,
            I => \N__23715\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__23715\,
            I => n2593
        );

    \I__2499\ : InMux
    port map (
            O => \N__23712\,
            I => \N__23708\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__23711\,
            I => \N__23705\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__23708\,
            I => \N__23701\
        );

    \I__2496\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23698\
        );

    \I__2495\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23695\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__23701\,
            I => n2422
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__23698\,
            I => n2422
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__23695\,
            I => n2422
        );

    \I__2491\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23685\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__2489\ : Span4Mux_h
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__23679\,
            I => n2489
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__2486\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23669\
        );

    \I__2485\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23666\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__23669\,
            I => \N__23663\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__23666\,
            I => n2521
        );

    \I__2482\ : Odrv12
    port map (
            O => \N__23663\,
            I => n2521
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__2480\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23650\
        );

    \I__2479\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23645\
        );

    \I__2478\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23645\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__23650\,
            I => n2526
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__23645\,
            I => n2526
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__23640\,
            I => \n2521_cascade_\
        );

    \I__2474\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23634\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__23634\,
            I => n14312
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__23631\,
            I => \N__23628\
        );

    \I__2471\ : InMux
    port map (
            O => \N__23628\,
            I => \N__23624\
        );

    \I__2470\ : InMux
    port map (
            O => \N__23627\,
            I => \N__23620\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__23624\,
            I => \N__23617\
        );

    \I__2468\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23614\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__23620\,
            I => n2423
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__23617\,
            I => n2423
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__23614\,
            I => n2423
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__23607\,
            I => \n2425_cascade_\
        );

    \I__2463\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23601\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__23601\,
            I => n14632
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__23598\,
            I => \N__23594\
        );

    \I__2460\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23591\
        );

    \I__2459\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23588\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__23591\,
            I => \N__23585\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__23588\,
            I => \N__23582\
        );

    \I__2456\ : Span4Mux_v
    port map (
            O => \N__23585\,
            I => \N__23578\
        );

    \I__2455\ : Span4Mux_s3_h
    port map (
            O => \N__23582\,
            I => \N__23575\
        );

    \I__2454\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23572\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__23578\,
            I => n2419
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__23575\,
            I => n2419
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__23572\,
            I => n2419
        );

    \I__2450\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23561\
        );

    \I__2449\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23557\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23554\
        );

    \I__2447\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23551\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__23557\,
            I => n2415
        );

    \I__2445\ : Odrv12
    port map (
            O => \N__23554\,
            I => n2415
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__23551\,
            I => n2415
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__23544\,
            I => \n14456_cascade_\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__23541\,
            I => \n2346_cascade_\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__23538\,
            I => \N__23534\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__23537\,
            I => \N__23531\
        );

    \I__2439\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23528\
        );

    \I__2438\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23525\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__23528\,
            I => \N__23521\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__23525\,
            I => \N__23518\
        );

    \I__2435\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23515\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__23521\,
            I => n2417
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__23518\,
            I => n2417
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__23515\,
            I => n2417
        );

    \I__2431\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23503\
        );

    \I__2430\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23500\
        );

    \I__2429\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23497\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__23503\,
            I => \N__23494\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__23500\,
            I => \N__23491\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__23497\,
            I => n2414
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__23494\,
            I => n2414
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__23491\,
            I => n2414
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__23484\,
            I => \N__23481\
        );

    \I__2422\ : InMux
    port map (
            O => \N__23481\,
            I => \N__23478\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__23478\,
            I => \N__23475\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__23475\,
            I => n13790
        );

    \I__2419\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23469\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__23469\,
            I => n14318
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__23466\,
            I => \N__23463\
        );

    \I__2416\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23456\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__23459\,
            I => \N__23453\
        );

    \I__2413\ : Span4Mux_v
    port map (
            O => \N__23456\,
            I => \N__23450\
        );

    \I__2412\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23447\
        );

    \I__2411\ : Span4Mux_s1_h
    port map (
            O => \N__23450\,
            I => \N__23441\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__23447\,
            I => \N__23441\
        );

    \I__2409\ : InMux
    port map (
            O => \N__23446\,
            I => \N__23438\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__23441\,
            I => n2529
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__23438\,
            I => n2529
        );

    \I__2406\ : InMux
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__23430\,
            I => n11942
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__2403\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__23421\,
            I => n13816
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__23418\,
            I => \n14622_cascade_\
        );

    \I__2400\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__23412\,
            I => n14638
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__23409\,
            I => \N__23406\
        );

    \I__2397\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23402\
        );

    \I__2396\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23399\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23396\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__23399\,
            I => n2420
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__23396\,
            I => n2420
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__23391\,
            I => \n2420_cascade_\
        );

    \I__2391\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__23385\,
            I => n14612
        );

    \I__2389\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23379\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__23379\,
            I => n14616
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__23376\,
            I => \N__23373\
        );

    \I__2386\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23369\
        );

    \I__2385\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23365\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__23369\,
            I => \N__23362\
        );

    \I__2383\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23359\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__23365\,
            I => n2426
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__23362\,
            I => n2426
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__23359\,
            I => n2426
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__23352\,
            I => \N__23348\
        );

    \I__2378\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23345\
        );

    \I__2377\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23342\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23338\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23335\
        );

    \I__2374\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23332\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__23338\,
            I => n2421
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__23335\,
            I => n2421
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__23332\,
            I => n2421
        );

    \I__2370\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23321\
        );

    \I__2369\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23318\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23315\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23311\
        );

    \I__2366\ : Span4Mux_s2_h
    port map (
            O => \N__23315\,
            I => \N__23308\
        );

    \I__2365\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23305\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__23311\,
            I => n2413
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__23308\,
            I => n2413
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__23305\,
            I => n2413
        );

    \I__2361\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23294\
        );

    \I__2360\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23291\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__23294\,
            I => \debounce.cnt_reg_9\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__23291\,
            I => \debounce.cnt_reg_9\
        );

    \I__2357\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23282\
        );

    \I__2356\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23279\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__23282\,
            I => \debounce.cnt_reg_8\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__23279\,
            I => \debounce.cnt_reg_8\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__2352\ : InMux
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__23268\,
            I => \N__23264\
        );

    \I__2350\ : InMux
    port map (
            O => \N__23267\,
            I => \N__23261\
        );

    \I__2349\ : Span4Mux_s1_v
    port map (
            O => \N__23264\,
            I => \N__23258\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__23261\,
            I => \debounce.cnt_reg_4\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__23258\,
            I => \debounce.cnt_reg_4\
        );

    \I__2346\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23249\
        );

    \I__2345\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23246\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__23249\,
            I => \debounce.cnt_reg_5\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__23246\,
            I => \debounce.cnt_reg_5\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__23241\,
            I => \N__23238\
        );

    \I__2341\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23235\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__23235\,
            I => n2976
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__23232\,
            I => \N__23228\
        );

    \I__2338\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23225\
        );

    \I__2337\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__23225\,
            I => \N__23217\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__23222\,
            I => \N__23217\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__23217\,
            I => n2432
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__23214\,
            I => \n2432_cascade_\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__23211\,
            I => \N__23208\
        );

    \I__2331\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23204\
        );

    \I__2330\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23201\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__23204\,
            I => n2433
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__23201\,
            I => n2433
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__23196\,
            I => \N__23193\
        );

    \I__2326\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23188\
        );

    \I__2325\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23185\
        );

    \I__2324\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23182\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__23188\,
            I => n2431
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__23185\,
            I => n2431
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__23182\,
            I => n2431
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__23175\,
            I => \N__23171\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__23174\,
            I => \N__23167\
        );

    \I__2318\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23164\
        );

    \I__2317\ : InMux
    port map (
            O => \N__23170\,
            I => \N__23161\
        );

    \I__2316\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23158\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__23164\,
            I => n2430
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__23161\,
            I => n2430
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__23158\,
            I => n2430
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__23151\,
            I => \n11946_cascade_\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__23148\,
            I => \N__23145\
        );

    \I__2310\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23140\
        );

    \I__2309\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23137\
        );

    \I__2308\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23134\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__23140\,
            I => \N__23131\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__23137\,
            I => n2429
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__23134\,
            I => n2429
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__23131\,
            I => n2429
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__23124\,
            I => \N__23120\
        );

    \I__2302\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23117\
        );

    \I__2301\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23114\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23111\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__23114\,
            I => \N__23108\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__23111\,
            I => n2427
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__23108\,
            I => n2427
        );

    \I__2296\ : InMux
    port map (
            O => \N__23103\,
            I => \N__23099\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__23102\,
            I => \N__23096\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__23099\,
            I => \N__23092\
        );

    \I__2293\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23089\
        );

    \I__2292\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23086\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__23092\,
            I => n2424
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__23089\,
            I => n2424
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__23086\,
            I => n2424
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__23079\,
            I => \n2427_cascade_\
        );

    \I__2287\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23072\
        );

    \I__2286\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23069\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__23072\,
            I => \N__23066\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__23069\,
            I => \N__23063\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__23066\,
            I => n2428
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__23063\,
            I => n2428
        );

    \I__2281\ : InMux
    port map (
            O => \N__23058\,
            I => n12842
        );

    \I__2280\ : InMux
    port map (
            O => \N__23055\,
            I => n12843
        );

    \I__2279\ : InMux
    port map (
            O => \N__23052\,
            I => n12844
        );

    \I__2278\ : InMux
    port map (
            O => \N__23049\,
            I => n12845
        );

    \I__2277\ : InMux
    port map (
            O => \N__23046\,
            I => \bfn_2_32_0_\
        );

    \I__2276\ : InMux
    port map (
            O => \N__23043\,
            I => n12847
        );

    \I__2275\ : InMux
    port map (
            O => \N__23040\,
            I => n12848
        );

    \I__2274\ : InMux
    port map (
            O => \N__23037\,
            I => n12849
        );

    \I__2273\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23030\
        );

    \I__2272\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23027\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__23030\,
            I => \debounce.cnt_reg_0\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__23027\,
            I => \debounce.cnt_reg_0\
        );

    \I__2269\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23018\
        );

    \I__2268\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23015\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__23018\,
            I => \debounce.cnt_reg_7\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__23015\,
            I => \debounce.cnt_reg_7\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__23010\,
            I => \N__23006\
        );

    \I__2264\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23003\
        );

    \I__2263\ : InMux
    port map (
            O => \N__23006\,
            I => \N__23000\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__23003\,
            I => \debounce.cnt_reg_1\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__23000\,
            I => \debounce.cnt_reg_1\
        );

    \I__2260\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22991\
        );

    \I__2259\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22988\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__22991\,
            I => \debounce.cnt_reg_2\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__22988\,
            I => \debounce.cnt_reg_2\
        );

    \I__2256\ : InMux
    port map (
            O => \N__22983\,
            I => n12833
        );

    \I__2255\ : InMux
    port map (
            O => \N__22980\,
            I => n12834
        );

    \I__2254\ : InMux
    port map (
            O => \N__22977\,
            I => n12835
        );

    \I__2253\ : InMux
    port map (
            O => \N__22974\,
            I => n12836
        );

    \I__2252\ : InMux
    port map (
            O => \N__22971\,
            I => n12837
        );

    \I__2251\ : InMux
    port map (
            O => \N__22968\,
            I => \bfn_2_31_0_\
        );

    \I__2250\ : InMux
    port map (
            O => \N__22965\,
            I => n12839
        );

    \I__2249\ : InMux
    port map (
            O => \N__22962\,
            I => n12840
        );

    \I__2248\ : InMux
    port map (
            O => \N__22959\,
            I => n12841
        );

    \I__2247\ : InMux
    port map (
            O => \N__22956\,
            I => n12824
        );

    \I__2246\ : InMux
    port map (
            O => \N__22953\,
            I => n12825
        );

    \I__2245\ : InMux
    port map (
            O => \N__22950\,
            I => n12826
        );

    \I__2244\ : InMux
    port map (
            O => \N__22947\,
            I => n12827
        );

    \I__2243\ : InMux
    port map (
            O => \N__22944\,
            I => n12828
        );

    \I__2242\ : InMux
    port map (
            O => \N__22941\,
            I => n12829
        );

    \I__2241\ : InMux
    port map (
            O => \N__22938\,
            I => \bfn_2_30_0_\
        );

    \I__2240\ : InMux
    port map (
            O => \N__22935\,
            I => n12831
        );

    \I__2239\ : InMux
    port map (
            O => \N__22932\,
            I => n12832
        );

    \I__2238\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__22926\,
            I => \N__22923\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__22923\,
            I => n2780
        );

    \I__2235\ : InMux
    port map (
            O => \N__22920\,
            I => \N__22916\
        );

    \I__2234\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22913\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22909\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__22913\,
            I => \N__22906\
        );

    \I__2231\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22903\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__22909\,
            I => n2817
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__22906\,
            I => n2817
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__22903\,
            I => n2817
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__22896\,
            I => \N__22893\
        );

    \I__2226\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22890\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__22890\,
            I => n2884
        );

    \I__2224\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__22884\,
            I => n2877
        );

    \I__2222\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__22875\,
            I => n2897
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__2218\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22861\
        );

    \I__2216\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22858\
        );

    \I__2215\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22855\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__22861\,
            I => n2830
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__22858\,
            I => n2830
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__22855\,
            I => n2830
        );

    \I__2211\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22844\
        );

    \I__2210\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22841\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__22844\,
            I => n2811
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__22841\,
            I => n2811
        );

    \I__2207\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__22833\,
            I => n2878
        );

    \I__2205\ : InMux
    port map (
            O => \N__22830\,
            I => \bfn_2_29_0_\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__22827\,
            I => \N__22824\
        );

    \I__2203\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22820\
        );

    \I__2202\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22817\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__22820\,
            I => n2933
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__22817\,
            I => n2933
        );

    \I__2199\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22809\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__22809\,
            I => n3000
        );

    \I__2197\ : InMux
    port map (
            O => \N__22806\,
            I => n12823
        );

    \I__2196\ : InMux
    port map (
            O => \N__22803\,
            I => \N__22800\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__22800\,
            I => \N__22797\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__22797\,
            I => n2789
        );

    \I__2193\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22789\
        );

    \I__2192\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22784\
        );

    \I__2191\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22784\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__22789\,
            I => \N__22779\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__22784\,
            I => \N__22779\
        );

    \I__2188\ : Odrv12
    port map (
            O => \N__22779\,
            I => n2711
        );

    \I__2187\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22773\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__22773\,
            I => \N__22770\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__22770\,
            I => n2778
        );

    \I__2184\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22764\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__22761\,
            I => n2781
        );

    \I__2181\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22753\
        );

    \I__2180\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22750\
        );

    \I__2179\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22747\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__22753\,
            I => n2714
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__22750\,
            I => n2714
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__22747\,
            I => n2714
        );

    \I__2175\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22737\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__2173\ : Odrv12
    port map (
            O => \N__22734\,
            I => n2800
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__2171\ : InMux
    port map (
            O => \N__22728\,
            I => \N__22724\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__22727\,
            I => \N__22720\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__22724\,
            I => \N__22717\
        );

    \I__2168\ : InMux
    port map (
            O => \N__22723\,
            I => \N__22714\
        );

    \I__2167\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22711\
        );

    \I__2166\ : Span4Mux_s3_v
    port map (
            O => \N__22717\,
            I => \N__22706\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__22714\,
            I => \N__22706\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__22711\,
            I => n2832
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__22706\,
            I => n2832
        );

    \I__2162\ : InMux
    port map (
            O => \N__22701\,
            I => \N__22698\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__2160\ : Odrv12
    port map (
            O => \N__22695\,
            I => n2794
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__22692\,
            I => \N__22689\
        );

    \I__2158\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22686\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__22686\,
            I => n2887
        );

    \I__2156\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22677\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__22677\,
            I => n2779
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__22674\,
            I => \n2811_cascade_\
        );

    \I__2152\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22668\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__22668\,
            I => \N__22665\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__22665\,
            I => n14708
        );

    \I__2149\ : InMux
    port map (
            O => \N__22662\,
            I => n12791
        );

    \I__2148\ : InMux
    port map (
            O => \N__22659\,
            I => n12792
        );

    \I__2147\ : InMux
    port map (
            O => \N__22656\,
            I => n12793
        );

    \I__2146\ : InMux
    port map (
            O => \N__22653\,
            I => n12794
        );

    \I__2145\ : InMux
    port map (
            O => \N__22650\,
            I => \bfn_2_26_0_\
        );

    \I__2144\ : InMux
    port map (
            O => \N__22647\,
            I => n12796
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__22644\,
            I => \n14158_cascade_\
        );

    \I__2142\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__22638\,
            I => \N__22635\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__22635\,
            I => n2790
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__22632\,
            I => \n2742_cascade_\
        );

    \I__2138\ : InMux
    port map (
            O => \N__22629\,
            I => n12783
        );

    \I__2137\ : InMux
    port map (
            O => \N__22626\,
            I => n12784
        );

    \I__2136\ : InMux
    port map (
            O => \N__22623\,
            I => n12785
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__22620\,
            I => \N__22617\
        );

    \I__2134\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22613\
        );

    \I__2133\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22610\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__22613\,
            I => n2719
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__22610\,
            I => n2719
        );

    \I__2130\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22602\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__22602\,
            I => n2786
        );

    \I__2128\ : InMux
    port map (
            O => \N__22599\,
            I => n12786
        );

    \I__2127\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22593\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__22593\,
            I => n2785
        );

    \I__2125\ : InMux
    port map (
            O => \N__22590\,
            I => \bfn_2_25_0_\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__2123\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__22581\,
            I => n2784
        );

    \I__2121\ : InMux
    port map (
            O => \N__22578\,
            I => n12788
        );

    \I__2120\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22572\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__22572\,
            I => n2783
        );

    \I__2118\ : InMux
    port map (
            O => \N__22569\,
            I => n12789
        );

    \I__2117\ : InMux
    port map (
            O => \N__22566\,
            I => \N__22563\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__22563\,
            I => n2782
        );

    \I__2115\ : InMux
    port map (
            O => \N__22560\,
            I => n12790
        );

    \I__2114\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22554\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__22554\,
            I => \N__22551\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__22551\,
            I => n2798
        );

    \I__2111\ : InMux
    port map (
            O => \N__22548\,
            I => n12774
        );

    \I__2110\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__22542\,
            I => \N__22539\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__22539\,
            I => n2797
        );

    \I__2107\ : InMux
    port map (
            O => \N__22536\,
            I => n12775
        );

    \I__2106\ : InMux
    port map (
            O => \N__22533\,
            I => n12776
        );

    \I__2105\ : InMux
    port map (
            O => \N__22530\,
            I => n12777
        );

    \I__2104\ : InMux
    port map (
            O => \N__22527\,
            I => n12778
        );

    \I__2103\ : InMux
    port map (
            O => \N__22524\,
            I => \bfn_2_24_0_\
        );

    \I__2102\ : InMux
    port map (
            O => \N__22521\,
            I => n12780
        );

    \I__2101\ : InMux
    port map (
            O => \N__22518\,
            I => n12781
        );

    \I__2100\ : InMux
    port map (
            O => \N__22515\,
            I => n12782
        );

    \I__2099\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22509\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__22509\,
            I => n2586
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__22506\,
            I => \N__22503\
        );

    \I__2096\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22500\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__22500\,
            I => \N__22496\
        );

    \I__2094\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22493\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__22496\,
            I => \N__22487\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22487\
        );

    \I__2091\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22484\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__22487\,
            I => \N__22481\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22478\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__22481\,
            I => n2519
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__22478\,
            I => n2519
        );

    \I__2086\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__22470\,
            I => \N__22467\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__22467\,
            I => \N__22464\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__22464\,
            I => n2484
        );

    \I__2082\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__22458\,
            I => n2583
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__22455\,
            I => \n2516_cascade_\
        );

    \I__2079\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__22449\,
            I => n2588
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__22446\,
            I => \N__22443\
        );

    \I__2076\ : InMux
    port map (
            O => \N__22443\,
            I => \N__22440\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__22440\,
            I => n2580
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__22437\,
            I => \n2612_cascade_\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__22434\,
            I => \N__22431\
        );

    \I__2072\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__22428\,
            I => \N__22425\
        );

    \I__2070\ : Sp12to4
    port map (
            O => \N__22425\,
            I => \N__22422\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__22422\,
            I => n2801
        );

    \I__2068\ : InMux
    port map (
            O => \N__22419\,
            I => \bfn_2_23_0_\
        );

    \I__2067\ : InMux
    port map (
            O => \N__22416\,
            I => n12772
        );

    \I__2066\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22410\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22407\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__22407\,
            I => n2799
        );

    \I__2063\ : InMux
    port map (
            O => \N__22404\,
            I => n12773
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__22401\,
            I => \n14650_cascade_\
        );

    \I__2061\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22395\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__22395\,
            I => n2595
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__2058\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22385\
        );

    \I__2057\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22382\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__22385\,
            I => \N__22378\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22375\
        );

    \I__2054\ : InMux
    port map (
            O => \N__22381\,
            I => \N__22372\
        );

    \I__2053\ : Odrv12
    port map (
            O => \N__22378\,
            I => n2528
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__22375\,
            I => n2528
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__22372\,
            I => n2528
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__22365\,
            I => \n2627_cascade_\
        );

    \I__2049\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22359\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__22359\,
            I => n14646
        );

    \I__2047\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22352\
        );

    \I__2046\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22349\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22343\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__22349\,
            I => \N__22343\
        );

    \I__2043\ : InMux
    port map (
            O => \N__22348\,
            I => \N__22340\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__22343\,
            I => n2520
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__22340\,
            I => n2520
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__2039\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__22329\,
            I => n2587
        );

    \I__2037\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__22323\,
            I => n2589
        );

    \I__2035\ : InMux
    port map (
            O => \N__22320\,
            I => \N__22316\
        );

    \I__2034\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22313\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22307\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22307\
        );

    \I__2031\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22304\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__22307\,
            I => n2522
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__22304\,
            I => n2522
        );

    \I__2028\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22296\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__22293\,
            I => n2596
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__22290\,
            I => \n2628_cascade_\
        );

    \I__2024\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__22284\,
            I => n14644
        );

    \I__2022\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22277\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__22280\,
            I => \N__22274\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__22277\,
            I => \N__22271\
        );

    \I__2019\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22268\
        );

    \I__2018\ : Odrv12
    port map (
            O => \N__22271\,
            I => n2527
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__22268\,
            I => n2527
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__22263\,
            I => \N__22260\
        );

    \I__2015\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22257\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__22257\,
            I => \N__22254\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__22254\,
            I => n2594
        );

    \I__2012\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22248\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__22248\,
            I => n2579
        );

    \I__2010\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__22239\,
            I => n2491
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__22236\,
            I => \N__22233\
        );

    \I__2006\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22230\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__22230\,
            I => n2481
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__22227\,
            I => \N__22224\
        );

    \I__2003\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22221\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__22221\,
            I => n14310
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__22218\,
            I => \N__22215\
        );

    \I__2000\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22212\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__22209\,
            I => n2494
        );

    \I__1997\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22203\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22200\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__22200\,
            I => n2483
        );

    \I__1994\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22192\
        );

    \I__1993\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22189\
        );

    \I__1992\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22186\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__22192\,
            I => n2416
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__22189\,
            I => n2416
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__22186\,
            I => n2416
        );

    \I__1988\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22176\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__22176\,
            I => n2480
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__22173\,
            I => \N__22170\
        );

    \I__1985\ : InMux
    port map (
            O => \N__22170\,
            I => \N__22167\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__22167\,
            I => n2482
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__22164\,
            I => \n2418_cascade_\
        );

    \I__1982\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22158\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__22158\,
            I => \N__22155\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__22155\,
            I => n2495
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__22152\,
            I => \n2428_cascade_\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__22149\,
            I => \n2527_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22143\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__22143\,
            I => n2488
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__1974\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22134\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__22134\,
            I => n2493
        );

    \I__1972\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22128\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__22128\,
            I => n2490
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__22125\,
            I => \N__22121\
        );

    \I__1969\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22118\
        );

    \I__1968\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22115\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__22118\,
            I => n2418
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__22115\,
            I => n2418
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__1964\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22104\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__22104\,
            I => n2485
        );

    \I__1962\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22098\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__22098\,
            I => n2498
        );

    \I__1960\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22092\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__22092\,
            I => n2487
        );

    \I__1958\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__22086\,
            I => n2497
        );

    \I__1956\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__22080\,
            I => n2499
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__1953\ : InMux
    port map (
            O => \N__22074\,
            I => \N__22071\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__22071\,
            I => n2496
        );

    \I__1951\ : InMux
    port map (
            O => \N__22068\,
            I => \debounce.n13020\
        );

    \I__1950\ : InMux
    port map (
            O => \N__22065\,
            I => \debounce.n13021\
        );

    \I__1949\ : InMux
    port map (
            O => \N__22062\,
            I => \debounce.n13022\
        );

    \I__1948\ : InMux
    port map (
            O => \N__22059\,
            I => \bfn_1_32_0_\
        );

    \I__1947\ : InMux
    port map (
            O => \N__22056\,
            I => \debounce.n13024\
        );

    \I__1946\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22050\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__22050\,
            I => n2501
        );

    \I__1944\ : InMux
    port map (
            O => \N__22047\,
            I => \N__22044\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__22044\,
            I => n2500
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__22041\,
            I => \n2433_cascade_\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__22038\,
            I => \n2532_cascade_\
        );

    \I__1940\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22032\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__22032\,
            I => \N__22029\
        );

    \I__1938\ : Odrv12
    port map (
            O => \N__22029\,
            I => n2900
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__22026\,
            I => \n2833_cascade_\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__22023\,
            I => \n2932_cascade_\
        );

    \I__1935\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22017\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__22017\,
            I => \N__22014\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__22014\,
            I => \N__22011\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__22011\,
            I => n2901
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__22008\,
            I => \n2933_cascade_\
        );

    \I__1930\ : InMux
    port map (
            O => \N__22005\,
            I => \bfn_1_31_0_\
        );

    \I__1929\ : InMux
    port map (
            O => \N__22002\,
            I => \debounce.n13016\
        );

    \I__1928\ : InMux
    port map (
            O => \N__21999\,
            I => \debounce.n13017\
        );

    \I__1927\ : InMux
    port map (
            O => \N__21996\,
            I => \debounce.n13018\
        );

    \I__1926\ : InMux
    port map (
            O => \N__21993\,
            I => \debounce.n13019\
        );

    \I__1925\ : InMux
    port map (
            O => \N__21990\,
            I => n12818
        );

    \I__1924\ : InMux
    port map (
            O => \N__21987\,
            I => n12819
        );

    \I__1923\ : InMux
    port map (
            O => \N__21984\,
            I => \bfn_1_29_0_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__1920\ : Odrv12
    port map (
            O => \N__21975\,
            I => n2876
        );

    \I__1919\ : InMux
    port map (
            O => \N__21972\,
            I => n12821
        );

    \I__1918\ : InMux
    port map (
            O => \N__21969\,
            I => n12822
        );

    \I__1917\ : InMux
    port map (
            O => \N__21966\,
            I => \N__21963\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__1915\ : Span4Mux_s1_h
    port map (
            O => \N__21960\,
            I => \N__21957\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__21957\,
            I => n11956
        );

    \I__1913\ : InMux
    port map (
            O => \N__21954\,
            I => \N__21951\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__21948\,
            I => n2899
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__21945\,
            I => \N__21942\
        );

    \I__1909\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21939\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__21939\,
            I => \N__21936\
        );

    \I__1907\ : Span4Mux_s1_h
    port map (
            O => \N__21936\,
            I => \N__21932\
        );

    \I__1906\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21929\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__21932\,
            I => n2833
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__21929\,
            I => n2833
        );

    \I__1903\ : InMux
    port map (
            O => \N__21924\,
            I => n12809
        );

    \I__1902\ : InMux
    port map (
            O => \N__21921\,
            I => n12810
        );

    \I__1901\ : InMux
    port map (
            O => \N__21918\,
            I => n12811
        );

    \I__1900\ : InMux
    port map (
            O => \N__21915\,
            I => \bfn_1_28_0_\
        );

    \I__1899\ : InMux
    port map (
            O => \N__21912\,
            I => n12813
        );

    \I__1898\ : InMux
    port map (
            O => \N__21909\,
            I => n12814
        );

    \I__1897\ : InMux
    port map (
            O => \N__21906\,
            I => n12815
        );

    \I__1896\ : InMux
    port map (
            O => \N__21903\,
            I => n12816
        );

    \I__1895\ : InMux
    port map (
            O => \N__21900\,
            I => n12817
        );

    \I__1894\ : InMux
    port map (
            O => \N__21897\,
            I => n12800
        );

    \I__1893\ : InMux
    port map (
            O => \N__21894\,
            I => n12801
        );

    \I__1892\ : InMux
    port map (
            O => \N__21891\,
            I => n12802
        );

    \I__1891\ : InMux
    port map (
            O => \N__21888\,
            I => n12803
        );

    \I__1890\ : InMux
    port map (
            O => \N__21885\,
            I => \bfn_1_27_0_\
        );

    \I__1889\ : InMux
    port map (
            O => \N__21882\,
            I => n12805
        );

    \I__1888\ : InMux
    port map (
            O => \N__21879\,
            I => n12806
        );

    \I__1887\ : InMux
    port map (
            O => \N__21876\,
            I => n12807
        );

    \I__1886\ : InMux
    port map (
            O => \N__21873\,
            I => n12808
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__21870\,
            I => \n13845_cascade_\
        );

    \I__1884\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21864\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__21864\,
            I => n14702
        );

    \I__1882\ : InMux
    port map (
            O => \N__21861\,
            I => \bfn_1_26_0_\
        );

    \I__1881\ : InMux
    port map (
            O => \N__21858\,
            I => n12797
        );

    \I__1880\ : InMux
    port map (
            O => \N__21855\,
            I => n12798
        );

    \I__1879\ : InMux
    port map (
            O => \N__21852\,
            I => n12799
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__21849\,
            I => \N__21846\
        );

    \I__1877\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__21843\,
            I => \N__21840\
        );

    \I__1875\ : Odrv12
    port map (
            O => \N__21840\,
            I => n2486
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__21837\,
            I => \n2816_cascade_\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__21834\,
            I => \n2829_cascade_\
        );

    \I__1872\ : InMux
    port map (
            O => \N__21831\,
            I => \bfn_1_22_0_\
        );

    \I__1871\ : InMux
    port map (
            O => \N__21828\,
            I => n12741
        );

    \I__1870\ : InMux
    port map (
            O => \N__21825\,
            I => n12742
        );

    \I__1869\ : InMux
    port map (
            O => \N__21822\,
            I => n12743
        );

    \I__1868\ : InMux
    port map (
            O => \N__21819\,
            I => n12744
        );

    \I__1867\ : InMux
    port map (
            O => \N__21816\,
            I => n12745
        );

    \I__1866\ : InMux
    port map (
            O => \N__21813\,
            I => n12746
        );

    \I__1865\ : InMux
    port map (
            O => \N__21810\,
            I => n12747
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__21807\,
            I => \n2719_cascade_\
        );

    \I__1863\ : InMux
    port map (
            O => \N__21804\,
            I => n12731
        );

    \I__1862\ : InMux
    port map (
            O => \N__21801\,
            I => \bfn_1_21_0_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__21798\,
            I => n12733
        );

    \I__1860\ : InMux
    port map (
            O => \N__21795\,
            I => n12734
        );

    \I__1859\ : InMux
    port map (
            O => \N__21792\,
            I => n12735
        );

    \I__1858\ : InMux
    port map (
            O => \N__21789\,
            I => n12736
        );

    \I__1857\ : InMux
    port map (
            O => \N__21786\,
            I => n12737
        );

    \I__1856\ : InMux
    port map (
            O => \N__21783\,
            I => n12738
        );

    \I__1855\ : InMux
    port map (
            O => \N__21780\,
            I => n12739
        );

    \I__1854\ : InMux
    port map (
            O => \N__21777\,
            I => n12723
        );

    \I__1853\ : InMux
    port map (
            O => \N__21774\,
            I => n12724
        );

    \I__1852\ : InMux
    port map (
            O => \N__21771\,
            I => \bfn_1_20_0_\
        );

    \I__1851\ : InMux
    port map (
            O => \N__21768\,
            I => n12725
        );

    \I__1850\ : InMux
    port map (
            O => \N__21765\,
            I => n12726
        );

    \I__1849\ : InMux
    port map (
            O => \N__21762\,
            I => n12727
        );

    \I__1848\ : InMux
    port map (
            O => \N__21759\,
            I => n12728
        );

    \I__1847\ : InMux
    port map (
            O => \N__21756\,
            I => n12729
        );

    \I__1846\ : InMux
    port map (
            O => \N__21753\,
            I => n12730
        );

    \I__1845\ : InMux
    port map (
            O => \N__21750\,
            I => n12714
        );

    \I__1844\ : InMux
    port map (
            O => \N__21747\,
            I => n12715
        );

    \I__1843\ : InMux
    port map (
            O => \N__21744\,
            I => n12716
        );

    \I__1842\ : InMux
    port map (
            O => \N__21741\,
            I => n12717
        );

    \I__1841\ : InMux
    port map (
            O => \N__21738\,
            I => \bfn_1_19_0_\
        );

    \I__1840\ : InMux
    port map (
            O => \N__21735\,
            I => n12719
        );

    \I__1839\ : InMux
    port map (
            O => \N__21732\,
            I => n12720
        );

    \I__1838\ : InMux
    port map (
            O => \N__21729\,
            I => n12721
        );

    \I__1837\ : InMux
    port map (
            O => \N__21726\,
            I => n12722
        );

    \I__1836\ : InMux
    port map (
            O => \N__21723\,
            I => n12705
        );

    \I__1835\ : InMux
    port map (
            O => \N__21720\,
            I => n12706
        );

    \I__1834\ : InMux
    port map (
            O => \N__21717\,
            I => n12707
        );

    \I__1833\ : InMux
    port map (
            O => \N__21714\,
            I => n12708
        );

    \I__1832\ : InMux
    port map (
            O => \N__21711\,
            I => n12709
        );

    \I__1831\ : InMux
    port map (
            O => \N__21708\,
            I => \bfn_1_18_0_\
        );

    \I__1830\ : InMux
    port map (
            O => \N__21705\,
            I => n12711
        );

    \I__1829\ : InMux
    port map (
            O => \N__21702\,
            I => n12712
        );

    \I__1828\ : InMux
    port map (
            O => \N__21699\,
            I => n12713
        );

    \I__1827\ : InMux
    port map (
            O => \N__21696\,
            I => \bfn_1_17_0_\
        );

    \I__1826\ : InMux
    port map (
            O => \N__21693\,
            I => n12703
        );

    \I__1825\ : InMux
    port map (
            O => \N__21690\,
            I => n12704
        );

    \I__1824\ : IoInMux
    port map (
            O => \N__21687\,
            I => \N__21684\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__21684\,
            I => \N__21681\
        );

    \I__1822\ : IoSpan4Mux
    port map (
            O => \N__21681\,
            I => \N__21678\
        );

    \I__1821\ : IoSpan4Mux
    port map (
            O => \N__21678\,
            I => \N__21675\
        );

    \I__1820\ : IoSpan4Mux
    port map (
            O => \N__21675\,
            I => \N__21672\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__21672\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_7_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_29_0_\
        );

    \IN_MUX_bfv_7_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12914,
            carryinitout => \bfn_7_30_0_\
        );

    \IN_MUX_bfv_7_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12922,
            carryinitout => \bfn_7_31_0_\
        );

    \IN_MUX_bfv_7_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12930,
            carryinitout => \bfn_7_32_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12442,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12450,
            carryinitout => \bfn_15_27_0_\
        );

    \IN_MUX_bfv_15_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12458,
            carryinitout => \bfn_15_28_0_\
        );

    \IN_MUX_bfv_9_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_30_0_\
        );

    \IN_MUX_bfv_9_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12419,
            carryinitout => \bfn_9_31_0_\
        );

    \IN_MUX_bfv_9_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12427,
            carryinitout => \bfn_9_32_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_17_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13006,
            carryinitout => \bfn_17_27_0_\
        );

    \IN_MUX_bfv_17_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13014,
            carryinitout => \bfn_17_28_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n13032\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n13040\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n13048\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_12_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_26_0_\
        );

    \IN_MUX_bfv_12_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12466,
            carryinitout => \bfn_12_27_0_\
        );

    \IN_MUX_bfv_12_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12474,
            carryinitout => \bfn_12_28_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12975,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12983,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12991,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12545,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12534,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12524,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12515,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12507,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_5_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12885,
            carryinitout => \bfn_5_26_0_\
        );

    \IN_MUX_bfv_5_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12893,
            carryinitout => \bfn_5_27_0_\
        );

    \IN_MUX_bfv_5_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12901,
            carryinitout => \bfn_5_28_0_\
        );

    \IN_MUX_bfv_3_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_29_0_\
        );

    \IN_MUX_bfv_3_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12857,
            carryinitout => \bfn_3_30_0_\
        );

    \IN_MUX_bfv_3_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12865,
            carryinitout => \bfn_3_31_0_\
        );

    \IN_MUX_bfv_3_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12873,
            carryinitout => \bfn_3_32_0_\
        );

    \IN_MUX_bfv_2_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_29_0_\
        );

    \IN_MUX_bfv_2_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12830,
            carryinitout => \bfn_2_30_0_\
        );

    \IN_MUX_bfv_2_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12838,
            carryinitout => \bfn_2_31_0_\
        );

    \IN_MUX_bfv_2_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12846,
            carryinitout => \bfn_2_32_0_\
        );

    \IN_MUX_bfv_1_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_26_0_\
        );

    \IN_MUX_bfv_1_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12804,
            carryinitout => \bfn_1_27_0_\
        );

    \IN_MUX_bfv_1_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12812,
            carryinitout => \bfn_1_28_0_\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12820,
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_2_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12779,
            carryinitout => \bfn_2_24_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12787,
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12795,
            carryinitout => \bfn_2_26_0_\
        );

    \IN_MUX_bfv_4_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_21_0_\
        );

    \IN_MUX_bfv_4_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12755,
            carryinitout => \bfn_4_22_0_\
        );

    \IN_MUX_bfv_4_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12763,
            carryinitout => \bfn_4_23_0_\
        );

    \IN_MUX_bfv_4_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12771,
            carryinitout => \bfn_4_24_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12732,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12740,
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12710,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12718,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12689,
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_4_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12697,
            carryinitout => \bfn_4_19_0_\
        );

    \IN_MUX_bfv_5_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_20_0_\
        );

    \IN_MUX_bfv_5_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12669,
            carryinitout => \bfn_5_21_0_\
        );

    \IN_MUX_bfv_5_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12677,
            carryinitout => \bfn_5_22_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12650,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_5_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12658,
            carryinitout => \bfn_5_19_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_7_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12632,
            carryinitout => \bfn_7_18_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12640,
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12615,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12623,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12599,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12607,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12584,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12570,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12557,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_15_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_31_0_\
        );

    \IN_MUX_bfv_1_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_31_0_\
        );

    \IN_MUX_bfv_1_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \debounce.n13023\,
            carryinitout => \bfn_1_32_0_\
        );

    \IN_MUX_bfv_11_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_29_0_\
        );

    \IN_MUX_bfv_11_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13094,
            carryinitout => \bfn_11_30_0_\
        );

    \IN_MUX_bfv_11_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13102,
            carryinitout => \bfn_11_31_0_\
        );

    \IN_MUX_bfv_11_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13110,
            carryinitout => \bfn_11_32_0_\
        );

    \IN_MUX_bfv_7_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_23_0_\
        );

    \IN_MUX_bfv_7_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12945,
            carryinitout => \bfn_7_24_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12953,
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_12_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_13_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n13063\,
            carryinitout => \bfn_13_27_0_\
        );

    \IN_MUX_bfv_13_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n13071\,
            carryinitout => \bfn_13_28_0_\
        );

    \IN_MUX_bfv_13_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n13079\,
            carryinitout => \bfn_13_29_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21687\,
            GLOBALBUFFEROUTPUT => \CLK_N\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_2_lut_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37816\,
            in2 => \_gnd_net_\,
            in3 => \N__21696\,
            lcout => n2501,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => n12703,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_3_lut_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53441\,
            in2 => \N__23211\,
            in3 => \N__21693\,
            lcout => n2500,
            ltout => OPEN,
            carryin => n12703,
            carryout => n12704,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_4_lut_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23232\,
            in3 => \N__21690\,
            lcout => n2499,
            ltout => OPEN,
            carryin => n12704,
            carryout => n12705,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_5_lut_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23191\,
            in2 => \N__53813\,
            in3 => \N__21723\,
            lcout => n2498,
            ltout => OPEN,
            carryin => n12705,
            carryout => n12706,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_6_lut_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23174\,
            in3 => \N__21720\,
            lcout => n2497,
            ltout => OPEN,
            carryin => n12706,
            carryout => n12707,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_7_lut_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23148\,
            in3 => \N__21717\,
            lcout => n2496,
            ltout => OPEN,
            carryin => n12707,
            carryout => n12708,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_8_lut_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23076\,
            in2 => \N__53812\,
            in3 => \N__21714\,
            lcout => n2495,
            ltout => OPEN,
            carryin => n12708,
            carryout => n12709,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_9_lut_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53445\,
            in2 => \N__23124\,
            in3 => \N__21711\,
            lcout => n2494,
            ltout => OPEN,
            carryin => n12709,
            carryout => n12710,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_10_lut_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53433\,
            in2 => \N__23376\,
            in3 => \N__21708\,
            lcout => n2493,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => n12711,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_11_lut_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53437\,
            in2 => \N__25689\,
            in3 => \N__21705\,
            lcout => n2492,
            ltout => OPEN,
            carryin => n12711,
            carryout => n12712,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_12_lut_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53434\,
            in2 => \N__23102\,
            in3 => \N__21702\,
            lcout => n2491,
            ltout => OPEN,
            carryin => n12712,
            carryout => n12713,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_13_lut_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53438\,
            in2 => \N__23631\,
            in3 => \N__21699\,
            lcout => n2490,
            ltout => OPEN,
            carryin => n12713,
            carryout => n12714,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_14_lut_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53435\,
            in2 => \N__23711\,
            in3 => \N__21750\,
            lcout => n2489,
            ltout => OPEN,
            carryin => n12714,
            carryout => n12715,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_15_lut_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53439\,
            in2 => \N__23352\,
            in3 => \N__21747\,
            lcout => n2488,
            ltout => OPEN,
            carryin => n12715,
            carryout => n12716,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_16_lut_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53436\,
            in2 => \N__23409\,
            in3 => \N__21744\,
            lcout => n2487,
            ltout => OPEN,
            carryin => n12716,
            carryout => n12717,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_17_lut_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53440\,
            in2 => \N__23598\,
            in3 => \N__21741\,
            lcout => n2486,
            ltout => OPEN,
            carryin => n12717,
            carryout => n12718,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_18_lut_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53418\,
            in2 => \N__22125\,
            in3 => \N__21738\,
            lcout => n2485,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => n12719,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_19_lut_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53425\,
            in2 => \N__23537\,
            in3 => \N__21735\,
            lcout => n2484,
            ltout => OPEN,
            carryin => n12719,
            carryout => n12720,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_20_lut_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22196\,
            in2 => \N__53810\,
            in3 => \N__21732\,
            lcout => n2483,
            ltout => OPEN,
            carryin => n12720,
            carryout => n12721,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_21_lut_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23565\,
            in2 => \N__53808\,
            in3 => \N__21729\,
            lcout => n2482,
            ltout => OPEN,
            carryin => n12721,
            carryout => n12722,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_22_lut_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23508\,
            in2 => \N__53811\,
            in3 => \N__21726\,
            lcout => n2481,
            ltout => OPEN,
            carryin => n12722,
            carryout => n12723,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_23_lut_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23325\,
            in2 => \N__53809\,
            in3 => \N__21777\,
            lcout => n2480,
            ltout => OPEN,
            carryin => n12723,
            carryout => n12724,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_24_lut_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53432\,
            in1 => \N__33024\,
            in2 => \N__25521\,
            in3 => \N__21774\,
            lcout => n2511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_2_lut_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28671\,
            in2 => \_gnd_net_\,
            in3 => \N__21771\,
            lcout => n2601,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => n12725,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_3_lut_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53412\,
            in2 => \N__28637\,
            in3 => \N__21768\,
            lcout => n2600,
            ltout => OPEN,
            carryin => n12725,
            carryout => n12726,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_4_lut_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28586\,
            in3 => \N__21765\,
            lcout => n2599,
            ltout => OPEN,
            carryin => n12726,
            carryout => n12727,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_5_lut_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53413\,
            in2 => \N__24113\,
            in3 => \N__21762\,
            lcout => n2598,
            ltout => OPEN,
            carryin => n12727,
            carryout => n12728,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_6_lut_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23850\,
            in3 => \N__21759\,
            lcout => n2597,
            ltout => OPEN,
            carryin => n12728,
            carryout => n12729,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_7_lut_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23459\,
            in3 => \N__21756\,
            lcout => n2596,
            ltout => OPEN,
            carryin => n12729,
            carryout => n12730,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_8_lut_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22388\,
            in2 => \N__53807\,
            in3 => \N__21753\,
            lcout => n2595,
            ltout => OPEN,
            carryin => n12730,
            carryout => n12731,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_9_lut_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53417\,
            in2 => \N__22280\,
            in3 => \N__21804\,
            lcout => n2594,
            ltout => OPEN,
            carryin => n12731,
            carryout => n12732,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_10_lut_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54529\,
            in2 => \N__23658\,
            in3 => \N__21801\,
            lcout => n2593,
            ltout => OPEN,
            carryin => \bfn_1_21_0_\,
            carryout => n12733,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_11_lut_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54534\,
            in2 => \N__24188\,
            in3 => \N__21798\,
            lcout => n2592,
            ltout => OPEN,
            carryin => n12733,
            carryout => n12734,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_12_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54530\,
            in2 => \N__25665\,
            in3 => \N__21795\,
            lcout => n2591,
            ltout => OPEN,
            carryin => n12734,
            carryout => n12735,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_13_lut_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54535\,
            in2 => \N__23892\,
            in3 => \N__21792\,
            lcout => n2590,
            ltout => OPEN,
            carryin => n12735,
            carryout => n12736,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_14_lut_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22319\,
            in2 => \N__54545\,
            in3 => \N__21789\,
            lcout => n2589,
            ltout => OPEN,
            carryin => n12736,
            carryout => n12737,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_15_lut_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54539\,
            in2 => \N__23676\,
            in3 => \N__21786\,
            lcout => n2588,
            ltout => OPEN,
            carryin => n12737,
            carryout => n12738,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_16_lut_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22355\,
            in2 => \N__54546\,
            in3 => \N__21783\,
            lcout => n2587,
            ltout => OPEN,
            carryin => n12738,
            carryout => n12739,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_17_lut_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22499\,
            in2 => \N__54544\,
            in3 => \N__21780\,
            lcout => n2586,
            ltout => OPEN,
            carryin => n12739,
            carryout => n12740,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_18_lut_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24016\,
            in2 => \N__54185\,
            in3 => \N__21831\,
            lcout => n2585,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => n12741,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_19_lut_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53925\,
            in2 => \N__23766\,
            in3 => \N__21828\,
            lcout => n2584,
            ltout => OPEN,
            carryin => n12741,
            carryout => n12742,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_20_lut_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52886\,
            in2 => \N__23979\,
            in3 => \N__21825\,
            lcout => n2583,
            ltout => OPEN,
            carryin => n12742,
            carryout => n12743,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_21_lut_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53926\,
            in2 => \N__24143\,
            in3 => \N__21822\,
            lcout => n2582,
            ltout => OPEN,
            carryin => n12743,
            carryout => n12744,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_22_lut_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24287\,
            in2 => \N__54186\,
            in3 => \N__21819\,
            lcout => n2581,
            ltout => OPEN,
            carryin => n12744,
            carryout => n12745,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_23_lut_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23936\,
            in2 => \N__53195\,
            in3 => \N__21816\,
            lcout => n2580,
            ltout => OPEN,
            carryin => n12745,
            carryout => n12746,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_24_lut_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23962\,
            in2 => \N__54187\,
            in3 => \N__21813\,
            lcout => n2579,
            ltout => OPEN,
            carryin => n12746,
            carryout => n12747,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_25_lut_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__52890\,
            in1 => \N__23912\,
            in2 => \N__33188\,
            in3 => \N__21810\,
            lcout => n2610,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1783_3_lut_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26219\,
            in2 => \N__26199\,
            in3 => \N__33349\,
            lcout => n2719,
            ltout => \n2719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_145_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24061\,
            in2 => \N__21807\,
            in3 => \N__24649\,
            lcout => n14138,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13096_1_lut_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33170\,
            lcout => n15821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1646_3_lut_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23597\,
            in2 => \N__21849\,
            in3 => \N__33000\,
            lcout => n2518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i0_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47662\,
            in1 => \N__34854\,
            in2 => \_gnd_net_\,
            in3 => \N__39543\,
            lcout => h3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55773\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1908_3_lut_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24897\,
            in1 => \N__21981\,
            in2 => \_gnd_net_\,
            in3 => \N__33713\,
            lcout => n2908,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1848_3_lut_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24498\,
            in2 => \N__22587\,
            in3 => \N__33517\,
            lcout => n2816,
            ltout => \n2816_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_40_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26998\,
            in1 => \N__24985\,
            in2 => \N__21837\,
            in3 => \N__21867\,
            lcout => n14708,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1850_3_lut_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22605\,
            in2 => \N__22620\,
            in3 => \N__33516\,
            lcout => n2818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1861_3_lut_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26474\,
            in2 => \N__33522\,
            in3 => \N__22545\,
            lcout => n2829,
            ltout => \n2829_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_38_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__24730\,
            in1 => \N__22864\,
            in2 => \N__21834\,
            in3 => \N__21966\,
            lcout => OPEN,
            ltout => \n13845_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_39_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27037\,
            in1 => \N__22912\,
            in2 => \N__21870\,
            in3 => \N__26577\,
            lcout => n14702,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1862_3_lut_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22557\,
            in2 => \N__26514\,
            in3 => \N__33492\,
            lcout => n2830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1846_3_lut_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24405\,
            in1 => \_gnd_net_\,
            in2 => \N__33523\,
            in3 => \N__22566\,
            lcout => n2814,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1847_3_lut_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22575\,
            in1 => \N__24435\,
            in2 => \_gnd_net_\,
            in3 => \N__33502\,
            lcout => n2815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1849_3_lut_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24477\,
            in1 => \_gnd_net_\,
            in2 => \N__33521\,
            in3 => \N__22596\,
            lcout => n2817,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1863_3_lut_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22413\,
            in2 => \N__26901\,
            in3 => \N__33491\,
            lcout => n2831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_2_lut_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38956\,
            in2 => \_gnd_net_\,
            in3 => \N__21861\,
            lcout => n2901,
            ltout => OPEN,
            carryin => \bfn_1_26_0_\,
            carryout => n12797,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_3_lut_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53028\,
            in2 => \N__21945\,
            in3 => \N__21858\,
            lcout => n2900,
            ltout => OPEN,
            carryin => n12797,
            carryout => n12798,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_4_lut_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22727\,
            in3 => \N__21855\,
            lcout => n2899,
            ltout => OPEN,
            carryin => n12798,
            carryout => n12799,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_5_lut_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53029\,
            in2 => \N__24737\,
            in3 => \N__21852\,
            lcout => n2898,
            ltout => OPEN,
            carryin => n12799,
            carryout => n12800,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_6_lut_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22865\,
            in2 => \_gnd_net_\,
            in3 => \N__21897\,
            lcout => n2897,
            ltout => OPEN,
            carryin => n12800,
            carryout => n12801,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_7_lut_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24680\,
            in3 => \N__21894\,
            lcout => n2896,
            ltout => OPEN,
            carryin => n12801,
            carryout => n12802,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_8_lut_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53031\,
            in2 => \N__27099\,
            in3 => \N__21891\,
            lcout => n2895,
            ltout => OPEN,
            carryin => n12802,
            carryout => n12803,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_9_lut_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53030\,
            in2 => \N__26787\,
            in3 => \N__21888\,
            lcout => n2894,
            ltout => OPEN,
            carryin => n12803,
            carryout => n12804,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_10_lut_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54415\,
            in2 => \N__25031\,
            in3 => \N__21885\,
            lcout => n2893,
            ltout => OPEN,
            carryin => \bfn_1_27_0_\,
            carryout => n12805,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_11_lut_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54422\,
            in2 => \N__27885\,
            in3 => \N__21882\,
            lcout => n2892,
            ltout => OPEN,
            carryin => n12805,
            carryout => n12806,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_12_lut_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54416\,
            in2 => \N__30710\,
            in3 => \N__21879\,
            lcout => n2891,
            ltout => OPEN,
            carryin => n12806,
            carryout => n12807,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_13_lut_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54423\,
            in2 => \N__24822\,
            in3 => \N__21876\,
            lcout => n2890,
            ltout => OPEN,
            carryin => n12807,
            carryout => n12808,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_14_lut_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54417\,
            in2 => \N__24540\,
            in3 => \N__21873\,
            lcout => n2889,
            ltout => OPEN,
            carryin => n12808,
            carryout => n12809,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_15_lut_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54424\,
            in2 => \N__24519\,
            in3 => \N__21924\,
            lcout => n2888,
            ltout => OPEN,
            carryin => n12809,
            carryout => n12810,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_16_lut_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54418\,
            in2 => \N__26616\,
            in3 => \N__21921\,
            lcout => n2887,
            ltout => OPEN,
            carryin => n12810,
            carryout => n12811,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_17_lut_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26826\,
            in2 => \N__54507\,
            in3 => \N__21918\,
            lcout => n2886,
            ltout => OPEN,
            carryin => n12811,
            carryout => n12812,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_18_lut_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27044\,
            in2 => \N__54508\,
            in3 => \N__21915\,
            lcout => n2885,
            ltout => OPEN,
            carryin => \bfn_1_28_0_\,
            carryout => n12813,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_19_lut_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22919\,
            in2 => \N__54512\,
            in3 => \N__21912\,
            lcout => n2884,
            ltout => OPEN,
            carryin => n12813,
            carryout => n12814,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_20_lut_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26282\,
            in2 => \N__54509\,
            in3 => \N__21909\,
            lcout => n2883,
            ltout => OPEN,
            carryin => n12814,
            carryout => n12815,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_21_lut_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24992\,
            in2 => \N__54513\,
            in3 => \N__21906\,
            lcout => n2882,
            ltout => OPEN,
            carryin => n12815,
            carryout => n12816,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_22_lut_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27005\,
            in2 => \N__54510\,
            in3 => \N__21903\,
            lcout => n2881,
            ltout => OPEN,
            carryin => n12816,
            carryout => n12817,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_23_lut_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24971\,
            in2 => \N__54514\,
            in3 => \N__21900\,
            lcout => n2880,
            ltout => OPEN,
            carryin => n12817,
            carryout => n12818,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_24_lut_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24704\,
            in2 => \N__54511\,
            in3 => \N__21990\,
            lcout => n2879,
            ltout => OPEN,
            carryin => n12818,
            carryout => n12819,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_25_lut_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22847\,
            in2 => \N__54515\,
            in3 => \N__21987\,
            lcout => n2878,
            ltout => OPEN,
            carryin => n12819,
            carryout => n12820,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_26_lut_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24872\,
            in2 => \N__54516\,
            in3 => \N__21984\,
            lcout => n2877,
            ltout => OPEN,
            carryin => \bfn_1_29_0_\,
            carryout => n12821,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_27_lut_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24896\,
            in2 => \N__54517\,
            in3 => \N__21972\,
            lcout => n2876,
            ltout => OPEN,
            carryin => n12821,
            carryout => n12822,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_28_lut_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__24849\,
            in1 => \N__54455\,
            in2 => \N__33731\,
            in3 => \N__21969\,
            lcout => n2907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9988_3_lut_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38957\,
            in1 => \N__22723\,
            in2 => \_gnd_net_\,
            in3 => \N__21935\,
            lcout => n11956,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i1_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34823\,
            lcout => \reg_B_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1931_3_lut_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21954\,
            in2 => \N__22731\,
            in3 => \N__33707\,
            lcout => n2931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1865_3_lut_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44866\,
            in2 => \N__22434\,
            in3 => \N__33524\,
            lcout => n2833,
            ltout => \n2833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1932_3_lut_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22035\,
            in2 => \N__22026\,
            in3 => \N__33708\,
            lcout => n2932,
            ltout => \n2932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10070_4_lut_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__32432\,
            in1 => \N__27445\,
            in2 => \N__22023\,
            in3 => \N__22823\,
            lcout => n12038,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1933_3_lut_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22020\,
            in1 => \_gnd_net_\,
            in2 => \N__38961\,
            in3 => \N__33706\,
            lcout => n2933,
            ltout => \n2933_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2000_3_lut_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22812\,
            in2 => \N__22008\,
            in3 => \N__33886\,
            lcout => n3032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.cnt_reg_662__i0_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23034\,
            in2 => \_gnd_net_\,
            in3 => \N__22005\,
            lcout => \debounce.cnt_reg_0\,
            ltout => OPEN,
            carryin => \bfn_1_31_0_\,
            carryout => \debounce.n13016\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i1_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23009\,
            in2 => \_gnd_net_\,
            in3 => \N__22002\,
            lcout => \debounce.cnt_reg_1\,
            ltout => OPEN,
            carryin => \debounce.n13016\,
            carryout => \debounce.n13017\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i2_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22995\,
            in2 => \_gnd_net_\,
            in3 => \N__21999\,
            lcout => \debounce.cnt_reg_2\,
            ltout => OPEN,
            carryin => \debounce.n13017\,
            carryout => \debounce.n13018\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i3_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25154\,
            in2 => \_gnd_net_\,
            in3 => \N__21996\,
            lcout => \debounce.cnt_reg_3\,
            ltout => OPEN,
            carryin => \debounce.n13018\,
            carryout => \debounce.n13019\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i4_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23267\,
            in2 => \_gnd_net_\,
            in3 => \N__21993\,
            lcout => \debounce.cnt_reg_4\,
            ltout => OPEN,
            carryin => \debounce.n13019\,
            carryout => \debounce.n13020\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i5_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23253\,
            in2 => \_gnd_net_\,
            in3 => \N__22068\,
            lcout => \debounce.cnt_reg_5\,
            ltout => OPEN,
            carryin => \debounce.n13020\,
            carryout => \debounce.n13021\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i6_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25181\,
            in2 => \_gnd_net_\,
            in3 => \N__22065\,
            lcout => \debounce.cnt_reg_6\,
            ltout => OPEN,
            carryin => \debounce.n13021\,
            carryout => \debounce.n13022\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i7_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23022\,
            in2 => \_gnd_net_\,
            in3 => \N__22062\,
            lcout => \debounce.cnt_reg_7\,
            ltout => OPEN,
            carryin => \debounce.n13022\,
            carryout => \debounce.n13023\,
            clk => \N__55781\,
            ce => 'H',
            sr => \N__27978\
        );

    \debounce.cnt_reg_662__i8_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23286\,
            in2 => \_gnd_net_\,
            in3 => \N__22059\,
            lcout => \debounce.cnt_reg_8\,
            ltout => OPEN,
            carryin => \bfn_1_32_0_\,
            carryout => \debounce.n13024\,
            clk => \N__55785\,
            ce => 'H',
            sr => \N__27974\
        );

    \debounce.cnt_reg_662__i9_LC_1_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23298\,
            in2 => \_gnd_net_\,
            in3 => \N__22056\,
            lcout => \debounce.cnt_reg_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55785\,
            ce => 'H',
            sr => \N__27974\
        );

    \encoder0_position_31__I_0_i1661_3_lut_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37818\,
            in1 => \N__22053\,
            in2 => \_gnd_net_\,
            in3 => \N__32904\,
            lcout => n2533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1593_3_lut_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30579\,
            in1 => \N__25134\,
            in2 => \_gnd_net_\,
            in3 => \N__32818\,
            lcout => n2433,
            ltout => \n2433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1660_3_lut_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22047\,
            in2 => \N__22041\,
            in3 => \N__32905\,
            lcout => n2532,
            ltout => \n2532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9974_3_lut_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28670\,
            in2 => \N__22038\,
            in3 => \N__28618\,
            lcout => n11942,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1658_3_lut_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22101\,
            in2 => \N__23196\,
            in3 => \N__32907\,
            lcout => n2530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1647_3_lut_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23405\,
            in1 => \_gnd_net_\,
            in2 => \N__32952\,
            in3 => \N__22095\,
            lcout => n2519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1657_3_lut_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22089\,
            in2 => \N__23175\,
            in3 => \N__32906\,
            lcout => n2529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1659_3_lut_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22083\,
            in2 => \N__32953\,
            in3 => \N__23231\,
            lcout => n2531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1591_3_lut_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30098\,
            in2 => \N__32820\,
            in3 => \N__25347\,
            lcout => n2431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1584_3_lut_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28143\,
            in2 => \N__25215\,
            in3 => \N__32782\,
            lcout => n2424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1590_3_lut_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28713\,
            in2 => \N__32821\,
            in3 => \N__25332\,
            lcout => n2430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1656_3_lut_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23144\,
            in2 => \N__22077\,
            in3 => \N__32946\,
            lcout => n2528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1582_3_lut_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29703\,
            in2 => \N__32819\,
            in3 => \N__25425\,
            lcout => n2422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1578_3_lut_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25386\,
            in2 => \N__25599\,
            in3 => \N__32792\,
            lcout => n2418,
            ltout => \n2418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_121_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23560\,
            in1 => \N__22195\,
            in2 => \N__22164\,
            in3 => \N__23604\,
            lcout => n14638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1588_3_lut_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25278\,
            in2 => \N__25304\,
            in3 => \N__32768\,
            lcout => n2428,
            ltout => \n2428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1655_3_lut_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22161\,
            in1 => \_gnd_net_\,
            in2 => \N__22152\,
            in3 => \N__32941\,
            lcout => n2527,
            ltout => \n2527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_127_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24174\,
            in1 => \N__22312\,
            in2 => \N__22149\,
            in3 => \N__22381\,
            lcout => n14310,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1576_3_lut_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30247\,
            in1 => \_gnd_net_\,
            in2 => \N__32812\,
            in3 => \N__25365\,
            lcout => n2416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1648_3_lut_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22146\,
            in1 => \_gnd_net_\,
            in2 => \N__32977\,
            in3 => \N__23351\,
            lcout => n2520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1653_3_lut_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23372\,
            in2 => \N__22140\,
            in3 => \N__32940\,
            lcout => n2525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1650_3_lut_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23627\,
            in2 => \N__32976\,
            in3 => \N__22131\,
            lcout => n2522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1645_3_lut_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22124\,
            in2 => \N__22110\,
            in3 => \N__32945\,
            lcout => n2517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1651_3_lut_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23103\,
            in2 => \N__32984\,
            in3 => \N__22245\,
            lcout => n2523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1641_3_lut_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__23506\,
            in1 => \_gnd_net_\,
            in2 => \N__22236\,
            in3 => \N__32965\,
            lcout => n2513,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_128_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22348\,
            in1 => \N__22492\,
            in2 => \N__22227\,
            in3 => \N__23637\,
            lcout => n14318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1654_3_lut_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23123\,
            in2 => \N__22218\,
            in3 => \N__32954\,
            lcout => n2526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1643_3_lut_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22206\,
            in2 => \N__32986\,
            in3 => \N__22197\,
            lcout => n2515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1720_3_lut_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24178\,
            in2 => \N__24209\,
            in3 => \N__33095\,
            lcout => n2624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1640_3_lut_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22179\,
            in2 => \N__32985\,
            in3 => \N__23324\,
            lcout => n2512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1642_3_lut_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23564\,
            in2 => \N__22173\,
            in3 => \N__32958\,
            lcout => n2514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_138_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25762\,
            in1 => \N__25729\,
            in2 => \N__26242\,
            in3 => \N__22287\,
            lcout => OPEN,
            ltout => \n14650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_139_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26215\,
            in1 => \N__26173\,
            in2 => \N__22401\,
            in3 => \N__22362\,
            lcout => n14656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1723_3_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22398\,
            in2 => \N__22392\,
            in3 => \N__33135\,
            lcout => n2627,
            ltout => \n2627_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_137_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25858\,
            in2 => \N__22365\,
            in3 => \N__25828\,
            lcout => n14646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1715_3_lut_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22356\,
            in2 => \N__22335\,
            in3 => \N__33136\,
            lcout => n2619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1717_3_lut_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22326\,
            in1 => \_gnd_net_\,
            in2 => \N__33159\,
            in3 => \N__22320\,
            lcout => n2621,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1724_3_lut_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22299\,
            in2 => \N__23466\,
            in3 => \N__33131\,
            lcout => n2628,
            ltout => \n2628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_135_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22290\,
            in3 => \N__25796\,
            lcout => n14644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1722_3_lut_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22281\,
            in2 => \N__22263\,
            in3 => \N__33121\,
            lcout => n2626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1707_3_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22251\,
            in1 => \_gnd_net_\,
            in2 => \N__33158\,
            in3 => \N__23963\,
            lcout => n2611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1714_3_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22512\,
            in2 => \N__22506\,
            in3 => \N__33125\,
            lcout => n2618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1644_3_lut_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22473\,
            in2 => \N__23538\,
            in3 => \N__32997\,
            lcout => n2516,
            ltout => \n2516_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1711_3_lut_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22461\,
            in1 => \_gnd_net_\,
            in2 => \N__22455\,
            in3 => \N__33126\,
            lcout => n2615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1716_3_lut_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23672\,
            in2 => \N__33157\,
            in3 => \N__22452\,
            lcout => n2620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1708_3_lut_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23937\,
            in2 => \N__22446\,
            in3 => \N__33127\,
            lcout => n2612,
            ltout => \n2612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1775_3_lut_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26391\,
            in2 => \N__22437\,
            in3 => \N__33344\,
            lcout => n2711,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_2_lut_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44870\,
            in2 => \_gnd_net_\,
            in3 => \N__22419\,
            lcout => n2801,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => n12772,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_3_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53708\,
            in2 => \N__26928\,
            in3 => \N__22416\,
            lcout => n2800,
            ltout => OPEN,
            carryin => n12772,
            carryout => n12773,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_4_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26893\,
            in3 => \N__22404\,
            lcout => n2799,
            ltout => OPEN,
            carryin => n12773,
            carryout => n12774,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_5_lut_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53709\,
            in2 => \N__26513\,
            in3 => \N__22548\,
            lcout => n2798,
            ltout => OPEN,
            carryin => n12774,
            carryout => n12775,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_6_lut_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26478\,
            in3 => \N__22536\,
            lcout => n2797,
            ltout => OPEN,
            carryin => n12775,
            carryout => n12776,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_7_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26862\,
            in3 => \N__22533\,
            lcout => n2796,
            ltout => OPEN,
            carryin => n12776,
            carryout => n12777,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_8_lut_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24329\,
            in2 => \N__54009\,
            in3 => \N__22530\,
            lcout => n2795,
            ltout => OPEN,
            carryin => n12777,
            carryout => n12778,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_9_lut_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53713\,
            in2 => \N__24062\,
            in3 => \N__22527\,
            lcout => n2794,
            ltout => OPEN,
            carryin => n12778,
            carryout => n12779,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_10_lut_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53783\,
            in2 => \N__26718\,
            in3 => \N__22524\,
            lcout => n2793,
            ltout => OPEN,
            carryin => \bfn_2_24_0_\,
            carryout => n12780,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_11_lut_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53792\,
            in2 => \N__24650\,
            in3 => \N__22521\,
            lcout => n2792,
            ltout => OPEN,
            carryin => n12780,
            carryout => n12781,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_12_lut_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53784\,
            in2 => \N__26696\,
            in3 => \N__22518\,
            lcout => n2791,
            ltout => OPEN,
            carryin => n12781,
            carryout => n12782,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_13_lut_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53793\,
            in2 => \N__26669\,
            in3 => \N__22515\,
            lcout => n2790,
            ltout => OPEN,
            carryin => n12782,
            carryout => n12783,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_14_lut_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53785\,
            in2 => \N__24374\,
            in3 => \N__22629\,
            lcout => n2789,
            ltout => OPEN,
            carryin => n12783,
            carryout => n12784,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_15_lut_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24611\,
            in2 => \N__54079\,
            in3 => \N__22626\,
            lcout => n2788,
            ltout => OPEN,
            carryin => n12784,
            carryout => n12785,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_16_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26735\,
            in2 => \N__54081\,
            in3 => \N__22623\,
            lcout => n2787,
            ltout => OPEN,
            carryin => n12785,
            carryout => n12786,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_17_lut_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22616\,
            in2 => \N__54080\,
            in3 => \N__22599\,
            lcout => n2786,
            ltout => OPEN,
            carryin => n12786,
            carryout => n12787,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_18_lut_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53616\,
            in2 => \N__24476\,
            in3 => \N__22590\,
            lcout => n2785,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => n12788,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_19_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24494\,
            in2 => \N__53981\,
            in3 => \N__22578\,
            lcout => n2784,
            ltout => OPEN,
            carryin => n12788,
            carryout => n12789,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_20_lut_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53620\,
            in2 => \N__24434\,
            in3 => \N__22569\,
            lcout => n2783,
            ltout => OPEN,
            carryin => n12789,
            carryout => n12790,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_21_lut_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24401\,
            in2 => \N__53982\,
            in3 => \N__22560\,
            lcout => n2782,
            ltout => OPEN,
            carryin => n12790,
            carryout => n12791,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_22_lut_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22757\,
            in2 => \N__53985\,
            in3 => \N__22662\,
            lcout => n2781,
            ltout => OPEN,
            carryin => n12791,
            carryout => n12792,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_23_lut_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24232\,
            in2 => \N__53983\,
            in3 => \N__22659\,
            lcout => n2780,
            ltout => OPEN,
            carryin => n12792,
            carryout => n12793,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_24_lut_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24310\,
            in2 => \N__53986\,
            in3 => \N__22656\,
            lcout => n2779,
            ltout => OPEN,
            carryin => n12793,
            carryout => n12794,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_25_lut_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22794\,
            in2 => \N__53984\,
            in3 => \N__22653\,
            lcout => n2778,
            ltout => OPEN,
            carryin => n12794,
            carryout => n12795,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_26_lut_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24911\,
            in2 => \N__53411\,
            in3 => \N__22650\,
            lcout => n2777,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => n12796,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_27_lut_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54297\,
            in1 => \N__26298\,
            in2 => \N__33551\,
            in3 => \N__22647\,
            lcout => n2808,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22756\,
            in1 => \N__24233\,
            in2 => \N__24312\,
            in3 => \N__24381\,
            lcout => OPEN,
            ltout => \n14158_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12589_4_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24910\,
            in1 => \N__22792\,
            in2 => \N__22644\,
            in3 => \N__26297\,
            lcout => n2742,
            ltout => \n2742_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12449_3_lut_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22641\,
            in2 => \N__22632\,
            in3 => \N__26670\,
            lcout => n2822,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1853_3_lut_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22803\,
            in2 => \N__24375\,
            in3 => \N__33456\,
            lcout => n2821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1842_3_lut_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22793\,
            in1 => \_gnd_net_\,
            in2 => \N__33506\,
            in3 => \N__22776\,
            lcout => n2810,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1778_3_lut_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26013\,
            in1 => \_gnd_net_\,
            in2 => \N__33351\,
            in3 => \N__26043\,
            lcout => n2714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1845_3_lut_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22767\,
            in1 => \N__22758\,
            in2 => \_gnd_net_\,
            in3 => \N__33452\,
            lcout => n2813,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1864_3_lut_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26927\,
            in2 => \N__33503\,
            in3 => \N__22740\,
            lcout => n2832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1858_3_lut_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22701\,
            in2 => \N__24069\,
            in3 => \N__33445\,
            lcout => n2826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1919_3_lut_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26609\,
            in2 => \N__22692\,
            in3 => \N__33647\,
            lcout => n2919,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1843_3_lut_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22683\,
            in2 => \N__33505\,
            in3 => \N__24311\,
            lcout => n2811,
            ltout => \n2811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_41_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24703\,
            in1 => \N__24970\,
            in2 => \N__22674\,
            in3 => \N__22671\,
            lcout => n14714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1844_3_lut_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24234\,
            in2 => \N__33504\,
            in3 => \N__22929\,
            lcout => n2812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1916_3_lut_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22920\,
            in2 => \N__22896\,
            in3 => \N__33667\,
            lcout => n2916,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1909_3_lut_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22887\,
            in2 => \N__33701\,
            in3 => \N__24873\,
            lcout => n2909,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1929_3_lut_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22881\,
            in2 => \N__22872\,
            in3 => \N__33668\,
            lcout => n2929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2054_3_lut_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__27575\,
            in1 => \_gnd_net_\,
            in2 => \N__25110\,
            in3 => \N__37219\,
            lcout => n3118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12621_1_lut_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33669\,
            lcout => n15346,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1910_3_lut_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22848\,
            in2 => \N__33700\,
            in3 => \N__22836\,
            lcout => n2910,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_2_lut_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32433\,
            in2 => \_gnd_net_\,
            in3 => \N__22830\,
            lcout => n3001,
            ltout => OPEN,
            carryin => \bfn_2_29_0_\,
            carryout => n12823,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_3_lut_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53763\,
            in2 => \N__22827\,
            in3 => \N__22806\,
            lcout => n3000,
            ltout => OPEN,
            carryin => n12823,
            carryout => n12824,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_4_lut_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29417\,
            in3 => \N__22956\,
            lcout => n2999,
            ltout => OPEN,
            carryin => n12824,
            carryout => n12825,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_5_lut_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53764\,
            in2 => \N__27452\,
            in3 => \N__22953\,
            lcout => n2998,
            ltout => OPEN,
            carryin => n12825,
            carryout => n12826,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_6_lut_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27167\,
            in3 => \N__22950\,
            lcout => n2997,
            ltout => OPEN,
            carryin => n12826,
            carryout => n12827,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_7_lut_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27285\,
            in3 => \N__22947\,
            lcout => n2996,
            ltout => OPEN,
            carryin => n12827,
            carryout => n12828,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_8_lut_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54062\,
            in2 => \N__27198\,
            in3 => \N__22944\,
            lcout => n2995,
            ltout => OPEN,
            carryin => n12828,
            carryout => n12829,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_9_lut_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53765\,
            in2 => \N__27378\,
            in3 => \N__22941\,
            lcout => n2994,
            ltout => OPEN,
            carryin => n12829,
            carryout => n12830,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_10_lut_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54010\,
            in2 => \N__28917\,
            in3 => \N__22938\,
            lcout => n2993,
            ltout => OPEN,
            carryin => \bfn_2_30_0_\,
            carryout => n12831,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_11_lut_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54354\,
            in2 => \N__28986\,
            in3 => \N__22935\,
            lcout => n2992,
            ltout => OPEN,
            carryin => n12831,
            carryout => n12832,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_12_lut_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54011\,
            in2 => \N__27837\,
            in3 => \N__22932\,
            lcout => n2991,
            ltout => OPEN,
            carryin => n12832,
            carryout => n12833,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_13_lut_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30671\,
            in2 => \N__54262\,
            in3 => \N__22983\,
            lcout => n2990,
            ltout => OPEN,
            carryin => n12833,
            carryout => n12834,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_14_lut_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27551\,
            in2 => \N__54458\,
            in3 => \N__22980\,
            lcout => n2989,
            ltout => OPEN,
            carryin => n12834,
            carryout => n12835,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_15_lut_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27249\,
            in2 => \N__54263\,
            in3 => \N__22977\,
            lcout => n2988,
            ltout => OPEN,
            carryin => n12835,
            carryout => n12836,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_16_lut_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54018\,
            in2 => \N__24792\,
            in3 => \N__22974\,
            lcout => n2987,
            ltout => OPEN,
            carryin => n12836,
            carryout => n12837,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_17_lut_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54358\,
            in2 => \N__27686\,
            in3 => \N__22971\,
            lcout => n2986,
            ltout => OPEN,
            carryin => n12837,
            carryout => n12838,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_18_lut_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27933\,
            in2 => \N__54272\,
            in3 => \N__22968\,
            lcout => n2985,
            ltout => OPEN,
            carryin => \bfn_2_31_0_\,
            carryout => n12839,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_19_lut_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27482\,
            in2 => \N__54278\,
            in3 => \N__22965\,
            lcout => n2984,
            ltout => OPEN,
            carryin => n12839,
            carryout => n12840,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_20_lut_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29356\,
            in2 => \N__54273\,
            in3 => \N__22962\,
            lcout => n2983,
            ltout => OPEN,
            carryin => n12840,
            carryout => n12841,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_21_lut_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27762\,
            in2 => \N__54279\,
            in3 => \N__22959\,
            lcout => n2982,
            ltout => OPEN,
            carryin => n12841,
            carryout => n12842,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_22_lut_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27617\,
            in2 => \N__54274\,
            in3 => \N__23058\,
            lcout => n2981,
            ltout => OPEN,
            carryin => n12842,
            carryout => n12843,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_23_lut_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54052\,
            in2 => \N__27804\,
            in3 => \N__23055\,
            lcout => n2980,
            ltout => OPEN,
            carryin => n12843,
            carryout => n12844,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_24_lut_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27716\,
            in2 => \N__54275\,
            in3 => \N__23052\,
            lcout => n2979,
            ltout => OPEN,
            carryin => n12844,
            carryout => n12845,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_25_lut_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27911\,
            in2 => \N__54280\,
            in3 => \N__23049\,
            lcout => n2978,
            ltout => OPEN,
            carryin => n12845,
            carryout => n12846,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_26_lut_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28031\,
            in2 => \N__54283\,
            in3 => \N__23046\,
            lcout => n2977,
            ltout => OPEN,
            carryin => \bfn_2_32_0_\,
            carryout => n12847,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_27_lut_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27335\,
            in2 => \N__54285\,
            in3 => \N__23043\,
            lcout => n2976,
            ltout => OPEN,
            carryin => n12847,
            carryout => n12848,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_28_lut_LC_2_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28086\,
            in2 => \N__54284\,
            in3 => \N__23040\,
            lcout => n2975,
            ltout => OPEN,
            carryin => n12848,
            carryout => n12849,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_29_lut_LC_2_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54091\,
            in1 => \N__27311\,
            in2 => \N__32306\,
            in3 => \N__23037\,
            lcout => n3006,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i6_4_lut_LC_2_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__23033\,
            in1 => \N__23021\,
            in2 => \N__23010\,
            in3 => \N__22994\,
            lcout => \debounce.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12653_1_lut_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33895\,
            lcout => n15378,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i7_4_lut_LC_2_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__23297\,
            in1 => \N__23285\,
            in2 => \N__23274\,
            in3 => \N__23252\,
            lcout => \debounce.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1976_3_lut_LC_2_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27336\,
            in2 => \N__23241\,
            in3 => \N__33896\,
            lcout => n3008,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1592_3_lut_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25122\,
            in2 => \N__28458\,
            in3 => \N__32813\,
            lcout => n2432,
            ltout => \n2432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9978_3_lut_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37817\,
            in2 => \N__23214\,
            in3 => \N__23207\,
            lcout => OPEN,
            ltout => \n11946_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_114_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__23192\,
            in1 => \N__23170\,
            in2 => \N__23151\,
            in3 => \N__23143\,
            lcout => n13816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1589_3_lut_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29873\,
            in1 => \_gnd_net_\,
            in2 => \N__25317\,
            in3 => \N__32817\,
            lcout => n2429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1587_3_lut_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25262\,
            in1 => \_gnd_net_\,
            in2 => \N__32828\,
            in3 => \N__25245\,
            lcout => n2427,
            ltout => \n2427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_111_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23095\,
            in1 => \N__23368\,
            in2 => \N__23079\,
            in3 => \N__23075\,
            lcout => n14612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_129_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__23446\,
            in1 => \N__23833\,
            in2 => \N__24106\,
            in3 => \N__23433\,
            lcout => n13790,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_123_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23314\,
            in1 => \N__23524\,
            in2 => \N__23427\,
            in3 => \N__23382\,
            lcout => OPEN,
            ltout => \n14622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13070_4_lut_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23507\,
            in1 => \N__25514\,
            in2 => \N__23418\,
            in3 => \N__23415\,
            lcout => n2445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1580_3_lut_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25404\,
            in2 => \N__28755\,
            in3 => \N__32798\,
            lcout => n2420,
            ltout => \n2420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_113_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23341\,
            in2 => \N__23391\,
            in3 => \N__23388\,
            lcout => n14616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1586_3_lut_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25236\,
            in2 => \N__25485\,
            in3 => \N__32793\,
            lcout => n2426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1581_3_lut_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30056\,
            in2 => \N__32822\,
            in3 => \N__25413\,
            lcout => n2421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1583_3_lut_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25434\,
            in2 => \N__29817\,
            in3 => \N__32794\,
            lcout => n2423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1573_3_lut_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25533\,
            in1 => \_gnd_net_\,
            in2 => \N__32823\,
            in3 => \N__25503\,
            lcout => n2413,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1585_3_lut_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32805\,
            in1 => \_gnd_net_\,
            in2 => \N__25227\,
            in3 => \N__25460\,
            lcout => n2425,
            ltout => \n2425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_112_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23581\,
            in1 => \N__23623\,
            in2 => \N__23607\,
            in3 => \N__23704\,
            lcout => n14632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1579_3_lut_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25619\,
            in2 => \N__32824\,
            in3 => \N__25395\,
            lcout => n2419,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1575_3_lut_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32806\,
            in2 => \N__32511\,
            in3 => \N__25353\,
            lcout => n2415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_110_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32500\,
            in1 => \N__25636\,
            in2 => \N__30251\,
            in3 => \N__23730\,
            lcout => OPEN,
            ltout => \n14456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13043_4_lut_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28162\,
            in1 => \N__25501\,
            in2 => \N__23544\,
            in3 => \N__28389\,
            lcout => n2346,
            ltout => \n2346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1577_3_lut_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25637\,
            in2 => \N__23541\,
            in3 => \N__25374\,
            lcout => n2417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1574_3_lut_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25542\,
            in2 => \N__28167\,
            in3 => \N__32807\,
            lcout => n2414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_130_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24024\,
            in1 => \N__23755\,
            in2 => \N__23484\,
            in3 => \N__23472\,
            lcout => n14324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1521_3_lut_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28338\,
            in2 => \N__28236\,
            in3 => \N__32664\,
            lcout => n2329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1520_3_lut_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__28221\,
            in1 => \N__30003\,
            in2 => \N__32682\,
            in3 => \_gnd_net_\,
            lcout => n2328,
            ltout => \n2328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_107_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28744\,
            in1 => \N__29701\,
            in2 => \N__23739\,
            in3 => \N__29815\,
            lcout => OPEN,
            ltout => \n14442_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_108_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25585\,
            in1 => \N__25615\,
            in2 => \N__23736\,
            in3 => \N__25440\,
            lcout => OPEN,
            ltout => \n14448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_109_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__25297\,
            in1 => \N__29872\,
            in2 => \N__23733\,
            in3 => \N__28683\,
            lcout => n14450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1721_3_lut_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23654\,
            in2 => \N__23724\,
            in3 => \N__33119\,
            lcout => n2625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1649_3_lut_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23712\,
            in2 => \N__32998\,
            in3 => \N__23688\,
            lcout => n2521,
            ltout => \n2521_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_125_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23887\,
            in1 => \N__23653\,
            in2 => \N__23640\,
            in3 => \N__25654\,
            lcout => n14312,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_131_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24280\,
            in1 => \N__24130\,
            in2 => \N__23988\,
            in3 => \N__23975\,
            lcout => OPEN,
            ltout => \n14330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13099_4_lut_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23964\,
            in1 => \N__23929\,
            in2 => \N__23916\,
            in3 => \N__23913\,
            lcout => n2544,
            ltout => \n2544_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1718_rep_16_3_lut_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23888\,
            in2 => \N__23874\,
            in3 => \N__23871\,
            lcout => n2622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1719_3_lut_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25655\,
            in2 => \N__23862\,
            in3 => \N__33120\,
            lcout => n2623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1725_3_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23849\,
            in2 => \N__23817\,
            in3 => \N__33114\,
            lcout => n2629,
            ltout => \n2629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_140_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__26530\,
            in1 => \N__28482\,
            in2 => \N__23799\,
            in3 => \N__23796\,
            lcout => n14658,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1729_3_lut_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23790\,
            in1 => \N__28669\,
            in2 => \_gnd_net_\,
            in3 => \N__33110\,
            lcout => n2633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1782_3_lut_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26177\,
            in2 => \N__26157\,
            in3 => \N__33343\,
            lcout => n2718,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1712_3_lut_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23775\,
            in2 => \N__33156\,
            in3 => \N__23765\,
            lcout => n2616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1710_3_lut_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24153\,
            in2 => \N__24144\,
            in3 => \N__33118\,
            lcout => n2614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1726_3_lut_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__24114\,
            in1 => \N__24081\,
            in2 => \N__33155\,
            in3 => \_gnd_net_\,
            lcout => n2630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1791_3_lut_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25940\,
            in1 => \_gnd_net_\,
            in2 => \N__33328\,
            in3 => \N__25920\,
            lcout => n2727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1796_3_lut_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25566\,
            in2 => \N__28535\,
            in3 => \N__33273\,
            lcout => n2732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1780_3_lut_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26085\,
            in1 => \_gnd_net_\,
            in2 => \N__33329\,
            in3 => \N__26099\,
            lcout => n2716,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1713_3_lut_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24036\,
            in2 => \N__33165\,
            in3 => \N__24023\,
            lcout => n2617,
            ltout => \n2617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_141_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26075\,
            in1 => \N__23997\,
            in2 => \N__23991\,
            in3 => \N__26125\,
            lcout => n14664,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1788_3_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25833\,
            in1 => \N__25812\,
            in2 => \_gnd_net_\,
            in3 => \N__33278\,
            lcout => n2724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1789_3_lut_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25842\,
            in2 => \N__25866\,
            in3 => \N__33274\,
            lcout => n2725,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1781_3_lut_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26109\,
            in2 => \N__26145\,
            in3 => \N__33301\,
            lcout => n2717,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1792_3_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25971\,
            in1 => \_gnd_net_\,
            in2 => \N__33339\,
            in3 => \N__25953\,
            lcout => n2728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1709_3_lut_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24291\,
            in2 => \N__24264\,
            in3 => \N__33148\,
            lcout => n2613,
            ltout => \n2613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_142_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26032\,
            in1 => \N__25997\,
            in2 => \N__24249\,
            in3 => \N__24246\,
            lcout => OPEN,
            ltout => \n14670_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13130_4_lut_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26408\,
            in1 => \N__26368\,
            in2 => \N__24240\,
            in3 => \N__26321\,
            lcout => n2643,
            ltout => \n2643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1777_3_lut_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25980\,
            in1 => \_gnd_net_\,
            in2 => \N__24237\,
            in3 => \N__25998\,
            lcout => n2713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1720_rep_14_3_lut_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24213\,
            in2 => \N__25785\,
            in3 => \N__33296\,
            lcout => OPEN,
            ltout => \n14889_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1787_3_lut_4_lut_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__33297\,
            in1 => \N__33166\,
            in2 => \N__24192\,
            in3 => \N__24189\,
            lcout => n2723,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1779_3_lut_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26055\,
            in1 => \_gnd_net_\,
            in2 => \N__33341\,
            in3 => \N__26076\,
            lcout => n2715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1790_3_lut_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25908\,
            in2 => \N__25884\,
            in3 => \N__33302\,
            lcout => n2726,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1785_3_lut_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25713\,
            in1 => \_gnd_net_\,
            in2 => \N__33340\,
            in3 => \N__25734\,
            lcout => n2721,
            ltout => \n2721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_146_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24367\,
            in1 => \N__24328\,
            in2 => \N__24501\,
            in3 => \N__26646\,
            lcout => OPEN,
            ltout => \n14140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_147_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24493\,
            in1 => \N__24469\,
            in2 => \N__24450\,
            in3 => \N__24447\,
            lcout => OPEN,
            ltout => \n14146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_149_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24427\,
            in1 => \N__24400\,
            in2 => \N__24384\,
            in3 => \N__26445\,
            lcout => n14152,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1786_3_lut_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25746\,
            in2 => \N__25770\,
            in3 => \N__33303\,
            lcout => n2722,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1851_3_lut_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26736\,
            in2 => \N__33515\,
            in3 => \N__24351\,
            lcout => n2819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1859_3_lut_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24342\,
            in2 => \N__33512\,
            in3 => \N__24333\,
            lcout => n2827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1776_3_lut_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26439\,
            in1 => \N__26424\,
            in2 => \_gnd_net_\,
            in3 => \N__33334\,
            lcout => n2712,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1856_3_lut_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24651\,
            in1 => \_gnd_net_\,
            in2 => \N__33513\,
            in3 => \N__24624\,
            lcout => n2824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1774_3_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26375\,
            in2 => \N__26346\,
            in3 => \N__33335\,
            lcout => n2710,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12515_3_lut_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24612\,
            in1 => \_gnd_net_\,
            in2 => \N__33514\,
            in3 => \N__24600\,
            lcout => n2820,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1857_3_lut_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26717\,
            in2 => \N__24591\,
            in3 => \N__33470\,
            lcout => n2825,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1921_3_lut_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__24536\,
            in1 => \_gnd_net_\,
            in2 => \N__24579\,
            in3 => \N__33646\,
            lcout => n2921,
            ltout => \n2921_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_43_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27544\,
            in1 => \N__27673\,
            in2 => \N__24567\,
            in3 => \N__24784\,
            lcout => n14346,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1920_3_lut_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24515\,
            in2 => \N__24564\,
            in3 => \N__33645\,
            lcout => n2920,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1855_3_lut_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26697\,
            in1 => \_gnd_net_\,
            in2 => \N__24552\,
            in3 => \N__33463\,
            lcout => n2823,
            ltout => \n2823_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_28_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24535\,
            in1 => \N__25024\,
            in2 => \N__24522\,
            in3 => \N__24514\,
            lcout => n14690,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1841_3_lut_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24921\,
            in1 => \_gnd_net_\,
            in2 => \N__24915\,
            in3 => \N__33464\,
            lcout => n2809,
            ltout => \n2809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12625_4_lut_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24871\,
            in1 => \N__24842\,
            in2 => \N__24831\,
            in3 => \N__24828\,
            lcout => n2841,
            ltout => \n2841_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1922_3_lut_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24818\,
            in1 => \_gnd_net_\,
            in2 => \N__24804\,
            in3 => \N__24801\,
            lcout => n2922,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1987_3_lut_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24788\,
            in2 => \N__24768\,
            in3 => \N__33845\,
            lcout => n3019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1930_3_lut_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24756\,
            in2 => \N__24744\,
            in3 => \N__33655\,
            lcout => n2930,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1911_3_lut_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24714\,
            in2 => \N__33698\,
            in3 => \N__24705\,
            lcout => n2911,
            ltout => \n2911_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_48_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28024\,
            in1 => \N__27709\,
            in2 => \N__24687\,
            in3 => \N__26961\,
            lcout => n14372,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1928_3_lut_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24684\,
            in2 => \N__33697\,
            in3 => \N__24663\,
            lcout => n2928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1925_3_lut_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25044\,
            in2 => \N__25032\,
            in3 => \N__33651\,
            lcout => n2925,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1914_3_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__33656\,
            in1 => \_gnd_net_\,
            in2 => \N__25008\,
            in3 => \N__24996\,
            lcout => n2914,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1912_3_lut_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24972\,
            in2 => \N__24954\,
            in3 => \N__33657\,
            lcout => n2912,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_2_lut_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42225\,
            in2 => \_gnd_net_\,
            in3 => \N__24939\,
            lcout => n3101,
            ltout => OPEN,
            carryin => \bfn_3_29_0_\,
            carryout => n12850,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_3_lut_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53714\,
            in2 => \N__29118\,
            in3 => \N__24936\,
            lcout => n3100,
            ltout => OPEN,
            carryin => n12850,
            carryout => n12851,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_4_lut_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29097\,
            in3 => \N__24933\,
            lcout => n3099,
            ltout => OPEN,
            carryin => n12851,
            carryout => n12852,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_5_lut_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53715\,
            in2 => \N__29400\,
            in3 => \N__24930\,
            lcout => n3098,
            ltout => OPEN,
            carryin => n12852,
            carryout => n12853,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_6_lut_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29052\,
            in3 => \N__24927\,
            lcout => n3097,
            ltout => OPEN,
            carryin => n12853,
            carryout => n12854,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_7_lut_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29037\,
            in3 => \N__24924\,
            lcout => n3096,
            ltout => OPEN,
            carryin => n12854,
            carryout => n12855,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_8_lut_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53717\,
            in2 => \N__29235\,
            in3 => \N__25071\,
            lcout => n3095,
            ltout => OPEN,
            carryin => n12855,
            carryout => n12856,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_9_lut_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53716\,
            in2 => \N__28877\,
            in3 => \N__25068\,
            lcout => n3094,
            ltout => OPEN,
            carryin => n12856,
            carryout => n12857,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_10_lut_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31385\,
            in2 => \N__54456\,
            in3 => \N__25065\,
            lcout => n3093,
            ltout => OPEN,
            carryin => \bfn_3_30_0_\,
            carryout => n12858,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_11_lut_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54345\,
            in2 => \N__29475\,
            in3 => \N__25062\,
            lcout => n3092,
            ltout => OPEN,
            carryin => n12858,
            carryout => n12859,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_12_lut_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54352\,
            in2 => \N__37269\,
            in3 => \N__25059\,
            lcout => n3091,
            ltout => OPEN,
            carryin => n12859,
            carryout => n12860,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_13_lut_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54346\,
            in2 => \N__31169\,
            in3 => \N__25056\,
            lcout => n3090,
            ltout => OPEN,
            carryin => n12860,
            carryout => n12861,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_14_lut_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29264\,
            in2 => \N__54457\,
            in3 => \N__25053\,
            lcout => n3089,
            ltout => OPEN,
            carryin => n12861,
            carryout => n12862,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_15_lut_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54350\,
            in2 => \N__31496\,
            in3 => \N__25050\,
            lcout => n3088,
            ltout => OPEN,
            carryin => n12862,
            carryout => n12863,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_16_lut_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54353\,
            in2 => \N__27405\,
            in3 => \N__25047\,
            lcout => n3087,
            ltout => OPEN,
            carryin => n12863,
            carryout => n12864,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_17_lut_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54351\,
            in2 => \N__27579\,
            in3 => \N__25098\,
            lcout => n3086,
            ltout => OPEN,
            carryin => n12864,
            carryout => n12865,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_18_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29540\,
            in2 => \N__54264\,
            in3 => \N__25095\,
            lcout => n3085,
            ltout => OPEN,
            carryin => \bfn_3_31_0_\,
            carryout => n12866,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_19_lut_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29504\,
            in2 => \N__54268\,
            in3 => \N__25092\,
            lcout => n3084,
            ltout => OPEN,
            carryin => n12866,
            carryout => n12867,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_20_lut_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27641\,
            in2 => \N__54265\,
            in3 => \N__25089\,
            lcout => n3083,
            ltout => OPEN,
            carryin => n12867,
            carryout => n12868,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_21_lut_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29313\,
            in2 => \N__54269\,
            in3 => \N__25086\,
            lcout => n3082,
            ltout => OPEN,
            carryin => n12868,
            carryout => n12869,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_22_lut_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29171\,
            in2 => \N__54266\,
            in3 => \N__25083\,
            lcout => n3081,
            ltout => OPEN,
            carryin => n12869,
            carryout => n12870,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_23_lut_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34331\,
            in2 => \N__54270\,
            in3 => \N__25080\,
            lcout => n3080,
            ltout => OPEN,
            carryin => n12870,
            carryout => n12871,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_24_lut_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29570\,
            in2 => \N__54267\,
            in3 => \N__25077\,
            lcout => n3079,
            ltout => OPEN,
            carryin => n12871,
            carryout => n12872,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_25_lut_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29207\,
            in2 => \N__54271\,
            in3 => \N__25074\,
            lcout => n3078,
            ltout => OPEN,
            carryin => n12872,
            carryout => n12873,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_26_lut_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29753\,
            in2 => \N__54281\,
            in3 => \N__25200\,
            lcout => n3077,
            ltout => OPEN,
            carryin => \bfn_3_32_0_\,
            carryout => n12874,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_27_lut_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29666\,
            in2 => \N__54276\,
            in3 => \N__25197\,
            lcout => n3076,
            ltout => OPEN,
            carryin => n12874,
            carryout => n12875,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_28_lut_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29623\,
            in2 => \N__54282\,
            in3 => \N__25194\,
            lcout => n3075,
            ltout => OPEN,
            carryin => n12875,
            carryout => n12876,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_29_lut_LC_3_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29649\,
            in2 => \N__54277\,
            in3 => \N__25191\,
            lcout => n3074,
            ltout => OPEN,
            carryin => n12876,
            carryout => n12877,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_30_lut_LC_3_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54078\,
            in1 => \N__29597\,
            in2 => \N__32336\,
            in3 => \N__25188\,
            lcout => n3105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i9_4_lut_LC_3_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__25185\,
            in1 => \N__25167\,
            in2 => \N__25161\,
            in3 => \N__25140\,
            lcout => n14125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i2_LC_3_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27996\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \reg_B_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_2_lut_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30578\,
            in2 => \_gnd_net_\,
            in3 => \N__25125\,
            lcout => n2401,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => n12682,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_3_lut_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28454\,
            in2 => \N__54505\,
            in3 => \N__25113\,
            lcout => n2400,
            ltout => OPEN,
            carryin => n12682,
            carryout => n12683,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_4_lut_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30099\,
            in3 => \N__25335\,
            lcout => n2399,
            ltout => OPEN,
            carryin => n12683,
            carryout => n12684,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_5_lut_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28712\,
            in2 => \N__54506\,
            in3 => \N__25320\,
            lcout => n2398,
            ltout => OPEN,
            carryin => n12684,
            carryout => n12685,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_6_lut_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29874\,
            in3 => \N__25308\,
            lcout => n2397,
            ltout => OPEN,
            carryin => n12685,
            carryout => n12686,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_7_lut_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25305\,
            in3 => \N__25266\,
            lcout => n2396,
            ltout => OPEN,
            carryin => n12686,
            carryout => n12687,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_8_lut_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54413\,
            in2 => \N__25263\,
            in3 => \N__25239\,
            lcout => n2395,
            ltout => OPEN,
            carryin => n12687,
            carryout => n12688,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_9_lut_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54414\,
            in2 => \N__25484\,
            in3 => \N__25230\,
            lcout => n2394,
            ltout => OPEN,
            carryin => n12688,
            carryout => n12689,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_10_lut_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54519\,
            in2 => \N__25461\,
            in3 => \N__25218\,
            lcout => n2393,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => n12690,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_11_lut_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54526\,
            in2 => \N__28139\,
            in3 => \N__25203\,
            lcout => n2392,
            ltout => OPEN,
            carryin => n12690,
            carryout => n12691,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_12_lut_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54520\,
            in2 => \N__29816\,
            in3 => \N__25428\,
            lcout => n2391,
            ltout => OPEN,
            carryin => n12691,
            carryout => n12692,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_13_lut_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54527\,
            in2 => \N__29702\,
            in3 => \N__25416\,
            lcout => n2390,
            ltout => OPEN,
            carryin => n12692,
            carryout => n12693,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_14_lut_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54521\,
            in2 => \N__30057\,
            in3 => \N__25407\,
            lcout => n2389,
            ltout => OPEN,
            carryin => n12693,
            carryout => n12694,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_15_lut_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54528\,
            in2 => \N__28754\,
            in3 => \N__25398\,
            lcout => n2388,
            ltout => OPEN,
            carryin => n12694,
            carryout => n12695,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_16_lut_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54522\,
            in2 => \N__25623\,
            in3 => \N__25389\,
            lcout => n2387,
            ltout => OPEN,
            carryin => n12695,
            carryout => n12696,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_17_lut_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25592\,
            in2 => \N__54543\,
            in3 => \N__25377\,
            lcout => n2386,
            ltout => OPEN,
            carryin => n12696,
            carryout => n12697,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_18_lut_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54096\,
            in2 => \N__25641\,
            in3 => \N__25368\,
            lcout => n2385,
            ltout => OPEN,
            carryin => \bfn_4_19_0_\,
            carryout => n12698,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_19_lut_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53916\,
            in2 => \N__30252\,
            in3 => \N__25356\,
            lcout => n2384,
            ltout => OPEN,
            carryin => n12698,
            carryout => n12699,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_20_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54097\,
            in2 => \N__32507\,
            in3 => \N__25545\,
            lcout => n2383,
            ltout => OPEN,
            carryin => n12699,
            carryout => n12700,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_21_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53917\,
            in2 => \N__28166\,
            in3 => \N__25536\,
            lcout => n2382,
            ltout => OPEN,
            carryin => n12700,
            carryout => n12701,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_22_lut_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25502\,
            in2 => \N__54184\,
            in3 => \N__25527\,
            lcout => n2381,
            ltout => OPEN,
            carryin => n12701,
            carryout => n12702,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_23_lut_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54098\,
            in1 => \N__28388\,
            in2 => \N__32846\,
            in3 => \N__25524\,
            lcout => n2412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1506_3_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28407\,
            in2 => \N__32685\,
            in3 => \N__29925\,
            lcout => n2314_adj_622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1518_3_lut_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30451\,
            in2 => \N__28197\,
            in3 => \N__32676\,
            lcout => n2326,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13040_1_lut_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32808\,
            lcout => n15765,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1519_3_lut_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30507\,
            in2 => \N__28209\,
            in3 => \N__32656\,
            lcout => n2327,
            ltout => \n2327_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_106_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30046\,
            in1 => \N__28132\,
            in2 => \N__25464\,
            in3 => \N__25456\,
            lcout => n14440,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1652_3_lut_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25701\,
            in2 => \N__25685\,
            in3 => \N__32966\,
            lcout => n2524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1510_3_lut_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28266\,
            in2 => \N__32681\,
            in3 => \N__30153\,
            lcout => n2318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1512_3_lut_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28284\,
            in1 => \_gnd_net_\,
            in2 => \N__30357\,
            in3 => \N__32660\,
            lcout => n2320,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1511_3_lut_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28275\,
            in1 => \_gnd_net_\,
            in2 => \N__32680\,
            in3 => \N__30327\,
            lcout => n2319,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_2_lut_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40117\,
            in2 => \_gnd_net_\,
            in3 => \N__25569\,
            lcout => n2701,
            ltout => OPEN,
            carryin => \bfn_4_21_0_\,
            carryout => n12748,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_3_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54460\,
            in2 => \N__28534\,
            in3 => \N__25557\,
            lcout => n2700,
            ltout => OPEN,
            carryin => n12748,
            carryout => n12749,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_4_lut_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28503\,
            in2 => \_gnd_net_\,
            in3 => \N__25554\,
            lcout => n2699,
            ltout => OPEN,
            carryin => n12749,
            carryout => n12750,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_5_lut_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28551\,
            in2 => \N__54518\,
            in3 => \N__25551\,
            lcout => n2698,
            ltout => OPEN,
            carryin => n12750,
            carryout => n12751,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_6_lut_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26537\,
            in3 => \N__25548\,
            lcout => n2697,
            ltout => OPEN,
            carryin => n12751,
            carryout => n12752,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_7_lut_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25970\,
            in3 => \N__25944\,
            lcout => n2696,
            ltout => OPEN,
            carryin => n12752,
            carryout => n12753,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_8_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54465\,
            in2 => \N__25941\,
            in3 => \N__25911\,
            lcout => n2695,
            ltout => OPEN,
            carryin => n12753,
            carryout => n12754,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_9_lut_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54461\,
            in2 => \N__25904\,
            in3 => \N__25869\,
            lcout => n2694,
            ltout => OPEN,
            carryin => n12754,
            carryout => n12755,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_10_lut_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25865\,
            in2 => \N__53187\,
            in3 => \N__25836\,
            lcout => n2693,
            ltout => OPEN,
            carryin => \bfn_4_22_0_\,
            carryout => n12756,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_11_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25829\,
            in2 => \N__53191\,
            in3 => \N__25806\,
            lcout => n2692,
            ltout => OPEN,
            carryin => n12756,
            carryout => n12757,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_12_lut_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25803\,
            in2 => \N__53188\,
            in3 => \N__25773\,
            lcout => n2691,
            ltout => OPEN,
            carryin => n12757,
            carryout => n12758,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_13_lut_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25763\,
            in2 => \N__53192\,
            in3 => \N__25737\,
            lcout => n2690,
            ltout => OPEN,
            carryin => n12758,
            carryout => n12759,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_14_lut_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25730\,
            in2 => \N__53189\,
            in3 => \N__25704\,
            lcout => n2689,
            ltout => OPEN,
            carryin => n12759,
            carryout => n12760,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_15_lut_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26249\,
            in2 => \N__53193\,
            in3 => \N__26223\,
            lcout => n2688,
            ltout => OPEN,
            carryin => n12760,
            carryout => n12761,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_16_lut_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26220\,
            in2 => \N__53190\,
            in3 => \N__26184\,
            lcout => n2687,
            ltout => OPEN,
            carryin => n12761,
            carryout => n12762,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_17_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26181\,
            in2 => \N__53194\,
            in3 => \N__26148\,
            lcout => n2686,
            ltout => OPEN,
            carryin => n12762,
            carryout => n12763,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_18_lut_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26138\,
            in2 => \N__54092\,
            in3 => \N__26103\,
            lcout => n2685,
            ltout => OPEN,
            carryin => \bfn_4_23_0_\,
            carryout => n12764,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_19_lut_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53818\,
            in2 => \N__26100\,
            in3 => \N__26079\,
            lcout => n2684,
            ltout => OPEN,
            carryin => n12764,
            carryout => n12765,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_20_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26074\,
            in2 => \N__54093\,
            in3 => \N__26046\,
            lcout => n2683,
            ltout => OPEN,
            carryin => n12765,
            carryout => n12766,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_21_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26039\,
            in2 => \N__54176\,
            in3 => \N__26001\,
            lcout => n2682,
            ltout => OPEN,
            carryin => n12766,
            carryout => n12767,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_22_lut_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25996\,
            in2 => \N__54094\,
            in3 => \N__25974\,
            lcout => n2681,
            ltout => OPEN,
            carryin => n12767,
            carryout => n12768,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_23_lut_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26435\,
            in2 => \N__54177\,
            in3 => \N__26415\,
            lcout => n2680,
            ltout => OPEN,
            carryin => n12768,
            carryout => n12769,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_24_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26412\,
            in2 => \N__54095\,
            in3 => \N__26379\,
            lcout => n2679,
            ltout => OPEN,
            carryin => n12769,
            carryout => n12770,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_25_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26376\,
            in2 => \N__54178\,
            in3 => \N__26331\,
            lcout => n2678,
            ltout => OPEN,
            carryin => n12770,
            carryout => n12771,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_26_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53814\,
            in1 => \N__33362\,
            in2 => \N__26328\,
            in3 => \N__26301\,
            lcout => n2709,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13066_1_lut_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32987\,
            lcout => n15791,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i13_3_lut_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38697\,
            in1 => \N__46200\,
            in2 => \_gnd_net_\,
            in3 => \N__36609\,
            lcout => n307,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13127_1_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33345\,
            in3 => \_gnd_net_\,
            lcout => n15852,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1915_3_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26283\,
            in2 => \N__26265\,
            in3 => \N__33709\,
            lcout => n2915,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1784_3_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26250\,
            in2 => \N__26748\,
            in3 => \N__33321\,
            lcout => n2720,
            ltout => \n2720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_143_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26713\,
            in1 => \N__26689\,
            in2 => \N__26673\,
            in3 => \N__26662\,
            lcout => n14136,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1795_3_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28502\,
            in2 => \N__26640\,
            in3 => \N__33310\,
            lcout => n2731,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1794_3_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28550\,
            in2 => \N__33342\,
            in3 => \N__26625\,
            lcout => n2730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_27_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27868\,
            in1 => \N__26779\,
            in2 => \N__30697\,
            in3 => \N__27091\,
            lcout => OPEN,
            ltout => \n14688_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_29_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26605\,
            in1 => \N__26818\,
            in2 => \N__26589\,
            in3 => \N__26586\,
            lcout => n14696,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_new_i0_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26568\,
            lcout => \quad_counter0.b_new_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55775\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1793_3_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26550\,
            in2 => \N__26541\,
            in3 => \N__33314\,
            lcout => n2729,
            ltout => \n2729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_148_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__26497\,
            in1 => \N__26467\,
            in2 => \N__26448\,
            in3 => \N__26868\,
            lcout => n13796,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2062_3_lut_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28878\,
            in2 => \N__26955\,
            in3 => \N__37210\,
            lcout => n3126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1797_3_lut_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26940\,
            in1 => \N__40125\,
            in2 => \_gnd_net_\,
            in3 => \N__33330\,
            lcout => n2733,
            ltout => \n2733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9968_3_lut_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44871\,
            in2 => \N__26904\,
            in3 => \N__26894\,
            lcout => n11936,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12585_1_lut_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33511\,
            lcout => n15310,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1860_3_lut_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26855\,
            in1 => \_gnd_net_\,
            in2 => \N__26841\,
            in3 => \N__33510\,
            lcout => n2828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1918_3_lut_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26822\,
            in2 => \N__26802\,
            in3 => \N__33662\,
            lcout => n2918,
            ltout => \n2918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28975\,
            in2 => \N__26790\,
            in3 => \N__27367\,
            lcout => n14350,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1926_3_lut_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26783\,
            in2 => \N__26763\,
            in3 => \N__33663\,
            lcout => n2926,
            ltout => \n2926_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_42_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27120\,
            in3 => \N__27193\,
            lcout => OPEN,
            ltout => \n14336_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_44_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30664\,
            in1 => \N__27117\,
            in2 => \N__27111\,
            in3 => \N__27833\,
            lcout => OPEN,
            ltout => \n14352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_45_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27469\,
            in1 => \N__29360\,
            in2 => \N__27108\,
            in3 => \N__27105\,
            lcout => n14358,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1927_3_lut_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27095\,
            in2 => \N__27075\,
            in3 => \N__33661\,
            lcout => n2927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1917_3_lut_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27060\,
            in1 => \_gnd_net_\,
            in2 => \N__33699\,
            in3 => \N__27048\,
            lcout => n2917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1913_3_lut_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27021\,
            in1 => \_gnd_net_\,
            in2 => \N__27012\,
            in3 => \N__33676\,
            lcout => n2913,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_46_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__27160\,
            in1 => \N__27283\,
            in2 => \N__26985\,
            in3 => \N__26970\,
            lcout => OPEN,
            ltout => \n14360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_47_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27610\,
            in1 => \N__27790\,
            in2 => \N__26964\,
            in3 => \N__27751\,
            lcout => n14366,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i0_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34874\,
            lcout => \reg_B_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1994_3_lut_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27371\,
            in2 => \N__27351\,
            in3 => \N__33795\,
            lcout => n3026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12657_4_lut_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27334\,
            in1 => \N__28075\,
            in2 => \N__27315\,
            in3 => \N__27291\,
            lcout => n2940,
            ltout => \n2940_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1996_3_lut_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27284\,
            in1 => \_gnd_net_\,
            in2 => \N__27264\,
            in3 => \N__27261\,
            lcout => n3028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1988_3_lut_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27248\,
            in2 => \N__33850\,
            in3 => \N__27228\,
            lcout => n3020,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2051_3_lut_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27642\,
            in2 => \N__37223\,
            in3 => \N__27216\,
            lcout => n3115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1995_3_lut_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27207\,
            in1 => \_gnd_net_\,
            in2 => \N__33849\,
            in3 => \N__27197\,
            lcout => n3027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1997_3_lut_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27177\,
            in2 => \N__27168\,
            in3 => \N__33803\,
            lcout => n3029,
            ltout => \n3029_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2064_3_lut_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27144\,
            in2 => \N__27138\,
            in3 => \N__37211\,
            lcout => n3128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1991_3_lut_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27829\,
            in2 => \N__27135\,
            in3 => \N__33804\,
            lcout => n3023,
            ltout => \n3023_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_68_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27400\,
            in1 => \N__27571\,
            in2 => \N__27555\,
            in3 => \N__28851\,
            lcout => n14738,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1989_3_lut_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27552\,
            in2 => \N__27528\,
            in3 => \N__33796\,
            lcout => n3021,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2046_3_lut_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37153\,
            in1 => \_gnd_net_\,
            in2 => \N__27513\,
            in3 => \N__29208\,
            lcout => n3110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2043_3_lut_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27504\,
            in2 => \N__29637\,
            in3 => \N__37154\,
            lcout => n3107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1984_3_lut_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27495\,
            in2 => \N__27483\,
            in3 => \N__33858\,
            lcout => n3016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1998_3_lut_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27453\,
            in2 => \N__27429\,
            in3 => \N__33854\,
            lcout => n3030,
            ltout => \n3030_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2065_3_lut_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27414\,
            in2 => \N__27408\,
            in3 => \N__37149\,
            lcout => n3129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2055_3_lut_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27404\,
            in2 => \N__37203\,
            in3 => \N__27384\,
            lcout => n3119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1985_3_lut_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27945\,
            in1 => \_gnd_net_\,
            in2 => \N__33887\,
            in3 => \N__27932\,
            lcout => n3017,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1978_3_lut_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27912\,
            in1 => \N__27894\,
            in2 => \_gnd_net_\,
            in3 => \N__33873\,
            lcout => n3010,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1924_3_lut_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__27884\,
            in1 => \_gnd_net_\,
            in2 => \N__27852\,
            in3 => \N__33705\,
            lcout => n2924,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1980_3_lut_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27800\,
            in2 => \N__27774\,
            in3 => \N__33871\,
            lcout => n3012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1982_3_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27761\,
            in2 => \N__27732\,
            in3 => \N__33867\,
            lcout => n3014,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1979_3_lut_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__27720\,
            in1 => \N__27696\,
            in2 => \N__33891\,
            in3 => \_gnd_net_\,
            lcout => n3011,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1986_3_lut_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27687\,
            in2 => \N__27657\,
            in3 => \N__33872\,
            lcout => n3018,
            ltout => \n3018_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_164_LC_4_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27640\,
            in2 => \N__27624\,
            in3 => \N__29170\,
            lcout => n14816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1981_3_lut_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27621\,
            in2 => \N__27594\,
            in3 => \N__33892\,
            lcout => n3013,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12687_1_lut_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37171\,
            lcout => n15412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1975_3_lut_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28085\,
            in2 => \N__28056\,
            in3 => \N__33894\,
            lcout => n3007,
            ltout => \n3007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2042_3_lut_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28044\,
            in2 => \N__28038\,
            in3 => \N__37172\,
            lcout => n3106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1977_3_lut_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28035\,
            in2 => \N__28008\,
            in3 => \N__33893\,
            lcout => n3009,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i3_4_lut_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111111"
        )
    port map (
            in0 => \N__39554\,
            in1 => \N__27995\,
            in2 => \N__34809\,
            in3 => \N__39516\,
            lcout => \debounce.cnt_next_9__N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_2_lut_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32184\,
            in2 => \_gnd_net_\,
            in3 => \N__27954\,
            lcout => n2201,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => n12643,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_3_lut_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54403\,
            in2 => \N__32214\,
            in3 => \N__27951\,
            lcout => n2200,
            ltout => OPEN,
            carryin => n12643,
            carryout => n12644,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_4_lut_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32460\,
            in3 => \N__27948\,
            lcout => n2199,
            ltout => OPEN,
            carryin => n12644,
            carryout => n12645,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_5_lut_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54404\,
            in2 => \N__31970\,
            in3 => \N__28116\,
            lcout => n2198,
            ltout => OPEN,
            carryin => n12645,
            carryout => n12646,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_6_lut_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31998\,
            in3 => \N__28113\,
            lcout => n2197,
            ltout => OPEN,
            carryin => n12646,
            carryout => n12647,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_7_lut_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31936\,
            in3 => \N__28110\,
            lcout => n2196,
            ltout => OPEN,
            carryin => n12647,
            carryout => n12648,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_8_lut_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54406\,
            in2 => \N__31823\,
            in3 => \N__28107\,
            lcout => n2195,
            ltout => OPEN,
            carryin => n12648,
            carryout => n12649,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_9_lut_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54405\,
            in2 => \N__32289\,
            in3 => \N__28104\,
            lcout => n2194,
            ltout => OPEN,
            carryin => n12649,
            carryout => n12650,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_10_lut_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53562\,
            in2 => \N__31644\,
            in3 => \N__28101\,
            lcout => n2193,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => n12651,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_11_lut_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53571\,
            in2 => \N__31848\,
            in3 => \N__28098\,
            lcout => n2192,
            ltout => OPEN,
            carryin => n12651,
            carryout => n12652,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_12_lut_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53563\,
            in2 => \N__31599\,
            in3 => \N__28095\,
            lcout => n2191,
            ltout => OPEN,
            carryin => n12652,
            carryout => n12653,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_13_lut_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53572\,
            in2 => \N__31670\,
            in3 => \N__28092\,
            lcout => n2190,
            ltout => OPEN,
            carryin => n12653,
            carryout => n12654,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_14_lut_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53564\,
            in2 => \N__31869\,
            in3 => \N__28089\,
            lcout => n2189,
            ltout => OPEN,
            carryin => n12654,
            carryout => n12655,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_15_lut_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31752\,
            in2 => \N__53933\,
            in3 => \N__28188\,
            lcout => n2188,
            ltout => OPEN,
            carryin => n12655,
            carryout => n12656,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_16_lut_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31793\,
            in2 => \N__53935\,
            in3 => \N__28185\,
            lcout => n2187,
            ltout => OPEN,
            carryin => n12656,
            carryout => n12657,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_17_lut_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31904\,
            in2 => \N__53934\,
            in3 => \N__28182\,
            lcout => n2186,
            ltout => OPEN,
            carryin => n12657,
            carryout => n12658,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_18_lut_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32061\,
            in2 => \N__54181\,
            in3 => \N__28179\,
            lcout => n2185,
            ltout => OPEN,
            carryin => \bfn_5_19_0_\,
            carryout => n12659,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_19_lut_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29957\,
            in2 => \N__54183\,
            in3 => \N__28176\,
            lcout => n2184,
            ltout => OPEN,
            carryin => n12659,
            carryout => n12660,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_20_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30030\,
            in2 => \N__54182\,
            in3 => \N__28173\,
            lcout => n2183,
            ltout => OPEN,
            carryin => n12660,
            carryout => n12661,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_21_lut_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53915\,
            in1 => \N__34184\,
            in2 => \N__31698\,
            in3 => \N__28170\,
            lcout => n2214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1507_3_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29939\,
            in1 => \_gnd_net_\,
            in2 => \N__32655\,
            in3 => \N__28419\,
            lcout => n2315,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1517_3_lut_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32250\,
            in2 => \N__28311\,
            in3 => \N__32614\,
            lcout => n2325,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1451_3_lut_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28257\,
            in2 => \N__31824\,
            in3 => \N__34127\,
            lcout => n2227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_2_lut_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32036\,
            in2 => \_gnd_net_\,
            in3 => \N__28248\,
            lcout => n2301,
            ltout => OPEN,
            carryin => \bfn_5_20_0_\,
            carryout => n12662,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_3_lut_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53902\,
            in2 => \N__32145\,
            in3 => \N__28245\,
            lcout => n2300,
            ltout => OPEN,
            carryin => n12662,
            carryout => n12663,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_4_lut_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32097\,
            in3 => \N__28242\,
            lcout => n2299,
            ltout => OPEN,
            carryin => n12663,
            carryout => n12664,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_5_lut_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53903\,
            in2 => \N__32123\,
            in3 => \N__28239\,
            lcout => n2298,
            ltout => OPEN,
            carryin => n12664,
            carryout => n12665,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_6_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28334\,
            in2 => \_gnd_net_\,
            in3 => \N__28224\,
            lcout => n2297,
            ltout => OPEN,
            carryin => n12665,
            carryout => n12666,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_7_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30002\,
            in3 => \N__28212\,
            lcout => n2296,
            ltout => OPEN,
            carryin => n12666,
            carryout => n12667,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_8_lut_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53905\,
            in2 => \N__30506\,
            in3 => \N__28200\,
            lcout => n2295,
            ltout => OPEN,
            carryin => n12667,
            carryout => n12668,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_9_lut_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53904\,
            in2 => \N__30453\,
            in3 => \N__28314\,
            lcout => n2294,
            ltout => OPEN,
            carryin => n12668,
            carryout => n12669,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_10_lut_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53890\,
            in2 => \N__32249\,
            in3 => \N__28299\,
            lcout => n2293,
            ltout => OPEN,
            carryin => \bfn_5_21_0_\,
            carryout => n12670,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_11_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53896\,
            in2 => \N__30426\,
            in3 => \N__28296\,
            lcout => n2292,
            ltout => OPEN,
            carryin => n12670,
            carryout => n12671,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_12_lut_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53891\,
            in2 => \N__30474\,
            in3 => \N__28293\,
            lcout => n2291,
            ltout => OPEN,
            carryin => n12671,
            carryout => n12672,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_13_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53897\,
            in2 => \N__30405\,
            in3 => \N__28290\,
            lcout => n2290,
            ltout => OPEN,
            carryin => n12672,
            carryout => n12673,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_14_lut_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53892\,
            in2 => \N__30381\,
            in3 => \N__28287\,
            lcout => n2289,
            ltout => OPEN,
            carryin => n12673,
            carryout => n12674,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_15_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53898\,
            in2 => \N__30353\,
            in3 => \N__28278\,
            lcout => n2288,
            ltout => OPEN,
            carryin => n12674,
            carryout => n12675,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_16_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30320\,
            in2 => \N__54180\,
            in3 => \N__28269\,
            lcout => n2287,
            ltout => OPEN,
            carryin => n12675,
            carryout => n12676,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_17_lut_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30146\,
            in2 => \N__54179\,
            in3 => \N__28260\,
            lcout => n2286,
            ltout => OPEN,
            carryin => n12676,
            carryout => n12677,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_18_lut_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53491\,
            in2 => \N__30177\,
            in3 => \N__28425\,
            lcout => n2285,
            ltout => OPEN,
            carryin => \bfn_5_22_0_\,
            carryout => n12678,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_19_lut_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32522\,
            in2 => \N__53888\,
            in3 => \N__28422\,
            lcout => n2284,
            ltout => OPEN,
            carryin => n12678,
            carryout => n12679,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_20_lut_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29940\,
            in2 => \N__53921\,
            in3 => \N__28410\,
            lcout => n2283,
            ltout => OPEN,
            carryin => n12679,
            carryout => n12680,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_21_lut_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29924\,
            in2 => \N__53889\,
            in3 => \N__28395\,
            lcout => n2282,
            ltout => OPEN,
            carryin => n12680,
            carryout => n12681,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_22_lut_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__53546\,
            in1 => \N__29901\,
            in2 => \N__32702\,
            in3 => \N__28392\,
            lcout => n2313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1523_3_lut_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28368\,
            in2 => \N__32671\,
            in3 => \N__32096\,
            lcout => n2331,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1452_3_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28359\,
            in2 => \N__31944\,
            in3 => \N__34159\,
            lcout => n2228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1454_3_lut_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28347\,
            in2 => \N__31977\,
            in3 => \N__34160\,
            lcout => n2230,
            ltout => \n2230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_103_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__30001\,
            in1 => \_gnd_net_\,
            in2 => \N__28317\,
            in3 => \_gnd_net_\,
            lcout => n14812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1513_3_lut_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30380\,
            in1 => \_gnd_net_\,
            in2 => \N__32684\,
            in3 => \N__28764\,
            lcout => n2321,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9986_4_lut_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__30565\,
            in1 => \N__30077\,
            in2 => \N__28705\,
            in3 => \N__28441\,
            lcout => n11954,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i9_3_lut_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38499\,
            in1 => \N__46182\,
            in2 => \_gnd_net_\,
            in3 => \N__36666\,
            lcout => n311,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1728_3_lut_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28638\,
            in2 => \N__28605\,
            in3 => \N__33163\,
            lcout => n2632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36665\,
            lcout => n25_adj_646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1727_3_lut_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28590\,
            in2 => \N__28566\,
            in3 => \N__33164\,
            lcout => n2631,
            ltout => \n2631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10076_4_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__40121\,
            in1 => \N__28536\,
            in2 => \N__28506\,
            in3 => \N__28498\,
            lcout => n12044,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1525_3_lut_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__32037\,
            in1 => \_gnd_net_\,
            in2 => \N__28470\,
            in3 => \N__32672\,
            lcout => n2333,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36570\,
            lcout => n20_adj_641,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_2_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40054\,
            in2 => \_gnd_net_\,
            in3 => \N__28791\,
            lcout => n3201,
            ltout => OPEN,
            carryin => \bfn_5_25_0_\,
            carryout => n12878,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_3_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53251\,
            in2 => \N__36933\,
            in3 => \N__28788\,
            lcout => n3200,
            ltout => OPEN,
            carryin => n12878,
            carryout => n12879,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_4_lut_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36906\,
            in3 => \N__28785\,
            lcout => n3199,
            ltout => OPEN,
            carryin => n12879,
            carryout => n12880,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_5_lut_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53252\,
            in2 => \N__36798\,
            in3 => \N__28782\,
            lcout => n3198,
            ltout => OPEN,
            carryin => n12880,
            carryout => n12881,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_6_lut_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36836\,
            in3 => \N__28779\,
            lcout => n3197,
            ltout => OPEN,
            carryin => n12881,
            carryout => n12882,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_7_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36876\,
            in3 => \N__28776\,
            lcout => n3196,
            ltout => OPEN,
            carryin => n12882,
            carryout => n12883,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_8_lut_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53254\,
            in2 => \N__34545\,
            in3 => \N__28773\,
            lcout => n3195,
            ltout => OPEN,
            carryin => n12883,
            carryout => n12884,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_9_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53253\,
            in2 => \N__34361\,
            in3 => \N__28770\,
            lcout => n3194,
            ltout => OPEN,
            carryin => n12884,
            carryout => n12885,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_10_lut_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53003\,
            in2 => \N__34243\,
            in3 => \N__28767\,
            lcout => n3193,
            ltout => OPEN,
            carryin => \bfn_5_26_0_\,
            carryout => n12886,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_11_lut_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53008\,
            in2 => \N__34920\,
            in3 => \N__28818\,
            lcout => n3192,
            ltout => OPEN,
            carryin => n12886,
            carryout => n12887,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_12_lut_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30953\,
            in2 => \N__53386\,
            in3 => \N__28815\,
            lcout => n3191,
            ltout => OPEN,
            carryin => n12887,
            carryout => n12888,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_13_lut_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53012\,
            in2 => \N__37044\,
            in3 => \N__28812\,
            lcout => n3190,
            ltout => OPEN,
            carryin => n12888,
            carryout => n12889,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_14_lut_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31138\,
            in2 => \N__53387\,
            in3 => \N__28809\,
            lcout => n3189,
            ltout => OPEN,
            carryin => n12889,
            carryout => n12890,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_15_lut_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53016\,
            in2 => \N__31005\,
            in3 => \N__28806\,
            lcout => n3188,
            ltout => OPEN,
            carryin => n12890,
            carryout => n12891,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_16_lut_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53004\,
            in2 => \N__31458\,
            in3 => \N__28803\,
            lcout => n3187,
            ltout => OPEN,
            carryin => n12891,
            carryout => n12892,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_17_lut_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34457\,
            in2 => \N__53385\,
            in3 => \N__28800\,
            lcout => n3186,
            ltout => OPEN,
            carryin => n12892,
            carryout => n12893,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_18_lut_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34780\,
            in2 => \N__54286\,
            in3 => \N__28797\,
            lcout => n3185,
            ltout => OPEN,
            carryin => \bfn_5_27_0_\,
            carryout => n12894,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_19_lut_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54102\,
            in2 => \N__34496\,
            in3 => \N__28794\,
            lcout => n3184,
            ltout => OPEN,
            carryin => n12894,
            carryout => n12895,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_20_lut_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30755\,
            in2 => \N__54287\,
            in3 => \N__28845\,
            lcout => n3183,
            ltout => OPEN,
            carryin => n12895,
            carryout => n12896,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_21_lut_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31076\,
            in2 => \N__54290\,
            in3 => \N__28842\,
            lcout => n3182,
            ltout => OPEN,
            carryin => n12896,
            carryout => n12897,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_22_lut_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31050\,
            in2 => \N__54288\,
            in3 => \N__28839\,
            lcout => n3181,
            ltout => OPEN,
            carryin => n12897,
            carryout => n12898,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_23_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30921\,
            in2 => \N__54291\,
            in3 => \N__28836\,
            lcout => n3180,
            ltout => OPEN,
            carryin => n12898,
            carryout => n12899,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_24_lut_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34956\,
            in2 => \N__54289\,
            in3 => \N__28833\,
            lcout => n3179,
            ltout => OPEN,
            carryin => n12899,
            carryout => n12900,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_25_lut_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31201\,
            in2 => \N__54292\,
            in3 => \N__28830\,
            lcout => n3178,
            ltout => OPEN,
            carryin => n12900,
            carryout => n12901,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_26_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54121\,
            in2 => \N__34292\,
            in3 => \N__28827\,
            lcout => n3177,
            ltout => OPEN,
            carryin => \bfn_5_28_0_\,
            carryout => n12902,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_27_lut_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43226\,
            in2 => \N__54293\,
            in3 => \N__28824\,
            lcout => n3176,
            ltout => OPEN,
            carryin => n12902,
            carryout => n12903,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_28_lut_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30893\,
            in2 => \N__54295\,
            in3 => \N__28821\,
            lcout => n3175,
            ltout => OPEN,
            carryin => n12903,
            carryout => n12904,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_29_lut_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30816\,
            in2 => \N__54294\,
            in3 => \N__29007\,
            lcout => n3174,
            ltout => OPEN,
            carryin => n12904,
            carryout => n12905,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_30_lut_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30848\,
            in2 => \N__54296\,
            in3 => \N__29004\,
            lcout => n3173,
            ltout => OPEN,
            carryin => n12905,
            carryout => n12906,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_31_lut_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__30873\,
            in1 => \N__54134\,
            in2 => \N__32366\,
            in3 => \N__29001\,
            lcout => n3204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2116_3_lut_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30919\,
            in2 => \N__28998\,
            in3 => \N__43146\,
            lcout => n3212,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1992_3_lut_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28985\,
            in2 => \N__28959\,
            in3 => \N__33844\,
            lcout => n3024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2067_3_lut_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29093\,
            in1 => \_gnd_net_\,
            in2 => \N__28944\,
            in3 => \N__37193\,
            lcout => n3131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2044_3_lut_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__37195\,
            in1 => \_gnd_net_\,
            in2 => \N__28932\,
            in3 => \N__29673\,
            lcout => n3108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1993_3_lut_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28913\,
            in2 => \N__28893\,
            in3 => \N__33865\,
            lcout => n3025,
            ltout => \n3025_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_67_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37255\,
            in1 => \N__28870\,
            in2 => \N__28854\,
            in3 => \N__29058\,
            lcout => n14736,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2049_3_lut_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29175\,
            in2 => \N__29154\,
            in3 => \N__37194\,
            lcout => n3113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2068_3_lut_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29114\,
            in2 => \N__37217\,
            in3 => \N__29139\,
            lcout => n3132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2001_3_lut_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__32425\,
            in1 => \_gnd_net_\,
            in2 => \N__29130\,
            in3 => \N__33866\,
            lcout => n3033,
            ltout => \n3033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9964_3_lut_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__42220\,
            in1 => \_gnd_net_\,
            in2 => \N__29100\,
            in3 => \N__29092\,
            lcout => n11932,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1990_3_lut_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30672\,
            in2 => \N__29073\,
            in3 => \N__33862\,
            lcout => n3022,
            ltout => \n3022_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_66_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29233\,
            in1 => \N__31489\,
            in2 => \N__29061\,
            in3 => \N__31384\,
            lcout => n14732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_69_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__29048\,
            in1 => \N__29033\,
            in2 => \N__29396\,
            in3 => \N__29022\,
            lcout => OPEN,
            ltout => \n13859_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_70_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29306\,
            in1 => \N__29503\,
            in2 => \N__29016\,
            in3 => \N__29013\,
            lcout => n14744,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1999_3_lut_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29436\,
            in2 => \N__29424\,
            in3 => \N__33863\,
            lcout => n3031,
            ltout => \n3031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2066_3_lut_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29376\,
            in2 => \N__29364\,
            in3 => \N__37155\,
            lcout => n3130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1983_3_lut_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29361\,
            in2 => \N__29328\,
            in3 => \N__33864\,
            lcout => n3015,
            ltout => \n3015_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2050_3_lut_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29295\,
            in2 => \N__29283\,
            in3 => \N__37156\,
            lcout => n3114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2057_3_lut_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29280\,
            in2 => \N__29268\,
            in3 => \N__37158\,
            lcout => n3121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2063_3_lut_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29247\,
            in2 => \N__37204\,
            in3 => \N__29234\,
            lcout => n3127,
            ltout => \n3127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_32_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34444\,
            in1 => \N__34534\,
            in2 => \N__29211\,
            in3 => \N__34245\,
            lcout => n14196,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_101_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29206\,
            in1 => \N__34330\,
            in2 => \N__29571\,
            in3 => \N__29190\,
            lcout => OPEN,
            ltout => \n14750_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_165_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29184\,
            in1 => \N__29752\,
            in2 => \N__29178\,
            in3 => \N__29665\,
            lcout => OPEN,
            ltout => \n14754_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12690_4_lut_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29648\,
            in1 => \N__29633\,
            in2 => \N__29604\,
            in3 => \N__29601\,
            lcout => n3039,
            ltout => \n3039_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2047_3_lut_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29583\,
            in2 => \N__29574\,
            in3 => \N__29569\,
            lcout => n3111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_30_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30946\,
            in1 => \N__34906\,
            in2 => \N__34782\,
            in3 => \N__31140\,
            lcout => OPEN,
            ltout => \n14194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_33_LC_5_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29514\,
            in1 => \N__30748\,
            in2 => \N__29553\,
            in3 => \N__29550\,
            lcout => n14204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2053_3_lut_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29544\,
            in1 => \_gnd_net_\,
            in2 => \N__37205\,
            in3 => \N__29529\,
            lcout => n3117,
            ltout => \n3117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_31_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30988\,
            in1 => \N__31441\,
            in2 => \N__29517\,
            in3 => \N__37039\,
            lcout => n14198,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2052_3_lut_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29508\,
            in2 => \N__37206\,
            in3 => \N__29487\,
            lcout => n3116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2060_3_lut_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29474\,
            in2 => \N__29451\,
            in3 => \N__37162\,
            lcout => n3124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2045_3_lut_LC_5_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29757\,
            in1 => \_gnd_net_\,
            in2 => \N__29736\,
            in3 => \N__37169\,
            lcout => n3109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1385_3_lut_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31410\,
            in2 => \N__37974\,
            in3 => \N__34024\,
            lcout => n2129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12989_1_lut_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34169\,
            in3 => \_gnd_net_\,
            lcout => n15714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1387_3_lut_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31422\,
            in2 => \N__38118\,
            in3 => \N__34025\,
            lcout => n2131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36608\,
            lcout => n21_adj_642,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1384_3_lut_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31401\,
            in2 => \N__36174\,
            in3 => \N__33985\,
            lcout => n2128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1448_3_lut_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__31847\,
            in1 => \_gnd_net_\,
            in2 => \N__29724\,
            in3 => \N__34154\,
            lcout => n2224,
            ltout => \n2224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1515_3_lut_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29715\,
            in2 => \N__29706\,
            in3 => \N__32653\,
            lcout => n2323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1382_3_lut_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31569\,
            in2 => \N__37677\,
            in3 => \N__33984\,
            lcout => n2126,
            ltout => \n2126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1449_3_lut_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29838\,
            in2 => \N__29832\,
            in3 => \N__34155\,
            lcout => n2225,
            ltout => \n2225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1516_3_lut_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29829\,
            in2 => \N__29820\,
            in3 => \N__32654\,
            lcout => n2324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1381_3_lut_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31560\,
            in2 => \N__36372\,
            in3 => \N__34002\,
            lcout => n2125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1372_3_lut_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36317\,
            in1 => \_gnd_net_\,
            in2 => \N__34027\,
            in3 => \N__31710\,
            lcout => n2116,
            ltout => \n2116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1439_3_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34153\,
            in1 => \_gnd_net_\,
            in2 => \N__29781\,
            in3 => \N__29778\,
            lcout => n2215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12967_4_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36316\,
            in1 => \N__36092\,
            in2 => \N__31629\,
            in3 => \N__36435\,
            lcout => n2049,
            ltout => \n2049_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1379_3_lut_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36203\,
            in2 => \N__29769\,
            in3 => \N__31548\,
            lcout => n2123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1442_3_lut_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31905\,
            in2 => \N__29766\,
            in3 => \N__34152\,
            lcout => n2218,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1376_3_lut_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31533\,
            in2 => \N__38028\,
            in3 => \N__34003\,
            lcout => n2120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1375_3_lut_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31524\,
            in2 => \N__34026\,
            in3 => \N__37886\,
            lcout => n2119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1514_3_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30403\,
            in2 => \N__30066\,
            in3 => \N__32613\,
            lcout => n2322,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1373_3_lut_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31628\,
            in2 => \N__31722\,
            in3 => \N__34015\,
            lcout => n2117,
            ltout => \n2117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12992_4_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31691\,
            in1 => \N__30029\,
            in2 => \N__30018\,
            in3 => \N__31884\,
            lcout => n2148,
            ltout => \n2148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1453_3_lut_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31991\,
            in2 => \N__30015\,
            in3 => \N__30012\,
            lcout => n2229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1445_3_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31862\,
            in2 => \N__29976\,
            in3 => \N__34148\,
            lcout => n2221,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1440_3_lut_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__29964\,
            in1 => \_gnd_net_\,
            in2 => \N__34168\,
            in3 => \N__29958\,
            lcout => n2216,
            ltout => \n2216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13017_4_lut_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29923\,
            in1 => \N__29897\,
            in2 => \N__29886\,
            in3 => \N__30126\,
            lcout => n2247,
            ltout => \n2247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1522_3_lut_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__29883\,
            in1 => \_gnd_net_\,
            in2 => \N__29877\,
            in3 => \N__32124\,
            lcout => n2330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1443_3_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__30285\,
            in1 => \_gnd_net_\,
            in2 => \N__34162\,
            in3 => \N__31797\,
            lcout => n2219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1455_3_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32453\,
            in2 => \N__30276\,
            in3 => \N__34128\,
            lcout => n2231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1509_3_lut_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__30173\,
            in1 => \_gnd_net_\,
            in2 => \N__30261\,
            in3 => \N__32635\,
            lcout => n2317,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1456_3_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32207\,
            in2 => \N__30216\,
            in3 => \N__34129\,
            lcout => n2232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1447_3_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31595\,
            in2 => \N__34161\,
            in3 => \N__30201\,
            lcout => n2223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1441_3_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32057\,
            in2 => \N__30192\,
            in3 => \N__34137\,
            lcout => n2217,
            ltout => \n2217_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_105_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30172\,
            in1 => \N__30145\,
            in2 => \N__30129\,
            in3 => \N__30291\,
            lcout => n14598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1444_3_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30120\,
            in2 => \N__31751\,
            in3 => \N__34133\,
            lcout => n2220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1524_3_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32138\,
            in2 => \N__30111\,
            in3 => \N__32636\,
            lcout => n2332,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1446_3_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__34163\,
            in1 => \N__31671\,
            in2 => \N__30522\,
            in3 => \_gnd_net_\,
            lcout => n2222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_99_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30499\,
            in3 => \N__30467\,
            lcout => OPEN,
            ltout => \n14578_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_100_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30452\,
            in1 => \N__32236\,
            in2 => \N__30429\,
            in3 => \N__30422\,
            lcout => OPEN,
            ltout => \n14582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_102_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30404\,
            in1 => \N__30376\,
            in2 => \N__30360\,
            in3 => \N__30352\,
            lcout => OPEN,
            ltout => \n14588_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_104_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__32076\,
            in1 => \N__30319\,
            in2 => \N__30303\,
            in3 => \N__30300\,
            lcout => n14592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13014_1_lut_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32637\,
            lcout => n15739,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41919\,
            in3 => \_gnd_net_\,
            lcout => n17_adj_638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12759_1_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32390\,
            lcout => n15484,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36718\,
            lcout => n19_adj_640,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i14_3_lut_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38661\,
            in1 => \N__46158\,
            in2 => \_gnd_net_\,
            in3 => \N__36569\,
            lcout => n306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i11_3_lut_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46159\,
            in1 => \N__38754\,
            in2 => \_gnd_net_\,
            in3 => \N__40007\,
            lcout => n309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12762_4_lut_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35754\,
            in1 => \N__30528\,
            in2 => \N__31347\,
            in3 => \N__30603\,
            lcout => n12034,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2198_3_lut_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35016\,
            in2 => \N__34992\,
            in3 => \N__34632\,
            lcout => OPEN,
            ltout => \n17_adj_710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_117_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__34633\,
            in1 => \N__35231\,
            in2 => \N__30543\,
            in3 => \N__35205\,
            lcout => n14236,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2197_3_lut_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35481\,
            in2 => \N__35457\,
            in3 => \N__34634\,
            lcout => OPEN,
            ltout => \n19_adj_711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_118_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__34635\,
            in1 => \N__35435\,
            in2 => \N__30540\,
            in3 => \N__35415\,
            lcout => OPEN,
            ltout => \n14230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_122_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30537\,
            in1 => \N__34254\,
            in2 => \N__30531\,
            in3 => \N__30615\,
            lcout => n14248,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2176_3_lut_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35820\,
            in1 => \N__35834\,
            in2 => \_gnd_net_\,
            in3 => \N__34656\,
            lcout => n61,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_152_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__35955\,
            in1 => \N__35969\,
            in2 => \N__34699\,
            in3 => \N__31296\,
            lcout => OPEN,
            ltout => \n14268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_153_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__35940\,
            in1 => \N__43006\,
            in2 => \N__30624\,
            in3 => \N__34655\,
            lcout => n14270,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_163_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35917\,
            in1 => \N__35968\,
            in2 => \N__43010\,
            in3 => \N__30726\,
            lcout => OPEN,
            ltout => \n14806_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12758_4_lut_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35875\,
            in1 => \N__35833\,
            in2 => \N__30621\,
            in3 => \N__35774\,
            lcout => n3237,
            ltout => \n3237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_115_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__35400\,
            in1 => \N__35376\,
            in2 => \N__30618\,
            in3 => \N__30774\,
            lcout => n14228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9894_4_lut_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__34565\,
            in1 => \N__35190\,
            in2 => \N__40563\,
            in3 => \N__34651\,
            lcout => n11861,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_154_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__35918\,
            in1 => \N__35898\,
            in2 => \N__34700\,
            in3 => \N__30609\,
            lcout => n14272,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2109_3_lut_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__30852\,
            in1 => \N__30597\,
            in2 => \N__43173\,
            in3 => \_gnd_net_\,
            lcout => n3205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2118_3_lut_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31077\,
            in2 => \N__30588\,
            in3 => \N__43152\,
            lcout => n3214,
            ltout => \n3214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_161_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35560\,
            in1 => \N__35618\,
            in2 => \N__30789\,
            in3 => \N__34389\,
            lcout => n14794,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2126_3_lut_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37043\,
            in2 => \N__30786\,
            in3 => \N__43150\,
            lcout => n3222,
            ltout => \n3222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2193_3_lut_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__35310\,
            in1 => \_gnd_net_\,
            in2 => \N__30777\,
            in3 => \N__34629\,
            lcout => n27_adj_713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2119_3_lut_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30768\,
            in2 => \N__30762\,
            in3 => \N__43151\,
            lcout => n3215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_162_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35524\,
            in1 => \N__36035\,
            in2 => \N__36013\,
            in3 => \N__30732\,
            lcout => n14800,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1923_3_lut_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30720\,
            in2 => \N__30711\,
            in3 => \N__33696\,
            lcout => n2923,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2123_3_lut_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30639\,
            in2 => \N__31457\,
            in3 => \N__43085\,
            lcout => n3219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2125_3_lut_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30633\,
            in2 => \N__43147\,
            in3 => \N__31139\,
            lcout => n3221,
            ltout => \n3221_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_155_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30627\,
            in3 => \N__35221\,
            lcout => n14764,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2111_3_lut_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31011\,
            in1 => \_gnd_net_\,
            in2 => \N__43149\,
            in3 => \N__30897\,
            lcout => n3207,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2124_3_lut_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31004\,
            in2 => \N__30972\,
            in3 => \N__43086\,
            lcout => n3220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2127_3_lut_LC_6_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30963\,
            in2 => \N__43148\,
            in3 => \N__30957\,
            lcout => n3223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2115_3_lut_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34952\,
            in2 => \N__30930\,
            in3 => \N__43093\,
            lcout => n3211,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_36_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31202\,
            in1 => \N__34948\,
            in2 => \N__30920\,
            in3 => \N__31017\,
            lcout => OPEN,
            ltout => \n14216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_37_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30892\,
            in1 => \N__34285\,
            in2 => \N__30876\,
            in3 => \N__43225\,
            lcout => OPEN,
            ltout => \n14222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12724_4_lut_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30814\,
            in1 => \N__30872\,
            in2 => \N__30855\,
            in3 => \N__30847\,
            lcout => n3138,
            ltout => \n3138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12720_1_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30819\,
            in3 => \_gnd_net_\,
            lcout => n15445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2110_3_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__30815\,
            in1 => \N__30795\,
            in2 => \N__43170\,
            in3 => \_gnd_net_\,
            lcout => n3206,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2137_3_lut_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31230\,
            in1 => \N__40055\,
            in2 => \_gnd_net_\,
            in3 => \N__43133\,
            lcout => n3233,
            ltout => \n3233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9958_4_lut_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__31215\,
            in1 => \N__35163\,
            in2 => \N__31206\,
            in3 => \N__34726\,
            lcout => n11926,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2114_3_lut_LC_6_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31203\,
            in2 => \N__31179\,
            in3 => \N__43134\,
            lcout => n3210,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2058_3_lut_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31170\,
            in2 => \N__37218\,
            in3 => \N__31152\,
            lcout => n3122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2117_3_lut_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31113\,
            in1 => \_gnd_net_\,
            in2 => \N__43172\,
            in3 => \N__31046\,
            lcout => n3213,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2135_3_lut_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36898\,
            in2 => \N__31104\,
            in3 => \N__43138\,
            lcout => n3231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2134_3_lut_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36787\,
            in2 => \N__43171\,
            in3 => \N__31089\,
            lcout => n3230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_35_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31072\,
            in1 => \N__31042\,
            in2 => \N__36768\,
            in3 => \N__31026\,
            lcout => n14210,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2069_3_lut_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31284\,
            in1 => \N__42224\,
            in2 => \_gnd_net_\,
            in3 => \N__37196\,
            lcout => n3133,
            ltout => \n3133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2136_3_lut_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31275\,
            in2 => \N__31263\,
            in3 => \N__43139\,
            lcout => n3232,
            ltout => \n3232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10062_4_lut_LC_6_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__40558\,
            in1 => \N__35174\,
            in2 => \N__31260\,
            in3 => \N__35125\,
            lcout => n12030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_119_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__35739\,
            in1 => \N__35718\,
            in2 => \N__34578\,
            in3 => \N__34703\,
            lcout => n14234,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16_4_lut_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__35127\,
            in1 => \N__35079\,
            in2 => \N__34728\,
            in3 => \N__35099\,
            lcout => n5_adj_703,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2188_3_lut_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35679\,
            in2 => \N__35709\,
            in3 => \N__34702\,
            lcout => n37_adj_715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2194_3_lut_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__35358\,
            in1 => \N__35337\,
            in2 => \N__34727\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n25_adj_712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_120_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__35025\,
            in1 => \N__35046\,
            in2 => \N__31257\,
            in3 => \N__34707\,
            lcout => OPEN,
            ltout => \n14238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_124_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31254\,
            in1 => \N__31248\,
            in2 => \N__31242\,
            in3 => \N__31239\,
            lcout => OPEN,
            ltout => \n14250_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_126_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__35670\,
            in1 => \N__35643\,
            in2 => \N__31392\,
            in3 => \N__34708\,
            lcout => n14252,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2061_3_lut_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31389\,
            in2 => \N__31362\,
            in3 => \N__37170\,
            lcout => n3125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2177_3_lut_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35879\,
            in2 => \N__34730\,
            in3 => \N__35850\,
            lcout => n59,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_132_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__34715\,
            in2 => \N__35634\,
            in3 => \N__31332\,
            lcout => OPEN,
            ltout => \n14254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_133_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__31305\,
            in1 => \N__31326\,
            in2 => \N__31320\,
            in3 => \N__31317\,
            lcout => OPEN,
            ltout => \n14256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_134_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__35597\,
            in1 => \N__35577\,
            in2 => \N__31308\,
            in3 => \N__34716\,
            lcout => n14258,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2203_3_lut_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35154\,
            in1 => \_gnd_net_\,
            in2 => \N__34729\,
            in3 => \N__35139\,
            lcout => n7_adj_708,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_150_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__36024\,
            in1 => \N__36051\,
            in2 => \N__34731\,
            in3 => \N__31506\,
            lcout => OPEN,
            ltout => \n14264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_151_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__36014\,
            in1 => \N__35982\,
            in2 => \N__31299\,
            in3 => \N__34725\,
            lcout => n14266,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_136_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__35568\,
            in1 => \N__34720\,
            in2 => \N__35538\,
            in3 => \N__31515\,
            lcout => OPEN,
            ltout => \n14260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_144_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__34721\,
            in1 => \N__35490\,
            in2 => \N__31509\,
            in3 => \N__35526\,
            lcout => n14262,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2056_3_lut_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31500\,
            in2 => \N__31473\,
            in3 => \N__37157\,
            lcout => n3120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_2_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38402\,
            in2 => \_gnd_net_\,
            in3 => \N__31428\,
            lcout => n2101,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => n12625,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_3_lut_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54399\,
            in2 => \N__38321\,
            in3 => \N__31425\,
            lcout => n2100,
            ltout => OPEN,
            carryin => n12625,
            carryout => n12626,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_4_lut_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38117\,
            in3 => \N__31416\,
            lcout => n2099,
            ltout => OPEN,
            carryin => n12626,
            carryout => n12627,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_5_lut_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54400\,
            in2 => \N__38427\,
            in3 => \N__31413\,
            lcout => n2098,
            ltout => OPEN,
            carryin => n12627,
            carryout => n12628,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_6_lut_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37973\,
            in3 => \N__31404\,
            lcout => n2097,
            ltout => OPEN,
            carryin => n12628,
            carryout => n12629,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_7_lut_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36173\,
            in3 => \N__31395\,
            lcout => n2096,
            ltout => OPEN,
            carryin => n12629,
            carryout => n12630,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_8_lut_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54402\,
            in2 => \N__38280\,
            in3 => \N__31572\,
            lcout => n2095,
            ltout => OPEN,
            carryin => n12630,
            carryout => n12631,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_9_lut_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54401\,
            in2 => \N__37676\,
            in3 => \N__31563\,
            lcout => n2094,
            ltout => OPEN,
            carryin => n12631,
            carryout => n12632,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_10_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54389\,
            in2 => \N__36371\,
            in3 => \N__31554\,
            lcout => n2093,
            ltout => OPEN,
            carryin => \bfn_7_18_0_\,
            carryout => n12633,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_11_lut_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53560\,
            in2 => \N__36273\,
            in3 => \N__31551\,
            lcout => n2092,
            ltout => OPEN,
            carryin => n12633,
            carryout => n12634,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_12_lut_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54390\,
            in2 => \N__36207\,
            in3 => \N__31542\,
            lcout => n2091,
            ltout => OPEN,
            carryin => n12634,
            carryout => n12635,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_13_lut_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53561\,
            in2 => \N__36414\,
            in3 => \N__31539\,
            lcout => n2090,
            ltout => OPEN,
            carryin => n12635,
            carryout => n12636,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_14_lut_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54391\,
            in2 => \N__36242\,
            in3 => \N__31536\,
            lcout => n2089,
            ltout => OPEN,
            carryin => n12636,
            carryout => n12637,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_15_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38024\,
            in2 => \N__54503\,
            in3 => \N__31527\,
            lcout => n2088,
            ltout => OPEN,
            carryin => n12637,
            carryout => n12638,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_16_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54395\,
            in2 => \N__37887\,
            in3 => \N__31518\,
            lcout => n2087,
            ltout => OPEN,
            carryin => n12638,
            carryout => n12639,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_17_lut_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36464\,
            in2 => \N__54504\,
            in3 => \N__31725\,
            lcout => n2086,
            ltout => OPEN,
            carryin => n12639,
            carryout => n12640,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_18_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31627\,
            in2 => \N__54459\,
            in3 => \N__31713\,
            lcout => n2085,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => n12641,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_19_lut_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36318\,
            in2 => \N__54502\,
            in3 => \N__31704\,
            lcout => n2084,
            ltout => OPEN,
            carryin => n12641,
            carryout => n12642,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_20_lut_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54365\,
            in1 => \N__36093\,
            in2 => \N__34046\,
            in3 => \N__31701\,
            lcout => n2115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1383_3_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38279\,
            in2 => \N__34016\,
            in3 => \N__31680\,
            lcout => n2127,
            ltout => \n2127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_94_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31663\,
            in1 => \N__31585\,
            in2 => \N__31647\,
            in3 => \N__31640\,
            lcout => n14384,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1306_3_lut_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39717\,
            in2 => \N__36117\,
            in3 => \N__38210\,
            lcout => n2018,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1380_3_lut_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36269\,
            in2 => \N__31608\,
            in3 => \N__33977\,
            lcout => n2124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12964_1_lut_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34017\,
            in3 => \_gnd_net_\,
            lcout => n15689,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1386_3_lut_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__38423\,
            in1 => \N__32007\,
            in2 => \N__34028\,
            in3 => \_gnd_net_\,
            lcout => n2130,
            ltout => \n2130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_97_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__31969\,
            in1 => \N__31940\,
            in2 => \N__31908\,
            in3 => \N__32190\,
            lcout => OPEN,
            ltout => \n13775_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_98_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31903\,
            in1 => \N__32053\,
            in2 => \N__31887\,
            in3 => \N__31767\,
            lcout => n14398,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1378_3_lut_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34011\,
            in1 => \N__31878\,
            in2 => \N__36413\,
            in3 => \_gnd_net_\,
            lcout => n2122,
            ltout => \n2122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_95_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31843\,
            in2 => \N__31827\,
            in3 => \N__31822\,
            lcout => OPEN,
            ltout => \n14386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_96_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31792\,
            in1 => \N__31741\,
            in2 => \N__31776\,
            in3 => \N__31773\,
            lcout => n14392,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1377_3_lut_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31761\,
            in2 => \N__36243\,
            in3 => \N__34010\,
            lcout => n2121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1450_3_lut_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32285\,
            in2 => \N__32265\,
            in3 => \N__34144\,
            lcout => n2226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1389_3_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32223\,
            in1 => \N__38398\,
            in2 => \_gnd_net_\,
            in3 => \N__34019\,
            lcout => n2133,
            ltout => \n2133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9925_3_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32182\,
            in2 => \N__32193\,
            in3 => \N__32449\,
            lcout => n11892,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1457_3_lut_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32183\,
            in1 => \_gnd_net_\,
            in2 => \N__34167\,
            in3 => \N__32157\,
            lcout => n2233,
            ltout => \n2233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9982_4_lut_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__32023\,
            in1 => \N__32116\,
            in2 => \N__32100\,
            in3 => \N__32092\,
            lcout => n11950,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1374_3_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32070\,
            in2 => \N__36468\,
            in3 => \N__34020\,
            lcout => n2118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37847\,
            lcout => n24_adj_645,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36633\,
            in1 => \N__38727\,
            in2 => \_gnd_net_\,
            in3 => \N__46160\,
            lcout => n308,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36632\,
            lcout => n22_adj_643,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1508_3_lut_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32535\,
            in2 => \N__32526\,
            in3 => \N__32652\,
            lcout => n2316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46164\,
            in1 => \N__36537\,
            in2 => \_gnd_net_\,
            in3 => \N__38079\,
            lcout => n319,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1388_3_lut_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32469\,
            in2 => \N__38322\,
            in3 => \N__34018\,
            lcout => n2132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36504\,
            in1 => \_gnd_net_\,
            in2 => \N__46195\,
            in3 => \N__38568\,
            lcout => n315,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i0_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__32397\,
            in1 => \N__42115\,
            in2 => \N__32391\,
            in3 => \N__32376\,
            lcout => encoder0_position_scaled_0,
            ltout => OPEN,
            carryin => \bfn_7_23_0_\,
            carryout => n12938,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i1_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35801\,
            in1 => \N__34701\,
            in2 => \N__42175\,
            in3 => \N__32373\,
            lcout => encoder0_position_scaled_1,
            ltout => OPEN,
            carryin => n12938,
            carryout => n12939,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i2_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__32370\,
            in1 => \N__43178\,
            in2 => \N__42178\,
            in3 => \N__32349\,
            lcout => encoder0_position_scaled_2,
            ltout => OPEN,
            carryin => n12939,
            carryout => n12940,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i3_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__32346\,
            in1 => \N__42128\,
            in2 => \N__37224\,
            in3 => \N__32319\,
            lcout => encoder0_position_scaled_3,
            ltout => OPEN,
            carryin => n12940,
            carryout => n12941,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i4_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__32316\,
            in1 => \N__33897\,
            in2 => \N__42179\,
            in3 => \N__33741\,
            lcout => encoder0_position_scaled_4,
            ltout => OPEN,
            carryin => n12941,
            carryout => n12942,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i5_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__33738\,
            in1 => \N__33714\,
            in2 => \N__42176\,
            in3 => \N__33555\,
            lcout => encoder0_position_scaled_5,
            ltout => OPEN,
            carryin => n12942,
            carryout => n12943,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i6_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__33552\,
            in1 => \N__33528\,
            in2 => \N__42180\,
            in3 => \N__33372\,
            lcout => encoder0_position_scaled_6,
            ltout => OPEN,
            carryin => n12943,
            carryout => n12944,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i7_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__33369\,
            in1 => \N__33350\,
            in2 => \N__42177\,
            in3 => \N__33198\,
            lcout => encoder0_position_scaled_7,
            ltout => OPEN,
            carryin => n12944,
            carryout => n12945,
            clk => \N__55778\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i8_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__33195\,
            in1 => \N__33171\,
            in2 => \N__42185\,
            in3 => \N__33027\,
            lcout => encoder0_position_scaled_8,
            ltout => OPEN,
            carryin => \bfn_7_24_0_\,
            carryout => n12946,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i9_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__33020\,
            in1 => \N__32999\,
            in2 => \N__42181\,
            in3 => \N__32853\,
            lcout => encoder0_position_scaled_9,
            ltout => OPEN,
            carryin => n12946,
            carryout => n12947,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i10_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__32850\,
            in1 => \N__32829\,
            in2 => \N__42186\,
            in3 => \N__32706\,
            lcout => encoder0_position_scaled_10,
            ltout => OPEN,
            carryin => n12947,
            carryout => n12948,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i11_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__32703\,
            in1 => \N__32683\,
            in2 => \N__42182\,
            in3 => \N__32538\,
            lcout => encoder0_position_scaled_11,
            ltout => OPEN,
            carryin => n12948,
            carryout => n12949,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i12_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34191\,
            in1 => \N__34170\,
            in2 => \N__42187\,
            in3 => \N__34053\,
            lcout => encoder0_position_scaled_12,
            ltout => OPEN,
            carryin => n12949,
            carryout => n12950,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i13_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34050\,
            in1 => \N__34029\,
            in2 => \N__42183\,
            in3 => \N__33921\,
            lcout => encoder0_position_scaled_13,
            ltout => OPEN,
            carryin => n12950,
            carryout => n12951,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i14_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37944\,
            in1 => \N__38217\,
            in2 => \N__42188\,
            in3 => \N__33918\,
            lcout => encoder0_position_scaled_14,
            ltout => OPEN,
            carryin => n12951,
            carryout => n12952,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i15_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39780\,
            in1 => \N__39888\,
            in2 => \N__42184\,
            in3 => \N__33915\,
            lcout => encoder0_position_scaled_15,
            ltout => OPEN,
            carryin => n12952,
            carryout => n12953,
            clk => \N__55779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i16_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__44550\,
            in1 => \N__41805\,
            in2 => \N__42171\,
            in3 => \N__33912\,
            lcout => encoder0_position_scaled_16,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => n12954,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i17_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47988\,
            in1 => \N__50202\,
            in2 => \N__42189\,
            in3 => \N__33909\,
            lcout => encoder0_position_scaled_17,
            ltout => OPEN,
            carryin => n12954,
            carryout => n12955,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i18_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45738\,
            in1 => \N__50676\,
            in2 => \N__42172\,
            in3 => \N__33906\,
            lcout => encoder0_position_scaled_18,
            ltout => OPEN,
            carryin => n12955,
            carryout => n12956,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i19_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__51324\,
            in1 => \N__51405\,
            in2 => \N__42190\,
            in3 => \N__33903\,
            lcout => encoder0_position_scaled_19,
            ltout => OPEN,
            carryin => n12956,
            carryout => n12957,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i20_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__48513\,
            in1 => \N__51300\,
            in2 => \N__42173\,
            in3 => \N__33900\,
            lcout => encoder0_position_scaled_20,
            ltout => OPEN,
            carryin => n12957,
            carryout => n12958,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i21_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__51531\,
            in1 => \N__51603\,
            in2 => \N__42191\,
            in3 => \N__34314\,
            lcout => encoder0_position_scaled_21,
            ltout => OPEN,
            carryin => n12958,
            carryout => n12959,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i22_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__52365\,
            in1 => \N__52275\,
            in2 => \N__42174\,
            in3 => \N__34311\,
            lcout => encoder0_position_scaled_22,
            ltout => OPEN,
            carryin => n12959,
            carryout => n12960,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i23_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46356\,
            in1 => \N__46425\,
            in2 => \N__42192\,
            in3 => \N__34308\,
            lcout => encoder0_position_scaled_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2113_3_lut_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34305\,
            in2 => \N__43174\,
            in3 => \N__34293\,
            lcout => n3209,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2191_3_lut_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__35261\,
            in1 => \_gnd_net_\,
            in2 => \N__35247\,
            in3 => \N__34630\,
            lcout => OPEN,
            ltout => \n31_adj_714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_116_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__34631\,
            in1 => \N__35291\,
            in2 => \N__34257\,
            in3 => \N__35277\,
            lcout => n14232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2129_3_lut_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34244\,
            in2 => \N__34215\,
            in3 => \N__43156\,
            lcout => n3225,
            ltout => \n3225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_156_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35008\,
            in1 => \N__35260\,
            in2 => \N__34203\,
            in3 => \N__35321\,
            lcout => OPEN,
            ltout => \n14776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_158_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35470\,
            in1 => \N__35350\,
            in2 => \N__34200\,
            in3 => \N__34197\,
            lcout => OPEN,
            ltout => \n14780_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_159_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34410\,
            in1 => \N__35659\,
            in2 => \N__34548\,
            in3 => \N__35704\,
            lcout => n14786,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2131_3_lut_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34544\,
            in2 => \N__34512\,
            in3 => \N__43125\,
            lcout => n3227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2120_3_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34497\,
            in2 => \N__43169\,
            in3 => \N__34467\,
            lcout => n3216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2122_3_lut_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34458\,
            in2 => \N__34428\,
            in3 => \N__43129\,
            lcout => n3218,
            ltout => \n3218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_157_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35392\,
            in2 => \N__34413\,
            in3 => \N__35041\,
            lcout => n14778,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_160_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__35100\,
            in1 => \N__34404\,
            in2 => \N__35070\,
            in3 => \N__34395\,
            lcout => n14788,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34383\,
            lcout => n13_adj_570,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2130_3_lut_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34374\,
            in2 => \N__43168\,
            in3 => \N__34362\,
            lcout => n3226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2048_3_lut_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34338\,
            in2 => \N__34971\,
            in3 => \N__37216\,
            lcout => n3112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2128_3_lut_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34932\,
            in2 => \N__43166\,
            in3 => \N__34916\,
            lcout => n3224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2132_3_lut_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36874\,
            in2 => \N__34890\,
            in3 => \N__43117\,
            lcout => n3228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12725_1_lut_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34664\,
            lcout => n15450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i2_4_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__34875\,
            in1 => \N__39426\,
            in2 => \N__34853\,
            in3 => \N__34824\,
            lcout => \debounce.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2121_3_lut_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34794\,
            in2 => \N__43167\,
            in3 => \N__34781\,
            lcout => n3217,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2133_3_lut_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36837\,
            in2 => \N__34749\,
            in3 => \N__43124\,
            lcout => n3229,
            ltout => \n3229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2200_3_lut_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35055\,
            in2 => \N__34734\,
            in3 => \N__34663\,
            lcout => n13_adj_709,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_2_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34566\,
            in2 => \N__53636\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_29_0_\,
            carryout => n12907,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40559\,
            in2 => \_gnd_net_\,
            in3 => \N__35178\,
            lcout => n3301,
            ltout => OPEN,
            carryin => n12907,
            carryout => n12908,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35175\,
            in2 => \N__53637\,
            in3 => \N__35157\,
            lcout => n3300,
            ltout => OPEN,
            carryin => n12908,
            carryout => n12909,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35150\,
            in2 => \_gnd_net_\,
            in3 => \N__35130\,
            lcout => n3299,
            ltout => OPEN,
            carryin => n12909,
            carryout => n12910,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35126\,
            in2 => \N__53638\,
            in3 => \N__35109\,
            lcout => n3298,
            ltout => OPEN,
            carryin => n12910,
            carryout => n12911,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__35106\,
            in1 => \N__35098\,
            in2 => \_gnd_net_\,
            in3 => \N__35073\,
            lcout => n15097,
            ltout => OPEN,
            carryin => n12911,
            carryout => n12912,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35069\,
            in2 => \_gnd_net_\,
            in3 => \N__35049\,
            lcout => n3296,
            ltout => OPEN,
            carryin => n12912,
            carryout => n12913,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35042\,
            in2 => \N__53639\,
            in3 => \N__35019\,
            lcout => n3295,
            ltout => OPEN,
            carryin => n12913,
            carryout => n12914,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35015\,
            in2 => \N__53987\,
            in3 => \N__34974\,
            lcout => n3294,
            ltout => OPEN,
            carryin => \bfn_7_30_0_\,
            carryout => n12915,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35477\,
            in2 => \N__54002\,
            in3 => \N__35439\,
            lcout => n3293,
            ltout => OPEN,
            carryin => n12915,
            carryout => n12916,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35436\,
            in2 => \N__53988\,
            in3 => \N__35403\,
            lcout => n3292,
            ltout => OPEN,
            carryin => n12916,
            carryout => n12917,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35399\,
            in2 => \N__54003\,
            in3 => \N__35361\,
            lcout => n3291,
            ltout => OPEN,
            carryin => n12917,
            carryout => n12918,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35357\,
            in2 => \N__53989\,
            in3 => \N__35331\,
            lcout => n3290,
            ltout => OPEN,
            carryin => n12918,
            carryout => n12919,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35328\,
            in2 => \N__54004\,
            in3 => \N__35298\,
            lcout => n3289,
            ltout => OPEN,
            carryin => n12919,
            carryout => n12920,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53694\,
            in2 => \N__35295\,
            in3 => \N__35268\,
            lcout => n3288,
            ltout => OPEN,
            carryin => n12920,
            carryout => n12921,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35265\,
            in2 => \N__54005\,
            in3 => \N__35235\,
            lcout => n3287,
            ltout => OPEN,
            carryin => n12921,
            carryout => n12922,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35232\,
            in2 => \N__53990\,
            in3 => \N__35193\,
            lcout => n3286,
            ltout => OPEN,
            carryin => \bfn_7_31_0_\,
            carryout => n12923,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35735\,
            in2 => \N__53994\,
            in3 => \N__35712\,
            lcout => n3285,
            ltout => OPEN,
            carryin => n12923,
            carryout => n12924,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35705\,
            in2 => \N__53991\,
            in3 => \N__35673\,
            lcout => n3284,
            ltout => OPEN,
            carryin => n12924,
            carryout => n12925,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35666\,
            in2 => \N__53995\,
            in3 => \N__35637\,
            lcout => n3283,
            ltout => OPEN,
            carryin => n12925,
            carryout => n12926,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35630\,
            in2 => \N__53992\,
            in3 => \N__35601\,
            lcout => n3282,
            ltout => OPEN,
            carryin => n12926,
            carryout => n12927,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35598\,
            in2 => \N__53996\,
            in3 => \N__35571\,
            lcout => n3281,
            ltout => OPEN,
            carryin => n12927,
            carryout => n12928,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35567\,
            in2 => \N__53993\,
            in3 => \N__35529\,
            lcout => n3280,
            ltout => OPEN,
            carryin => n12928,
            carryout => n12929,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35525\,
            in2 => \N__53997\,
            in3 => \N__35484\,
            lcout => n3279,
            ltout => OPEN,
            carryin => n12929,
            carryout => n12930,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36047\,
            in2 => \N__53998\,
            in3 => \N__36018\,
            lcout => n3278,
            ltout => OPEN,
            carryin => \bfn_7_32_0_\,
            carryout => n12931,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36015\,
            in2 => \N__54006\,
            in3 => \N__35976\,
            lcout => n3277,
            ltout => OPEN,
            carryin => n12931,
            carryout => n12932,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35973\,
            in2 => \N__53999\,
            in3 => \N__35943\,
            lcout => n3276,
            ltout => OPEN,
            carryin => n12932,
            carryout => n12933,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43011\,
            in2 => \N__54007\,
            in3 => \N__35928\,
            lcout => n3275,
            ltout => OPEN,
            carryin => n12933,
            carryout => n12934,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35925\,
            in2 => \N__54000\,
            in3 => \N__35883\,
            lcout => n3274,
            ltout => OPEN,
            carryin => n12934,
            carryout => n12935,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35880\,
            in2 => \N__54008\,
            in3 => \N__35844\,
            lcout => n3273,
            ltout => OPEN,
            carryin => n12935,
            carryout => n12936,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35841\,
            in2 => \N__54001\,
            in3 => \N__35805\,
            lcout => n3272,
            ltout => OPEN,
            carryin => n12936,
            carryout => n12937,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53707\,
            in1 => \N__35802\,
            in2 => \N__35781\,
            in3 => \N__35757\,
            lcout => n14873,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_2_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38359\,
            in2 => \_gnd_net_\,
            in3 => \N__36078\,
            lcout => n2001,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => n12608,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_3_lut_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38233\,
            in2 => \N__54360\,
            in3 => \N__36075\,
            lcout => n2000,
            ltout => OPEN,
            carryin => n12608,
            carryout => n12609,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_4_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38456\,
            in2 => \_gnd_net_\,
            in3 => \N__36072\,
            lcout => n1999,
            ltout => OPEN,
            carryin => n12609,
            carryout => n12610,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_5_lut_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54201\,
            in2 => \N__39954\,
            in3 => \N__36069\,
            lcout => n1998,
            ltout => OPEN,
            carryin => n12610,
            carryout => n12611,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_6_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39690\,
            in3 => \N__36066\,
            lcout => n1997,
            ltout => OPEN,
            carryin => n12611,
            carryout => n12612,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_7_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39662\,
            in3 => \N__36063\,
            lcout => n1996,
            ltout => OPEN,
            carryin => n12612,
            carryout => n12613,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_8_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54197\,
            in2 => \N__39618\,
            in3 => \N__36060\,
            lcout => n1995,
            ltout => OPEN,
            carryin => n12613,
            carryout => n12614,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_9_lut_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37787\,
            in2 => \N__54361\,
            in3 => \N__36057\,
            lcout => n1994,
            ltout => OPEN,
            carryin => n12614,
            carryout => n12615,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_10_lut_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53152\,
            in2 => \N__37748\,
            in3 => \N__36054\,
            lcout => n1993,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => n12616,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_11_lut_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53158\,
            in2 => \N__37641\,
            in3 => \N__36135\,
            lcout => n1992,
            ltout => OPEN,
            carryin => n12616,
            carryout => n12617,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_12_lut_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53153\,
            in2 => \N__37721\,
            in3 => \N__36132\,
            lcout => n1991,
            ltout => OPEN,
            carryin => n12617,
            carryout => n12618,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_13_lut_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53159\,
            in2 => \N__37769\,
            in3 => \N__36129\,
            lcout => n1990,
            ltout => OPEN,
            carryin => n12618,
            carryout => n12619,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_14_lut_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53154\,
            in2 => \N__38052\,
            in3 => \N__36126\,
            lcout => n1989,
            ltout => OPEN,
            carryin => n12619,
            carryout => n12620,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_15_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53160\,
            in2 => \N__37904\,
            in3 => \N__36123\,
            lcout => n1988,
            ltout => OPEN,
            carryin => n12620,
            carryout => n12621,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_16_lut_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39737\,
            in2 => \N__53559\,
            in3 => \N__36120\,
            lcout => n1987,
            ltout => OPEN,
            carryin => n12621,
            carryout => n12622,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_17_lut_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39716\,
            in2 => \N__53558\,
            in3 => \N__36102\,
            lcout => n1986,
            ltout => OPEN,
            carryin => n12622,
            carryout => n12623,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_18_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53452\,
            in2 => \N__39926\,
            in3 => \N__36099\,
            lcout => n1985,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => n12624,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_19_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53453\,
            in1 => \N__37937\,
            in2 => \N__37926\,
            in3 => \N__36096\,
            lcout => n2016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1313_3_lut_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36336\,
            in2 => \N__37752\,
            in3 => \N__38184\,
            lcout => n2025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1310_3_lut_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37770\,
            in2 => \N__38208\,
            in3 => \N__36330\,
            lcout => n2022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1305_3_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36324\,
            in2 => \N__39927\,
            in3 => \N__38195\,
            lcout => n2017,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1312_3_lut_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37639\,
            in2 => \N__38207\,
            in3 => \N__36297\,
            lcout => n2024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1317_3_lut_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39686\,
            in2 => \N__36291\,
            in3 => \N__38191\,
            lcout => n2029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1307_3_lut_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36279\,
            in2 => \N__38209\,
            in3 => \N__39741\,
            lcout => n2019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_90_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36352\,
            in1 => \N__36259\,
            in2 => \N__38269\,
            in3 => \N__37663\,
            lcout => OPEN,
            ltout => \n14550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_91_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36223\,
            in1 => \N__36199\,
            in2 => \N__36177\,
            in3 => \N__36397\,
            lcout => OPEN,
            ltout => \n14556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_92_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__36154\,
            in1 => \N__37966\,
            in2 => \N__36138\,
            in3 => \N__38367\,
            lcout => OPEN,
            ltout => \n14558_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_93_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37870\,
            in1 => \N__38011\,
            in2 => \N__36471\,
            in3 => \N__36451\,
            lcout => n14564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1311_3_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37722\,
            in1 => \_gnd_net_\,
            in2 => \N__38206\,
            in3 => \N__36423\,
            lcout => n2023,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1314_3_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36381\,
            in2 => \N__37797\,
            in3 => \N__38180\,
            lcout => n2026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42374\,
            lcout => n15_adj_636,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40579\,
            lcout => n32_adj_653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40072\,
            lcout => n31_adj_652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38977\,
            lcout => n28_adj_649,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36532\,
            lcout => n33_adj_654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44887\,
            lcout => n27_adj_648,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36499\,
            lcout => n29_adj_650,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40141\,
            lcout => n26_adj_647,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i0_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36536\,
            in2 => \_gnd_net_\,
            in3 => \N__36516\,
            lcout => encoder0_position_0,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \quad_counter0.n13025\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i1_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37367\,
            in2 => \N__40589\,
            in3 => \N__36513\,
            lcout => encoder0_position_1,
            ltout => OPEN,
            carryin => \quad_counter0.n13025\,
            carryout => \quad_counter0.n13026\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i2_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40076\,
            in2 => \N__37415\,
            in3 => \N__36510\,
            lcout => encoder0_position_2,
            ltout => OPEN,
            carryin => \quad_counter0.n13026\,
            carryout => \quad_counter0.n13027\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i3_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37371\,
            in2 => \N__42250\,
            in3 => \N__36507\,
            lcout => encoder0_position_3,
            ltout => OPEN,
            carryin => \quad_counter0.n13027\,
            carryout => \quad_counter0.n13028\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i4_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36503\,
            in2 => \N__37416\,
            in3 => \N__36483\,
            lcout => encoder0_position_4,
            ltout => OPEN,
            carryin => \quad_counter0.n13028\,
            carryout => \quad_counter0.n13029\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i5_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37375\,
            in2 => \N__38987\,
            in3 => \N__36480\,
            lcout => encoder0_position_5,
            ltout => OPEN,
            carryin => \quad_counter0.n13029\,
            carryout => \quad_counter0.n13030\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i6_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44891\,
            in2 => \N__37417\,
            in3 => \N__36477\,
            lcout => encoder0_position_6,
            ltout => OPEN,
            carryin => \quad_counter0.n13030\,
            carryout => \quad_counter0.n13031\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i7_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37379\,
            in2 => \N__40151\,
            in3 => \N__36474\,
            lcout => encoder0_position_7,
            ltout => OPEN,
            carryin => \quad_counter0.n13031\,
            carryout => \quad_counter0.n13032\,
            clk => \N__55780\,
            ce => \N__39117\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i8_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37380\,
            in2 => \N__36664\,
            in3 => \N__36642\,
            lcout => encoder0_position_8,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \quad_counter0.n13033\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i9_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37840\,
            in2 => \N__37418\,
            in3 => \N__36639\,
            lcout => encoder0_position_9,
            ltout => OPEN,
            carryin => \quad_counter0.n13033\,
            carryout => \quad_counter0.n13034\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i10_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37384\,
            in2 => \N__40008\,
            in3 => \N__36636\,
            lcout => encoder0_position_10,
            ltout => OPEN,
            carryin => \quad_counter0.n13034\,
            carryout => \quad_counter0.n13035\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i11_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36626\,
            in2 => \N__37419\,
            in3 => \N__36612\,
            lcout => encoder0_position_11,
            ltout => OPEN,
            carryin => \quad_counter0.n13035\,
            carryout => \quad_counter0.n13036\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i12_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37388\,
            in2 => \N__36601\,
            in3 => \N__36573\,
            lcout => encoder0_position_12,
            ltout => OPEN,
            carryin => \quad_counter0.n13036\,
            carryout => \quad_counter0.n13037\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i13_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36565\,
            in2 => \N__37420\,
            in3 => \N__36546\,
            lcout => encoder0_position_13,
            ltout => OPEN,
            carryin => \quad_counter0.n13037\,
            carryout => \quad_counter0.n13038\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i14_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37392\,
            in2 => \N__36720\,
            in3 => \N__36543\,
            lcout => encoder0_position_14,
            ltout => OPEN,
            carryin => \quad_counter0.n13038\,
            carryout => \quad_counter0.n13039\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i15_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42437\,
            in2 => \N__37421\,
            in3 => \N__36540\,
            lcout => encoder0_position_15,
            ltout => OPEN,
            carryin => \quad_counter0.n13039\,
            carryout => \quad_counter0.n13040\,
            clk => \N__55784\,
            ce => \N__39113\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i16_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41908\,
            in2 => \N__37422\,
            in3 => \N__36693\,
            lcout => encoder0_position_16,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \quad_counter0.n13041\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i17_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37399\,
            in2 => \N__42289\,
            in3 => \N__36690\,
            lcout => encoder0_position_17,
            ltout => OPEN,
            carryin => \quad_counter0.n13041\,
            carryout => \quad_counter0.n13042\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i18_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42373\,
            in2 => \N__37423\,
            in3 => \N__36687\,
            lcout => encoder0_position_18,
            ltout => OPEN,
            carryin => \quad_counter0.n13042\,
            carryout => \quad_counter0.n13043\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i19_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37403\,
            in2 => \N__45809\,
            in3 => \N__36684\,
            lcout => encoder0_position_19,
            ltout => OPEN,
            carryin => \quad_counter0.n13043\,
            carryout => \quad_counter0.n13044\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i20_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44605\,
            in2 => \N__37424\,
            in3 => \N__36681\,
            lcout => encoder0_position_20,
            ltout => OPEN,
            carryin => \quad_counter0.n13044\,
            carryout => \quad_counter0.n13045\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i21_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37407\,
            in2 => \N__46331\,
            in3 => \N__36678\,
            lcout => encoder0_position_21,
            ltout => OPEN,
            carryin => \quad_counter0.n13045\,
            carryout => \quad_counter0.n13046\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i22_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44798\,
            in2 => \N__37425\,
            in3 => \N__36675\,
            lcout => encoder0_position_22,
            ltout => OPEN,
            carryin => \quad_counter0.n13046\,
            carryout => \quad_counter0.n13047\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i23_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37411\,
            in2 => \N__41992\,
            in3 => \N__36672\,
            lcout => encoder0_position_23,
            ltout => OPEN,
            carryin => \quad_counter0.n13047\,
            carryout => \quad_counter0.n13048\,
            clk => \N__55786\,
            ce => \N__39111\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i24_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37353\,
            in2 => \N__44728\,
            in3 => \N__36669\,
            lcout => encoder0_position_24,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \quad_counter0.n13049\,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i25_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40355\,
            in2 => \N__37412\,
            in3 => \N__36753\,
            lcout => encoder0_position_25,
            ltout => OPEN,
            carryin => \quad_counter0.n13049\,
            carryout => \quad_counter0.n13050\,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i26_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37357\,
            in2 => \N__42724\,
            in3 => \N__36750\,
            lcout => encoder0_position_26,
            ltout => OPEN,
            carryin => \quad_counter0.n13050\,
            carryout => \quad_counter0.n13051\,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i27_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42813\,
            in2 => \N__37413\,
            in3 => \N__36747\,
            lcout => encoder0_position_27,
            ltout => OPEN,
            carryin => \quad_counter0.n13051\,
            carryout => \quad_counter0.n13052\,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i28_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37361\,
            in2 => \N__40428\,
            in3 => \N__36744\,
            lcout => encoder0_position_28,
            ltout => OPEN,
            carryin => \quad_counter0.n13052\,
            carryout => \quad_counter0.n13053\,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i29_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40735\,
            in2 => \N__37414\,
            in3 => \N__36741\,
            lcout => encoder0_position_29,
            ltout => OPEN,
            carryin => \quad_counter0.n13053\,
            carryout => \quad_counter0.n13054\,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i30_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37365\,
            in2 => \N__40665\,
            in3 => \N__36738\,
            lcout => encoder0_position_30,
            ltout => OPEN,
            carryin => \quad_counter0.n13054\,
            carryout => \quad_counter0.n13055\,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_656__i31_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37366\,
            in1 => \N__46061\,
            in2 => \_gnd_net_\,
            in3 => \N__36735\,
            lcout => encoder0_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55787\,
            ce => \N__39112\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36732\,
            lcout => n8_adj_575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44606\,
            lcout => n13_adj_634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38628\,
            in1 => \N__36719\,
            in2 => \_gnd_net_\,
            in3 => \N__46053\,
            lcout => n305,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i1_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__42932\,
            in1 => \N__55331\,
            in2 => \_gnd_net_\,
            in3 => \N__37530\,
            lcout => pwm_setpoint_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36969\,
            lcout => n21_adj_556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i0_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55330\,
            in1 => \N__37440\,
            in2 => \_gnd_net_\,
            in3 => \N__42968\,
            lcout => pwm_setpoint_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36957\,
            lcout => n20_adj_557,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.debounce_cnt_50_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__39162\,
            in1 => \N__36992\,
            in2 => \N__39080\,
            in3 => \N__38927\,
            lcout => \quad_counter0.debounce_cnt\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36945\,
            lcout => n3_adj_580,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_new_i1_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36993\,
            lcout => a_new_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9962_3_lut_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40056\,
            in2 => \N__36932\,
            in3 => \N__36905\,
            lcout => OPEN,
            ltout => \n11930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_34_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__36875\,
            in1 => \N__36835\,
            in2 => \N__36801\,
            in3 => \N__36794\,
            lcout => n13819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12559_4_lut_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__36991\,
            in1 => \N__39160\,
            in2 => \N__39081\,
            in3 => \N__38926\,
            lcout => \quad_counter0.a_prev_N_543\,
            ltout => \quad_counter0.a_prev_N_543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_52_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__39161\,
            in1 => \N__39045\,
            in2 => \N__37428\,
            in3 => \N__39135\,
            lcout => b_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_I_0_63_2_lut_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39070\,
            in2 => \_gnd_net_\,
            in3 => \N__39042\,
            lcout => \quad_counter0.direction_N_536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2059_3_lut_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37265\,
            in2 => \N__37239\,
            in3 => \N__37215\,
            lcout => n3123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i8_1_lut_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43392\,
            lcout => n18_adj_598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_new_i0_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37011\,
            lcout => \quad_counter0.a_new_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i3_1_lut_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42896\,
            lcout => n23_adj_603,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i2_1_lut_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42933\,
            lcout => n24_adj_604,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36981\,
            lcout => n4_adj_579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n6_adj_577,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i1_1_lut_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42969\,
            lcout => n25_adj_605,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i13_1_lut_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44094\,
            lcout => n13_adj_593,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i20_1_lut_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43907\,
            lcout => n6_adj_586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i9_1_lut_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46908\,
            lcout => n17_adj_597,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i4_1_lut_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43518\,
            lcout => n22_adj_602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i16_1_lut_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43634\,
            lcout => n10_adj_590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i12_1_lut_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44007\,
            lcout => n14_adj_594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_2_lut_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37449\,
            in2 => \_gnd_net_\,
            in3 => \N__37431\,
            lcout => \pwm_setpoint_23_N_171_0\,
            ltout => OPEN,
            carryin => \bfn_9_30_0_\,
            carryout => n12412,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_3_lut_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37539\,
            in2 => \_gnd_net_\,
            in3 => \N__37521\,
            lcout => \pwm_setpoint_23_N_171_1\,
            ltout => OPEN,
            carryin => n12412,
            carryout => n12413,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_4_lut_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37518\,
            in2 => \_gnd_net_\,
            in3 => \N__37509\,
            lcout => \pwm_setpoint_23_N_171_2\,
            ltout => OPEN,
            carryin => n12413,
            carryout => n12414,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_5_lut_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37506\,
            in2 => \_gnd_net_\,
            in3 => \N__37500\,
            lcout => \pwm_setpoint_23_N_171_3\,
            ltout => OPEN,
            carryin => n12414,
            carryout => n12415,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_6_lut_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39303\,
            in2 => \_gnd_net_\,
            in3 => \N__37497\,
            lcout => \pwm_setpoint_23_N_171_4\,
            ltout => OPEN,
            carryin => n12415,
            carryout => n12416,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_7_lut_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39321\,
            in2 => \_gnd_net_\,
            in3 => \N__37494\,
            lcout => \pwm_setpoint_23_N_171_5\,
            ltout => OPEN,
            carryin => n12416,
            carryout => n12417,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_8_lut_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39468\,
            in2 => \_gnd_net_\,
            in3 => \N__37491\,
            lcout => \pwm_setpoint_23_N_171_6\,
            ltout => OPEN,
            carryin => n12417,
            carryout => n12418,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_9_lut_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37488\,
            in2 => \_gnd_net_\,
            in3 => \N__37479\,
            lcout => \pwm_setpoint_23_N_171_7\,
            ltout => OPEN,
            carryin => n12418,
            carryout => n12419,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_10_lut_LC_9_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37476\,
            in2 => \_gnd_net_\,
            in3 => \N__37467\,
            lcout => \pwm_setpoint_23_N_171_8\,
            ltout => OPEN,
            carryin => \bfn_9_31_0_\,
            carryout => n12420,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_11_lut_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39315\,
            in2 => \_gnd_net_\,
            in3 => \N__37464\,
            lcout => \pwm_setpoint_23_N_171_9\,
            ltout => OPEN,
            carryin => n12420,
            carryout => n12421,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_12_lut_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39309\,
            in2 => \_gnd_net_\,
            in3 => \N__37593\,
            lcout => \pwm_setpoint_23_N_171_10\,
            ltout => OPEN,
            carryin => n12421,
            carryout => n12422,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_13_lut_LC_9_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37590\,
            in2 => \_gnd_net_\,
            in3 => \N__37581\,
            lcout => \pwm_setpoint_23_N_171_11\,
            ltout => OPEN,
            carryin => n12422,
            carryout => n12423,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_14_lut_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37578\,
            in2 => \_gnd_net_\,
            in3 => \N__37569\,
            lcout => \pwm_setpoint_23_N_171_12\,
            ltout => OPEN,
            carryin => n12423,
            carryout => n12424,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_15_lut_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39261\,
            in2 => \_gnd_net_\,
            in3 => \N__37566\,
            lcout => \pwm_setpoint_23_N_171_13\,
            ltout => OPEN,
            carryin => n12424,
            carryout => n12425,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_16_lut_LC_9_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39582\,
            in2 => \_gnd_net_\,
            in3 => \N__37563\,
            lcout => \pwm_setpoint_23_N_171_14\,
            ltout => OPEN,
            carryin => n12425,
            carryout => n12426,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_17_lut_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37560\,
            in2 => \_gnd_net_\,
            in3 => \N__37551\,
            lcout => \pwm_setpoint_23_N_171_15\,
            ltout => OPEN,
            carryin => n12426,
            carryout => n12427,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_18_lut_LC_9_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39564\,
            in2 => \_gnd_net_\,
            in3 => \N__37548\,
            lcout => \pwm_setpoint_23_N_171_16\,
            ltout => OPEN,
            carryin => \bfn_9_32_0_\,
            carryout => n12428,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_19_lut_LC_9_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41100\,
            in2 => \_gnd_net_\,
            in3 => \N__37545\,
            lcout => \pwm_setpoint_23_N_171_17\,
            ltout => OPEN,
            carryin => n12428,
            carryout => n12429,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_20_lut_LC_9_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39438\,
            in2 => \_gnd_net_\,
            in3 => \N__37542\,
            lcout => \pwm_setpoint_23_N_171_18\,
            ltout => OPEN,
            carryin => n12429,
            carryout => n12430,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_21_lut_LC_9_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37617\,
            in2 => \_gnd_net_\,
            in3 => \N__37608\,
            lcout => \pwm_setpoint_23_N_171_19\,
            ltout => OPEN,
            carryin => n12430,
            carryout => n12431,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_22_lut_LC_9_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41091\,
            in2 => \_gnd_net_\,
            in3 => \N__37605\,
            lcout => \pwm_setpoint_23_N_171_20\,
            ltout => OPEN,
            carryin => n12431,
            carryout => n12432,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_23_lut_LC_9_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44112\,
            in3 => \N__37602\,
            lcout => \pwm_setpoint_23_N_171_21\,
            ltout => OPEN,
            carryin => n12432,
            carryout => n12433,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_24_lut_LC_9_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39570\,
            in2 => \_gnd_net_\,
            in3 => \N__37599\,
            lcout => \pwm_setpoint_23_N_171_22\,
            ltout => OPEN,
            carryin => n12433,
            carryout => n12434,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i23_LC_9_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44339\,
            in2 => \_gnd_net_\,
            in3 => \N__37596\,
            lcout => pwm_setpoint_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55812\,
            ce => 'H',
            sr => \N__44340\
        );

    \i1_3_lut_adj_85_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39607\,
            in2 => \N__37640\,
            in3 => \N__37786\,
            lcout => n14408,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1246_3_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41226\,
            in2 => \N__41838\,
            in3 => \N__39839\,
            lcout => n1926,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1182_3_lut_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44250\,
            in2 => \N__41803\,
            in3 => \N__45690\,
            lcout => n1830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1253_3_lut_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41448\,
            in1 => \N__42423\,
            in2 => \_gnd_net_\,
            in3 => \N__39840\,
            lcout => n1933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38469\,
            in1 => \N__46181\,
            in2 => \_gnd_net_\,
            in3 => \N__37848\,
            lcout => n310,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1247_3_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41261\,
            in2 => \N__41241\,
            in3 => \N__39838\,
            lcout => n1927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1243_3_lut_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41626\,
            in2 => \N__39874\,
            in3 => \N__41604\,
            lcout => n1923,
            ltout => \n1923_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_86_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37741\,
            in2 => \N__37725\,
            in3 => \N__37714\,
            lcout => n14410,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1244_3_lut_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41660\,
            in2 => \N__39873\,
            in3 => \N__41640\,
            lcout => n1924,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1241_3_lut_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__39852\,
            in1 => \_gnd_net_\,
            in2 => \N__41523\,
            in3 => \N__41553\,
            lcout => n1921,
            ltout => \n1921_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_87_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38048\,
            in1 => \N__37698\,
            in2 => \N__37692\,
            in3 => \N__37689\,
            lcout => n14416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1315_3_lut_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37683\,
            in2 => \N__39617\,
            in3 => \N__38173\,
            lcout => n2027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1245_3_lut_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41676\,
            in2 => \N__41694\,
            in3 => \N__39845\,
            lcout => n1925,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1242_3_lut_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41591\,
            in2 => \N__41571\,
            in3 => \N__39867\,
            lcout => n1922,
            ltout => \n1922_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1309_3_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38037\,
            in2 => \N__38031\,
            in3 => \N__38197\,
            lcout => n2021,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_89_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__39730\,
            in1 => \N__37854\,
            in2 => \N__39630\,
            in3 => \N__37998\,
            lcout => OPEN,
            ltout => \n14420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12944_4_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39914\,
            in1 => \N__39703\,
            in2 => \N__37992\,
            in3 => \N__37922\,
            lcout => n1950,
            ltout => \n1950_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1318_3_lut_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39950\,
            in2 => \N__37989\,
            in3 => \N__37986\,
            lcout => n2030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12941_1_lut_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38198\,
            lcout => n15666,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1237_3_lut_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44523\,
            in2 => \N__41871\,
            in3 => \N__39868\,
            lcout => n1917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1308_3_lut_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37911\,
            in2 => \N__37905\,
            in3 => \N__38196\,
            lcout => n2020,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9998_4_lut_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__38360\,
            in1 => \N__39946\,
            in2 => \N__38457\,
            in3 => \N__38234\,
            lcout => n11966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1252_3_lut_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41412\,
            in2 => \N__39884\,
            in3 => \N__41432\,
            lcout => n1932,
            ltout => \n1932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1319_3_lut_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__38179\,
            in1 => \_gnd_net_\,
            in2 => \N__38439\,
            in3 => \N__38436\,
            lcout => n2031,
            ltout => \n2031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9996_4_lut_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__38403\,
            in1 => \N__38099\,
            in2 => \N__38370\,
            in3 => \N__38302\,
            lcout => n11964,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1321_3_lut_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__38361\,
            in1 => \N__38334\,
            in2 => \N__38205\,
            in3 => \_gnd_net_\,
            lcout => n2033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1316_3_lut_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38289\,
            in2 => \N__39663\,
            in3 => \N__38178\,
            lcout => n2028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1320_3_lut_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38250\,
            in2 => \N__38238\,
            in3 => \N__38174\,
            lcout => n2032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38088\,
            in3 => \N__38067\,
            lcout => n33,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => n12968,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38064\,
            in3 => \N__38055\,
            lcout => n32,
            ltout => OPEN,
            carryin => n12968,
            carryout => n12969,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38592\,
            in3 => \N__38583\,
            lcout => n31,
            ltout => OPEN,
            carryin => n12969,
            carryout => n12970,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40167\,
            in3 => \N__38580\,
            lcout => n30,
            ltout => OPEN,
            carryin => n12970,
            carryout => n12971,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38577\,
            in3 => \N__38556\,
            lcout => n29,
            ltout => OPEN,
            carryin => n12971,
            carryout => n12972,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38553\,
            in3 => \N__38544\,
            lcout => n28,
            ltout => OPEN,
            carryin => n12972,
            carryout => n12973,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38541\,
            in3 => \N__38532\,
            lcout => n27,
            ltout => OPEN,
            carryin => n12973,
            carryout => n12974,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38529\,
            in3 => \N__38520\,
            lcout => n26,
            ltout => OPEN,
            carryin => n12974,
            carryout => n12975,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38517\,
            in3 => \N__38484\,
            lcout => n25_adj_551,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => n12976,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38481\,
            in3 => \N__38460\,
            lcout => n24,
            ltout => OPEN,
            carryin => n12976,
            carryout => n12977,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39978\,
            in3 => \N__38739\,
            lcout => n23,
            ltout => OPEN,
            carryin => n12977,
            carryout => n12978,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38736\,
            in2 => \_gnd_net_\,
            in3 => \N__38718\,
            lcout => n22,
            ltout => OPEN,
            carryin => n12978,
            carryout => n12979,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38715\,
            in3 => \N__38682\,
            lcout => n21,
            ltout => OPEN,
            carryin => n12979,
            carryout => n12980,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38679\,
            in3 => \N__38646\,
            lcout => n20,
            ltout => OPEN,
            carryin => n12980,
            carryout => n12981,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38643\,
            in3 => \N__38616\,
            lcout => n19,
            ltout => OPEN,
            carryin => n12981,
            carryout => n12982,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41946\,
            in3 => \N__38613\,
            lcout => n18,
            ltout => OPEN,
            carryin => n12982,
            carryout => n12983,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38610\,
            in3 => \N__38598\,
            lcout => n17,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => n12984,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41709\,
            in3 => \N__38595\,
            lcout => n16,
            ltout => OPEN,
            carryin => n12984,
            carryout => n12985,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38805\,
            in3 => \N__38793\,
            lcout => n15,
            ltout => OPEN,
            carryin => n12985,
            carryout => n12986,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45789\,
            in3 => \N__38790\,
            lcout => n14,
            ltout => OPEN,
            carryin => n12986,
            carryout => n12987,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38787\,
            in3 => \N__38775\,
            lcout => n13,
            ltout => OPEN,
            carryin => n12987,
            carryout => n12988,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46305\,
            in3 => \N__38772\,
            lcout => n12,
            ltout => OPEN,
            carryin => n12988,
            carryout => n12989,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44784\,
            in3 => \N__38769\,
            lcout => n11,
            ltout => OPEN,
            carryin => n12989,
            carryout => n12990,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41961\,
            in3 => \N__38766\,
            lcout => n10,
            ltout => OPEN,
            carryin => n12990,
            carryout => n12991,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44706\,
            in3 => \N__38763\,
            lcout => n9,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => n12992,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38823\,
            in3 => \N__38760\,
            lcout => n8,
            ltout => OPEN,
            carryin => n12992,
            carryout => n12993,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38814\,
            in3 => \N__38757\,
            lcout => n7,
            ltout => OPEN,
            carryin => n12993,
            carryout => n12994,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38832\,
            in3 => \N__38856\,
            lcout => n6,
            ltout => OPEN,
            carryin => n12994,
            carryout => n12995,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38841\,
            in3 => \N__38853\,
            lcout => n5,
            ltout => OPEN,
            carryin => n12995,
            carryout => n12996,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39018\,
            in3 => \N__38850\,
            lcout => n4,
            ltout => OPEN,
            carryin => n12996,
            carryout => n12997,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39201\,
            in3 => \N__38847\,
            lcout => n3,
            ltout => OPEN,
            carryin => n12997,
            carryout => n12998,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42102\,
            in3 => \N__38844\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40416\,
            lcout => n5_adj_626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42814\,
            in3 => \_gnd_net_\,
            lcout => n6_adj_627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_166_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__46031\,
            in1 => \_gnd_net_\,
            in2 => \N__40689\,
            in3 => \N__40464\,
            lcout => n14574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40351\,
            lcout => n8_adj_629,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42709\,
            lcout => n7_adj_628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46029\,
            in2 => \N__42815\,
            in3 => \N__42865\,
            lcout => n292,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40728\,
            lcout => n4_adj_625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46030\,
            in2 => \N__40663\,
            in3 => \N__40684\,
            lcout => n403,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i4_4_lut_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__45180\,
            in1 => \N__39009\,
            in2 => \N__45201\,
            in3 => \N__39003\,
            lcout => n4_adj_655,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i6_3_lut_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38997\,
            in1 => \N__46060\,
            in2 => \_gnd_net_\,
            in3 => \N__38988\,
            lcout => n314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_new_i1_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38928\,
            lcout => \quad_counter0.b_new_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n25_adj_552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38880\,
            lcout => n10_adj_573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38868\,
            lcout => n12_adj_571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40653\,
            lcout => n3_adj_624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39189\,
            lcout => n23_adj_554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12508_3_lut_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43781\,
            in1 => \N__43762\,
            in2 => \_gnd_net_\,
            in3 => \N__39177\,
            lcout => n15233,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_prev_51_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__39144\,
            in1 => \N__39134\,
            in2 => \N__39171\,
            in3 => \N__39076\,
            lcout => \quad_counter0.a_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_I_0_65_2_lut_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39159\,
            in2 => \_gnd_net_\,
            in3 => \N__39043\,
            lcout => OPEN,
            ltout => \quad_counter0.direction_N_540_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001000"
        )
    port map (
            in0 => \N__39143\,
            in1 => \N__39133\,
            in2 => \N__39120\,
            in3 => \N__39074\,
            lcout => \direction_N_537\,
            ltout => \direction_N_537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.direction_57_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110010101100"
        )
    port map (
            in0 => \N__39075\,
            in1 => \N__39024\,
            in2 => \N__39048\,
            in3 => \N__39044\,
            lcout => n1302,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i29_2_lut_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__39212\,
            in1 => \N__46637\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n29_adj_672,
            ltout => \n29_adj_672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12509_3_lut_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39213\,
            in2 => \N__39291\,
            in3 => \N__39288\,
            lcout => n15234,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12457_3_lut_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39399\,
            in1 => \N__39382\,
            in2 => \_gnd_net_\,
            in3 => \N__39282\,
            lcout => n15182,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n9_adj_574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i33_2_lut_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46593\,
            in2 => \_gnd_net_\,
            in3 => \N__40911\,
            lcout => n33_adj_675,
            ltout => \n33_adj_675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12396_4_lut_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__39350\,
            in1 => \N__39383\,
            in2 => \N__39264\,
            in3 => \N__40782\,
            lcout => n15121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i14_1_lut_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43701\,
            lcout => n12_adj_592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i16_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43599\,
            in1 => \N__55307\,
            in2 => \_gnd_net_\,
            in3 => \N__39252\,
            lcout => pwm_setpoint_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i2_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__55306\,
            in1 => \_gnd_net_\,
            in2 => \N__39240\,
            in3 => \N__42897\,
            lcout => pwm_setpoint_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55794\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i14_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__43674\,
            in1 => \_gnd_net_\,
            in2 => \N__39228\,
            in3 => \N__55329\,
            lcout => pwm_setpoint_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55797\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i10_3_lut_3_lut_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__45306\,
            in1 => \N__45284\,
            in2 => \_gnd_net_\,
            in3 => \N__46713\,
            lcout => n10_adj_659,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12552_4_lut_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__39366\,
            in1 => \N__43821\,
            in2 => \N__39330\,
            in3 => \N__39360\,
            lcout => n15277,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12500_4_lut_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__39384\,
            in1 => \N__39354\,
            in2 => \N__43767\,
            in3 => \N__47379\,
            lcout => n15225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i30_3_lut_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43941\,
            in1 => \N__40929\,
            in2 => \_gnd_net_\,
            in3 => \N__43819\,
            lcout => OPEN,
            ltout => \n30_adj_673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12542_4_lut_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__43820\,
            in1 => \N__40881\,
            in2 => \N__39339\,
            in3 => \N__39336\,
            lcout => n15267,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i6_1_lut_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43448\,
            lcout => n20_adj_600,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i10_1_lut_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43352\,
            lcout => n16_adj_596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i11_1_lut_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43325\,
            lcout => n15_adj_595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i5_1_lut_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43478\,
            lcout => n21_adj_601,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i5_LC_10_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55323\,
            in1 => \N__39297\,
            in2 => \_gnd_net_\,
            in3 => \N__43449\,
            lcout => pwm_setpoint_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i7_1_lut_LC_10_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43421\,
            lcout => n19_adj_599,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i6_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55324\,
            in1 => \_gnd_net_\,
            in2 => \N__43425\,
            in3 => \N__39462\,
            lcout => pwm_setpoint_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i10_LC_10_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43326\,
            in1 => \N__55325\,
            in2 => \_gnd_net_\,
            in3 => \N__39456\,
            lcout => pwm_setpoint_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55801\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i9_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55326\,
            in1 => \N__39450\,
            in2 => \_gnd_net_\,
            in3 => \N__43353\,
            lcout => pwm_setpoint_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i4_LC_10_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43485\,
            in1 => \N__55328\,
            in2 => \_gnd_net_\,
            in3 => \N__39444\,
            lcout => pwm_setpoint_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i19_1_lut_LC_10_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43553\,
            lcout => n7_adj_587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i15_LC_10_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43635\,
            in1 => \N__55327\,
            in2 => \_gnd_net_\,
            in3 => \N__39432\,
            lcout => pwm_setpoint_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i1_LC_10_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47581\,
            in1 => \N__39425\,
            in2 => \_gnd_net_\,
            in3 => \N__39539\,
            lcout => h2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55806\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i31_2_lut_LC_10_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39395\,
            in2 => \_gnd_net_\,
            in3 => \N__46454\,
            lcout => n31_adj_674,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i15_1_lut_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43673\,
            lcout => n11_adj_591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i18_LC_10_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55332\,
            in1 => \N__43554\,
            in2 => \_gnd_net_\,
            in3 => \N__39576\,
            lcout => pwm_setpoint_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12212_4_lut_LC_10_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111100000"
        )
    port map (
            in0 => \N__41181\,
            in1 => \N__41145\,
            in2 => \N__41205\,
            in3 => \N__41163\,
            lcout => n14937,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i23_1_lut_LC_10_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43847\,
            lcout => n3_adj_583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i17_1_lut_LC_10_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43598\,
            lcout => n9_adj_589,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i2_LC_10_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__39558\,
            in1 => \N__39526\,
            in2 => \_gnd_net_\,
            in3 => \N__47621\,
            lcout => h1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12211_4_lut_LC_10_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010110000"
        )
    port map (
            in0 => \N__41180\,
            in1 => \N__41144\,
            in2 => \N__41204\,
            in3 => \N__41162\,
            lcout => OPEN,
            ltout => \n14936_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12213_3_lut_LC_10_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__39498\,
            in1 => \_gnd_net_\,
            in2 => \N__39492\,
            in3 => \N__41124\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i22_LC_10_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43848\,
            in1 => \N__55333\,
            in2 => \_gnd_net_\,
            in3 => \N__39474\,
            lcout => pwm_setpoint_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1181_3_lut_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44238\,
            in2 => \N__41804\,
            in3 => \N__45535\,
            lcout => n1829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12513_3_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49790\,
            in2 => \N__44466\,
            in3 => \N__41796\,
            lcout => n1826,
            ltout => \n1826_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_81_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41827\,
            in1 => \N__41257\,
            in2 => \N__39621\,
            in3 => \N__41656\,
            lcout => n14526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1248_3_lut_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41291\,
            in2 => \N__41274\,
            in3 => \N__39841\,
            lcout => n1928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_82_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41587\,
            in2 => \N__41627\,
            in3 => \N__39591\,
            lcout => OPEN,
            ltout => \n14530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_83_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__41320\,
            in1 => \N__41290\,
            in2 => \N__39585\,
            in3 => \N__39762\,
            lcout => n14532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1249_3_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41321\,
            in2 => \N__39872\,
            in3 => \N__41301\,
            lcout => n1929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_79_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45495\,
            in3 => \N__45537\,
            lcout => n14520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1180_3_lut_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45493\,
            in2 => \N__44226\,
            in3 => \N__41760\,
            lcout => n1828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1175_3_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44424\,
            in2 => \N__41790\,
            in3 => \N__50313\,
            lcout => n1823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1176_3_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50286\,
            in2 => \N__44439\,
            in3 => \N__41767\,
            lcout => n1824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12443_3_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50343\,
            in2 => \N__41789\,
            in3 => \N__44451\,
            lcout => n1825,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1171_3_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44562\,
            in2 => \N__44583\,
            in3 => \N__41768\,
            lcout => n1819,
            ltout => \n1819_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12922_4_lut_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40176\,
            in1 => \N__44519\,
            in2 => \N__39753\,
            in3 => \N__39750\,
            lcout => n1851,
            ltout => \n1851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1240_3_lut_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__41856\,
            in1 => \N__41508\,
            in2 => \N__39744\,
            in3 => \_gnd_net_\,
            lcout => n1920,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1239_3_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41495\,
            in1 => \_gnd_net_\,
            in2 => \N__39882\,
            in3 => \N__41481\,
            lcout => n1919,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1250_3_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41337\,
            in1 => \_gnd_net_\,
            in2 => \N__41363\,
            in3 => \N__39860\,
            lcout => n1930,
            ltout => \n1930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_88_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39666\,
            in3 => \N__39652\,
            lcout => n14540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1251_3_lut_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41376\,
            in2 => \N__41396\,
            in3 => \N__39859\,
            lcout => n1931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1238_3_lut_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41471\,
            in2 => \N__39881\,
            in3 => \N__41457\,
            lcout => n1918,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_80_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__44393\,
            in1 => \N__45609\,
            in2 => \N__39903\,
            in3 => \N__50223\,
            lcout => OPEN,
            ltout => \n14176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12901_4_lut_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44371\,
            in1 => \N__44578\,
            in2 => \N__39894\,
            in3 => \N__47942\,
            lcout => n1752,
            ltout => \n1752_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1183_3_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44265\,
            in2 => \N__39891\,
            in3 => \N__45597\,
            lcout => n1831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12919_1_lut_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39883\,
            lcout => n15644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1184_3_lut_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45669\,
            in2 => \N__44283\,
            in3 => \N__41770\,
            lcout => n1832,
            ltout => \n1832_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10000_4_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__41353\,
            in1 => \N__42406\,
            in2 => \N__39765\,
            in3 => \N__41431\,
            lcout => n11968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1185_3_lut_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44301\,
            in1 => \N__45634\,
            in2 => \_gnd_net_\,
            in3 => \N__41769\,
            lcout => n1833,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1172_3_lut_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44373\,
            in1 => \_gnd_net_\,
            in2 => \N__41792\,
            in3 => \N__44355\,
            lcout => n1820,
            ltout => \n1820_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_84_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41539\,
            in2 => \N__40179\,
            in3 => \N__41854\,
            lcout => n14538,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1174_3_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44412\,
            in2 => \N__41791\,
            in3 => \N__50253\,
            lcout => n1822,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42251\,
            lcout => n30_adj_651,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i8_3_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40158\,
            in1 => \N__46192\,
            in2 => \_gnd_net_\,
            in3 => \N__40152\,
            lcout => n312,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i3_3_lut_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46193\,
            in1 => \N__40086\,
            in2 => \_gnd_net_\,
            in3 => \N__40080\,
            lcout => n317,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40006\,
            lcout => n23_adj_644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39969\,
            lcout => n24_adj_553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_2_lut_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40329\,
            in3 => \N__39957\,
            lcout => n901,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => n12487,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_3_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52980\,
            in2 => \N__42687\,
            in3 => \N__40230\,
            lcout => n900,
            ltout => OPEN,
            carryin => n12487,
            carryout => n12488,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_4_lut_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42786\,
            in3 => \N__40227\,
            lcout => n899,
            ltout => OPEN,
            carryin => n12488,
            carryout => n12489,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_5_lut_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52981\,
            in2 => \N__40449\,
            in3 => \N__40224\,
            lcout => n898,
            ltout => OPEN,
            carryin => n12489,
            carryout => n12490,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_6_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40497\,
            in3 => \N__40221\,
            lcout => n897,
            ltout => OPEN,
            carryin => n12490,
            carryout => n12491,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_7_lut_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40629\,
            in3 => \N__40218\,
            lcout => n896,
            ltout => OPEN,
            carryin => n12491,
            carryout => n12492,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_8_lut_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__52982\,
            in1 => \N__40275\,
            in2 => \N__40296\,
            in3 => \N__40215\,
            lcout => n927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i573_3_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40327\,
            in2 => \N__40212\,
            in3 => \N__40262\,
            lcout => n933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i568_3_lut_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40628\,
            in2 => \N__40274\,
            in3 => \N__40200\,
            lcout => n928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i572_3_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42682\,
            in2 => \N__40194\,
            in3 => \N__40261\,
            lcout => n932,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i571_3_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42782\,
            in2 => \N__40273\,
            in3 => \N__40185\,
            lcout => n931,
            ltout => \n931_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9972_4_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__44756\,
            in1 => \N__42745\,
            in2 => \N__40383\,
            in3 => \N__44680\,
            lcout => n11940,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i24_3_lut_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46151\,
            in2 => \N__40380\,
            in3 => \N__41994\,
            lcout => n296,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i569_3_lut_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40493\,
            in2 => \N__40371\,
            in3 => \N__40263\,
            lcout => n929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i26_3_lut_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46150\,
            in2 => \N__40362\,
            in3 => \N__40335\,
            lcout => n294,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10044_4_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__42778\,
            in1 => \N__40328\,
            in2 => \N__42683\,
            in3 => \N__40441\,
            lcout => n12012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i500_4_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__43254\,
            in1 => \N__42326\,
            in2 => \N__40305\,
            in3 => \N__46154\,
            lcout => n828,
            ltout => \n828_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10130_4_lut_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__40489\,
            in1 => \N__40618\,
            in2 => \N__40284\,
            in3 => \N__40281\,
            lcout => n861,
            ltout => \n861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i570_3_lut_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40442\,
            in1 => \_gnd_net_\,
            in2 => \N__40242\,
            in3 => \N__40239\,
            lcout => n930,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10980_3_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40706\,
            in2 => \N__42849\,
            in3 => \N__43299\,
            lcout => OPEN,
            ltout => \n13644_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10981_3_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46153\,
            in2 => \N__40500\,
            in3 => \N__40740\,
            lcout => n830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10986_3_lut_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40473\,
            in1 => \_gnd_net_\,
            in2 => \N__42848\,
            in3 => \N__42630\,
            lcout => n13650,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i27_3_lut_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46152\,
            in2 => \N__42729\,
            in3 => \N__40472\,
            lcout => n293,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_64_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__40393\,
            in1 => \N__42866\,
            in2 => \N__40707\,
            in3 => \N__42641\,
            lcout => n5_adj_676,
            ltout => \n5_adj_676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_65_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40680\,
            in2 => \N__40458\,
            in3 => \N__42316\,
            lcout => n13641,
            ltout => \n13641_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10982_3_lut_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40397\,
            in1 => \_gnd_net_\,
            in2 => \N__40455\,
            in3 => \N__42588\,
            lcout => OPEN,
            ltout => \n13646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10983_3_lut_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46102\,
            in1 => \_gnd_net_\,
            in2 => \N__40452\,
            in3 => \N__40427\,
            lcout => n831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i29_3_lut_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40426\,
            in2 => \N__40398\,
            in3 => \N__46098\,
            lcout => n174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40736\,
            in2 => \N__46165\,
            in3 => \N__40705\,
            lcout => n404,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10978_3_lut_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42847\,
            in2 => \N__40688\,
            in3 => \N__43278\,
            lcout => OPEN,
            ltout => \n13642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10979_3_lut_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__46103\,
            in1 => \N__40664\,
            in2 => \N__40632\,
            in3 => \_gnd_net_\,
            lcout => n829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i2_3_lut_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46180\,
            in1 => \N__40602\,
            in2 => \_gnd_net_\,
            in3 => \N__40590\,
            lcout => n318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40524\,
            lcout => n11_adj_572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_50_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__49019\,
            in1 => \N__48940\,
            in2 => \N__49068\,
            in3 => \N__46866\,
            lcout => OPEN,
            ltout => \n10_adj_606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_52_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__48977\,
            in1 => \N__54806\,
            in2 => \N__40512\,
            in3 => \N__48896\,
            lcout => OPEN,
            ltout => \n15_adj_565_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_55_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49547\,
            in1 => \N__49380\,
            in2 => \N__40509\,
            in3 => \N__40506\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_51_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49435\,
            in2 => \_gnd_net_\,
            in3 => \N__54848\,
            lcout => n16_adj_564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40833\,
            lcout => n15_adj_568,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i3_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40821\,
            in1 => \N__43514\,
            in2 => \_gnd_net_\,
            in3 => \N__55263\,
            lcout => pwm_setpoint_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55795\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40809\,
            lcout => n14_adj_569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i13_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43697\,
            in1 => \N__55262\,
            in2 => \_gnd_net_\,
            in3 => \N__40797\,
            lcout => pwm_setpoint_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55795\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i15_2_lut_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46748\,
            in2 => \_gnd_net_\,
            in3 => \N__40896\,
            lcout => n15_adj_663,
            ltout => \n15_adj_663_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12400_4_lut_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__47445\,
            in1 => \N__47421\,
            in2 => \N__40785\,
            in3 => \N__43763\,
            lcout => n15125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40776\,
            lcout => n7_adj_576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40764\,
            lcout => n5_adj_578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40752\,
            lcout => n2_adj_581,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i12_3_lut_3_lut_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__46591\,
            in1 => \N__40909\,
            in2 => \_gnd_net_\,
            in3 => \N__40894\,
            lcout => n12_adj_661,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i37_2_lut_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46476\,
            lcout => n37,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i7_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43391\,
            in1 => \N__55261\,
            in2 => \_gnd_net_\,
            in3 => \N__40923\,
            lcout => pwm_setpoint_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55798\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12394_2_lut_4_lut_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__46592\,
            in1 => \N__40910\,
            in2 => \N__46752\,
            in3 => \N__40895\,
            lcout => n15119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i6_3_lut_3_lut_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__46841\,
            in1 => \N__46826\,
            in2 => \_gnd_net_\,
            in3 => \N__46797\,
            lcout => n6_adj_656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40875\,
            lcout => n16_adj_563,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i0_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40860\,
            in2 => \_gnd_net_\,
            in3 => \N__40854\,
            lcout => n26_adj_697,
            ltout => OPEN,
            carryin => \bfn_11_29_0_\,
            carryout => n13087,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i1_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40851\,
            in2 => \_gnd_net_\,
            in3 => \N__40845\,
            lcout => n25_adj_696,
            ltout => OPEN,
            carryin => n13087,
            carryout => n13088,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i2_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40842\,
            in2 => \_gnd_net_\,
            in3 => \N__40836\,
            lcout => n24_adj_695,
            ltout => OPEN,
            carryin => n13088,
            carryout => n13089,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i3_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41010\,
            in2 => \_gnd_net_\,
            in3 => \N__41004\,
            lcout => n23_adj_694,
            ltout => OPEN,
            carryin => n13089,
            carryout => n13090,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i4_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41001\,
            in2 => \_gnd_net_\,
            in3 => \N__40995\,
            lcout => n22_adj_693,
            ltout => OPEN,
            carryin => n13090,
            carryout => n13091,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i5_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40992\,
            in2 => \_gnd_net_\,
            in3 => \N__40986\,
            lcout => n21_adj_692,
            ltout => OPEN,
            carryin => n13091,
            carryout => n13092,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i6_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40983\,
            in2 => \_gnd_net_\,
            in3 => \N__40977\,
            lcout => n20_adj_691,
            ltout => OPEN,
            carryin => n13092,
            carryout => n13093,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i7_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40974\,
            in2 => \_gnd_net_\,
            in3 => \N__40968\,
            lcout => n19_adj_690,
            ltout => OPEN,
            carryin => n13093,
            carryout => n13094,
            clk => \N__55802\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i8_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40965\,
            in2 => \_gnd_net_\,
            in3 => \N__40959\,
            lcout => n18_adj_689,
            ltout => OPEN,
            carryin => \bfn_11_30_0_\,
            carryout => n13095,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i9_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40956\,
            in2 => \_gnd_net_\,
            in3 => \N__40950\,
            lcout => n17_adj_688,
            ltout => OPEN,
            carryin => n13095,
            carryout => n13096,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i10_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40947\,
            in2 => \_gnd_net_\,
            in3 => \N__40941\,
            lcout => n16_adj_687,
            ltout => OPEN,
            carryin => n13096,
            carryout => n13097,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i11_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40938\,
            in2 => \_gnd_net_\,
            in3 => \N__40932\,
            lcout => n15_adj_686,
            ltout => OPEN,
            carryin => n13097,
            carryout => n13098,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i12_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41082\,
            in2 => \_gnd_net_\,
            in3 => \N__41076\,
            lcout => n14_adj_685,
            ltout => OPEN,
            carryin => n13098,
            carryout => n13099,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i13_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41073\,
            in2 => \_gnd_net_\,
            in3 => \N__41067\,
            lcout => n13_adj_684,
            ltout => OPEN,
            carryin => n13099,
            carryout => n13100,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i14_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41064\,
            in2 => \_gnd_net_\,
            in3 => \N__41058\,
            lcout => n12_adj_683,
            ltout => OPEN,
            carryin => n13100,
            carryout => n13101,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i15_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41055\,
            in2 => \_gnd_net_\,
            in3 => \N__41049\,
            lcout => n11_adj_682,
            ltout => OPEN,
            carryin => n13101,
            carryout => n13102,
            clk => \N__55807\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i16_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41046\,
            in2 => \_gnd_net_\,
            in3 => \N__41040\,
            lcout => n10_adj_681,
            ltout => OPEN,
            carryin => \bfn_11_31_0_\,
            carryout => n13103,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i17_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41037\,
            in2 => \_gnd_net_\,
            in3 => \N__41031\,
            lcout => n9_adj_680,
            ltout => OPEN,
            carryin => n13103,
            carryout => n13104,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i18_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41028\,
            in2 => \_gnd_net_\,
            in3 => \N__41022\,
            lcout => n8_adj_679,
            ltout => OPEN,
            carryin => n13104,
            carryout => n13105,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i19_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41019\,
            in2 => \_gnd_net_\,
            in3 => \N__41013\,
            lcout => n7_adj_678,
            ltout => OPEN,
            carryin => n13105,
            carryout => n13106,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i20_LC_11_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41214\,
            in2 => \_gnd_net_\,
            in3 => \N__41208\,
            lcout => n6_adj_677,
            ltout => OPEN,
            carryin => n13106,
            carryout => n13107,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i21_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41197\,
            in2 => \_gnd_net_\,
            in3 => \N__41184\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n13107,
            carryout => n13108,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i22_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41179\,
            in2 => \_gnd_net_\,
            in3 => \N__41166\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n13108,
            carryout => n13109,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i23_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41161\,
            in2 => \_gnd_net_\,
            in3 => \N__41148\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n13109,
            carryout => n13110,
            clk => \N__55814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i24_LC_11_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41143\,
            in2 => \_gnd_net_\,
            in3 => \N__41130\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_11_32_0_\,
            carryout => n13111,
            clk => \N__55818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_660__i25_LC_11_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41120\,
            in2 => \_gnd_net_\,
            in3 => \N__41127\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i19_LC_11_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43908\,
            in1 => \N__55334\,
            in2 => \_gnd_net_\,
            in3 => \N__41109\,
            lcout => pwm_setpoint_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i18_1_lut_LC_11_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43974\,
            lcout => n8_adj_588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i21_1_lut_LC_11_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44138\,
            lcout => n5_adj_585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_2_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42419\,
            in2 => \_gnd_net_\,
            in3 => \N__41439\,
            lcout => n1901,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => n12592,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_3_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53101\,
            in2 => \N__41436\,
            in3 => \N__41400\,
            lcout => n1900,
            ltout => OPEN,
            carryin => n12592,
            carryout => n12593,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_4_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41397\,
            in3 => \N__41367\,
            lcout => n1899,
            ltout => OPEN,
            carryin => n12593,
            carryout => n12594,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_5_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53102\,
            in2 => \N__41364\,
            in3 => \N__41325\,
            lcout => n1898,
            ltout => OPEN,
            carryin => n12594,
            carryout => n12595,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_6_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41322\,
            in3 => \N__41295\,
            lcout => n1897,
            ltout => OPEN,
            carryin => n12595,
            carryout => n12596,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_7_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41292\,
            in3 => \N__41265\,
            lcout => n1896,
            ltout => OPEN,
            carryin => n12596,
            carryout => n12597,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_8_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53937\,
            in2 => \N__41262\,
            in3 => \N__41229\,
            lcout => n1895,
            ltout => OPEN,
            carryin => n12597,
            carryout => n12598,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_9_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53103\,
            in2 => \N__41834\,
            in3 => \N__41217\,
            lcout => n1894,
            ltout => OPEN,
            carryin => n12598,
            carryout => n12599,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_10_lut_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53577\,
            in2 => \N__41693\,
            in3 => \N__41664\,
            lcout => n1893,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => n12600,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_11_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53584\,
            in2 => \N__41661\,
            in3 => \N__41631\,
            lcout => n1892,
            ltout => OPEN,
            carryin => n12600,
            carryout => n12601,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_12_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53578\,
            in2 => \N__41628\,
            in3 => \N__41595\,
            lcout => n1891,
            ltout => OPEN,
            carryin => n12601,
            carryout => n12602,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_13_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53585\,
            in2 => \N__41592\,
            in3 => \N__41556\,
            lcout => n1890,
            ltout => OPEN,
            carryin => n12602,
            carryout => n12603,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_14_lut_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53579\,
            in2 => \N__41552\,
            in3 => \N__41511\,
            lcout => n1889,
            ltout => OPEN,
            carryin => n12603,
            carryout => n12604,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_15_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41855\,
            in2 => \N__53936\,
            in3 => \N__41502\,
            lcout => n1888,
            ltout => OPEN,
            carryin => n12604,
            carryout => n12605,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_16_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53583\,
            in2 => \N__41499\,
            in3 => \N__41475\,
            lcout => n1887,
            ltout => OPEN,
            carryin => n12605,
            carryout => n12606,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_17_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53586\,
            in2 => \N__41472\,
            in3 => \N__41451\,
            lcout => n1886,
            ltout => OPEN,
            carryin => n12606,
            carryout => n12607,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_18_lut_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52810\,
            in1 => \N__44518\,
            in2 => \_gnd_net_\,
            in3 => \N__41874\,
            lcout => n1885,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1104_3_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__48027\,
            in1 => \N__48003\,
            in2 => \N__50195\,
            in3 => \_gnd_net_\,
            lcout => n1720,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48112\,
            in2 => \N__48090\,
            in3 => \N__50187\,
            lcout => n1722,
            ltout => \n1722_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__41759\,
            in1 => \_gnd_net_\,
            in2 => \N__41859\,
            in3 => \N__44382\,
            lcout => n1821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1105_3_lut_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48072\,
            in2 => \N__48045\,
            in3 => \N__50188\,
            lcout => n1721,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1179_3_lut_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__44478\,
            in1 => \_gnd_net_\,
            in2 => \N__50109\,
            in3 => \N__41758\,
            lcout => n1827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12897_1_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41785\,
            lcout => n15622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1039_3_lut_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44640\,
            in2 => \N__48420\,
            in3 => \N__50672\,
            lcout => n1623_adj_610,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42290\,
            lcout => n16_adj_637,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2177_2_lut_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46196\,
            in2 => \_gnd_net_\,
            in3 => \N__42330\,
            lcout => n402,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i18_3_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46197\,
            in1 => \N__42303\,
            in2 => \_gnd_net_\,
            in3 => \N__42291\,
            lcout => n302,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i4_3_lut_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42267\,
            in1 => \N__46198\,
            in2 => \_gnd_net_\,
            in3 => \N__42255\,
            lcout => n316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46183\,
            lcout => n2_adj_623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42009\,
            lcout => n18_adj_559,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41993\,
            lcout => n10_adj_631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42443\,
            lcout => n18_adj_639,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46185\,
            in1 => \N__41931\,
            in2 => \_gnd_net_\,
            in3 => \N__41918\,
            lcout => n303,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i16_3_lut_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41886\,
            in1 => \N__46186\,
            in2 => \_gnd_net_\,
            in3 => \N__42444\,
            lcout => n304,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46184\,
            in1 => \N__42390\,
            in2 => \_gnd_net_\,
            in3 => \N__42378\,
            lcout => n301,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_2_lut_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44744\,
            in2 => \_gnd_net_\,
            in3 => \N__42351\,
            lcout => n1001,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => n12493,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_3_lut_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52901\,
            in2 => \N__44687\,
            in3 => \N__42348\,
            lcout => n1000,
            ltout => OPEN,
            carryin => n12493,
            carryout => n12494,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_4_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42752\,
            in3 => \N__42345\,
            lcout => n999,
            ltout => OPEN,
            carryin => n12494,
            carryout => n12495,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_5_lut_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52902\,
            in2 => \N__42473\,
            in3 => \N__42342\,
            lcout => n998,
            ltout => OPEN,
            carryin => n12495,
            carryout => n12496,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_6_lut_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42546\,
            in3 => \N__42339\,
            lcout => n997,
            ltout => OPEN,
            carryin => n12496,
            carryout => n12497,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_7_lut_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42516\,
            in3 => \N__42336\,
            lcout => n996,
            ltout => OPEN,
            carryin => n12497,
            carryout => n12498,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_8_lut_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52903\,
            in2 => \N__44987\,
            in3 => \N__42333\,
            lcout => n995,
            ltout => OPEN,
            carryin => n12498,
            carryout => n12499,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_9_lut_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__52904\,
            in1 => \N__42567\,
            in2 => \N__44964\,
            in3 => \N__42579\,
            lcout => n1026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i641_3_lut_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44757\,
            in2 => \N__42576\,
            in3 => \N__44952\,
            lcout => n1033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_167_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42515\,
            in3 => \N__42538\,
            lcout => OPEN,
            ltout => \n14466_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_169_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__44980\,
            in1 => \N__42566\,
            in2 => \N__42555\,
            in3 => \N__42552\,
            lcout => n960,
            ltout => \n960_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i637_3_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42539\,
            in2 => \N__42525\,
            in3 => \N__42522\,
            lcout => n1029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i636_3_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42511\,
            in2 => \N__42495\,
            in3 => \N__44954\,
            lcout => n1028,
            ltout => \n1028_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i703_3_lut_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46408\,
            in2 => \N__42486\,
            in3 => \N__45096\,
            lcout => n1127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i638_3_lut_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42483\,
            in2 => \N__42477\,
            in3 => \N__44953\,
            lcout => n1030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42456\,
            lcout => n17_adj_560,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10984_3_lut_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42870\,
            in2 => \N__42609\,
            in3 => \N__42846\,
            lcout => OPEN,
            ltout => \n13648_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10985_3_lut_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46173\,
            in2 => \N__42822\,
            in3 => \N__42819\,
            lcout => n832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i639_3_lut_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42762\,
            in2 => \N__42753\,
            in3 => \N__44955\,
            lcout => n1031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12441_3_lut_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42728\,
            in2 => \N__46199\,
            in3 => \N__42693\,
            lcout => n833,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42660\,
            lcout => n22_adj_555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_738_2_lut_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42645\,
            in3 => \N__42624\,
            lcout => n2542,
            ltout => OPEN,
            carryin => \bfn_12_25_0_\,
            carryout => n12482,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_738_3_lut_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52427\,
            in2 => \N__42621\,
            in3 => \N__42600\,
            lcout => n2541,
            ltout => OPEN,
            carryin => n12482,
            carryout => n12483,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_738_4_lut_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42597\,
            in3 => \N__42582\,
            lcout => n2540,
            ltout => OPEN,
            carryin => n12483,
            carryout => n12484,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_738_5_lut_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52428\,
            in2 => \N__43308\,
            in3 => \N__43293\,
            lcout => n2539,
            ltout => OPEN,
            carryin => n12484,
            carryout => n12485,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_738_6_lut_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43290\,
            in3 => \N__43272\,
            lcout => n2538,
            ltout => OPEN,
            carryin => n12485,
            carryout => n12486,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_738_7_lut_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43269\,
            in3 => \N__43257\,
            lcout => n2537,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43248\,
            lcout => n19_adj_558,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2112_3_lut_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43233\,
            in2 => \N__43197\,
            in3 => \N__43179\,
            lcout => n3208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i0_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42978\,
            in2 => \N__48825\,
            in3 => \N__42948\,
            lcout => duty_0,
            ltout => OPEN,
            carryin => \bfn_12_26_0_\,
            carryout => n12459,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i1_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42945\,
            in2 => \N__48792\,
            in3 => \N__42912\,
            lcout => duty_1,
            ltout => OPEN,
            carryin => n12459,
            carryout => n12460,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i2_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48756\,
            in2 => \N__42909\,
            in3 => \N__42873\,
            lcout => duty_2,
            ltout => OPEN,
            carryin => n12460,
            carryout => n12461,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i3_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43527\,
            in2 => \N__49170\,
            in3 => \N__43500\,
            lcout => duty_3,
            ltout => OPEN,
            carryin => n12461,
            carryout => n12462,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i4_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49137\,
            in2 => \N__43497\,
            in3 => \N__43461\,
            lcout => duty_4,
            ltout => OPEN,
            carryin => n12462,
            carryout => n12463,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i5_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43458\,
            in2 => \N__49104\,
            in3 => \N__43434\,
            lcout => duty_5,
            ltout => OPEN,
            carryin => n12463,
            carryout => n12464,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i6_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43431\,
            in2 => \N__49067\,
            in3 => \N__43407\,
            lcout => duty_6,
            ltout => OPEN,
            carryin => n12464,
            carryout => n12465,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i7_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49020\,
            in2 => \N__43404\,
            in3 => \N__43374\,
            lcout => duty_7,
            ltout => OPEN,
            carryin => n12465,
            carryout => n12466,
            clk => \N__55796\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i8_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43371\,
            in2 => \N__48984\,
            in3 => \N__43362\,
            lcout => duty_8,
            ltout => OPEN,
            carryin => \bfn_12_27_0_\,
            carryout => n12467,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i9_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43359\,
            in2 => \N__48945\,
            in3 => \N__43335\,
            lcout => duty_9,
            ltout => OPEN,
            carryin => n12467,
            carryout => n12468,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i10_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43332\,
            in2 => \N__48900\,
            in3 => \N__43311\,
            lcout => duty_10,
            ltout => OPEN,
            carryin => n12468,
            carryout => n12469,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i11_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43734\,
            in2 => \N__49488\,
            in3 => \N__43728\,
            lcout => duty_11,
            ltout => OPEN,
            carryin => n12469,
            carryout => n12470,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i12_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43725\,
            in2 => \N__49443\,
            in3 => \N__43716\,
            lcout => duty_12,
            ltout => OPEN,
            carryin => n12470,
            carryout => n12471,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i13_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43713\,
            in2 => \N__49392\,
            in3 => \N__43683\,
            lcout => duty_13,
            ltout => OPEN,
            carryin => n12471,
            carryout => n12472,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i14_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43680\,
            in2 => \N__49344\,
            in3 => \N__43656\,
            lcout => duty_14,
            ltout => OPEN,
            carryin => n12472,
            carryout => n12473,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i15_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54881\,
            in2 => \N__43653\,
            in3 => \N__43611\,
            lcout => duty_15,
            ltout => OPEN,
            carryin => n12473,
            carryout => n12474,
            clk => \N__55799\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i16_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43608\,
            in2 => \N__49296\,
            in3 => \N__43578\,
            lcout => duty_16,
            ltout => OPEN,
            carryin => \bfn_12_28_0_\,
            carryout => n12475,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i17_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43575\,
            in2 => \N__49257\,
            in3 => \N__43563\,
            lcout => duty_17,
            ltout => OPEN,
            carryin => n12475,
            carryout => n12476,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i18_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43560\,
            in2 => \N__49215\,
            in3 => \N__43530\,
            lcout => duty_18,
            ltout => OPEN,
            carryin => n12476,
            carryout => n12477,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i19_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43917\,
            in2 => \N__54810\,
            in3 => \N__43887\,
            lcout => duty_19,
            ltout => OPEN,
            carryin => n12477,
            carryout => n12478,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i20_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49590\,
            in2 => \N__43884\,
            in3 => \N__43875\,
            lcout => duty_20,
            ltout => OPEN,
            carryin => n12478,
            carryout => n12479,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i21_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43872\,
            in2 => \N__54852\,
            in3 => \N__43863\,
            lcout => duty_21,
            ltout => OPEN,
            carryin => n12479,
            carryout => n12480,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i22_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43860\,
            in2 => \N__49548\,
            in3 => \N__43833\,
            lcout => duty_22,
            ltout => OPEN,
            carryin => n12480,
            carryout => n12481,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i23_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54763\,
            in1 => \N__43830\,
            in2 => \_gnd_net_\,
            in3 => \N__43824\,
            lcout => duty_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i35_2_lut_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46558\,
            in2 => \_gnd_net_\,
            in3 => \N__43934\,
            lcout => n35,
            ltout => \n35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12540_4_lut_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43806\,
            in1 => \N__44064\,
            in2 => \N__43794\,
            in3 => \N__43791\,
            lcout => n15265,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i27_2_lut_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43782\,
            in2 => \_gnd_net_\,
            in3 => \N__46541\,
            lcout => n27_adj_671,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i12_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44093\,
            in1 => \N__55260\,
            in2 => \_gnd_net_\,
            in3 => \N__44076\,
            lcout => pwm_setpoint_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55808\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12553_3_lut_LC_12_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44063\,
            in1 => \N__44055\,
            in2 => \_gnd_net_\,
            in3 => \N__44031\,
            lcout => n15278,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12510_3_lut_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45270\,
            in1 => \N__47245\,
            in2 => \_gnd_net_\,
            in3 => \N__44022\,
            lcout => OPEN,
            ltout => \n15235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12511_3_lut_LC_12_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45471\,
            in2 => \N__44013\,
            in3 => \N__47744\,
            lcout => OPEN,
            ltout => \n15236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12455_3_lut_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__45458\,
            in1 => \_gnd_net_\,
            in2 => \N__44010\,
            in3 => \N__47723\,
            lcout => n15180,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i11_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55271\,
            in1 => \N__44006\,
            in2 => \_gnd_net_\,
            in3 => \N__43986\,
            lcout => pwm_setpoint_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i17_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55272\,
            in1 => \N__43973\,
            in2 => \_gnd_net_\,
            in3 => \N__43953\,
            lcout => pwm_setpoint_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55815\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12549_3_lut_LC_12_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45366\,
            in1 => \N__45348\,
            in2 => \_gnd_net_\,
            in3 => \N__43923\,
            lcout => n15274,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i8_3_lut_3_lut_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__47489\,
            in1 => \N__47364\,
            in2 => \_gnd_net_\,
            in3 => \N__47346\,
            lcout => OPEN,
            ltout => \n8_adj_657_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12494_4_lut_LC_12_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__44166\,
            in1 => \N__45390\,
            in2 => \N__44208\,
            in3 => \N__44193\,
            lcout => OPEN,
            ltout => \n15219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12530_4_lut_LC_12_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__44164\,
            in1 => \N__44205\,
            in2 => \N__44196\,
            in3 => \N__47706\,
            lcout => n15255,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i24_3_lut_LC_12_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44187\,
            in1 => \N__44163\,
            in2 => \_gnd_net_\,
            in3 => \N__44100\,
            lcout => n24_adj_669,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i45_2_lut_LC_12_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44186\,
            in2 => \_gnd_net_\,
            in3 => \N__46497\,
            lcout => n45,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12545_3_lut_LC_12_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45444\,
            in1 => \N__45432\,
            in2 => \_gnd_net_\,
            in3 => \N__44172\,
            lcout => OPEN,
            ltout => \n40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12532_4_lut_LC_12_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__44165\,
            in1 => \N__44148\,
            in2 => \N__44142\,
            in3 => \N__45414\,
            lcout => n15257,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i20_LC_12_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55309\,
            in1 => \N__44139\,
            in2 => \_gnd_net_\,
            in3 => \N__44121\,
            lcout => pwm_setpoint_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i22_1_lut_LC_12_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44312\,
            lcout => n4_adj_584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i16_3_lut_3_lut_LC_12_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__47188\,
            in1 => \N__45379\,
            in2 => \_gnd_net_\,
            in3 => \N__47306\,
            lcout => n16_adj_664,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2175_1_lut_LC_12_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55308\,
            lcout => \pwm_setpoint_23__N_195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_3_lut_LC_12_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111010"
        )
    port map (
            in0 => \N__47633\,
            in1 => \_gnd_net_\,
            in2 => \N__47598\,
            in3 => \N__47672\,
            lcout => n6_adj_717,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i21_LC_12_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44322\,
            in1 => \N__55310\,
            in2 => \_gnd_net_\,
            in3 => \N__44313\,
            lcout => pwm_setpoint_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_2_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45642\,
            in2 => \_gnd_net_\,
            in3 => \N__44286\,
            lcout => n1801,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => n12577,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_3_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52731\,
            in2 => \N__45665\,
            in3 => \N__44268\,
            lcout => n1800,
            ltout => OPEN,
            carryin => n12577,
            carryout => n12578,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45593\,
            in3 => \N__44253\,
            lcout => n1799,
            ltout => OPEN,
            carryin => n12578,
            carryout => n12579,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_5_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52732\,
            in2 => \N__45686\,
            in3 => \N__44241\,
            lcout => n1798,
            ltout => OPEN,
            carryin => n12579,
            carryout => n12580,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_6_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45536\,
            in3 => \N__44229\,
            lcout => n1797,
            ltout => OPEN,
            carryin => n12580,
            carryout => n12581,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_7_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45494\,
            in3 => \N__44211\,
            lcout => n1796,
            ltout => OPEN,
            carryin => n12581,
            carryout => n12582,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_8_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52734\,
            in2 => \N__50105\,
            in3 => \N__44469\,
            lcout => n1795,
            ltout => OPEN,
            carryin => n12582,
            carryout => n12583,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_9_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52733\,
            in2 => \N__49791\,
            in3 => \N__44454\,
            lcout => n1794,
            ltout => OPEN,
            carryin => n12583,
            carryout => n12584,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_10_lut_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52724\,
            in2 => \N__50339\,
            in3 => \N__44442\,
            lcout => n1793,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => n12585,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_11_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53085\,
            in2 => \N__50285\,
            in3 => \N__44427\,
            lcout => n1792,
            ltout => OPEN,
            carryin => n12585,
            carryout => n12586,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_12_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52725\,
            in2 => \N__50312\,
            in3 => \N__44415\,
            lcout => n1791,
            ltout => OPEN,
            carryin => n12586,
            carryout => n12587,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_13_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53086\,
            in2 => \N__50249\,
            in3 => \N__44400\,
            lcout => n1790,
            ltout => OPEN,
            carryin => n12587,
            carryout => n12588,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_14_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52726\,
            in2 => \N__44397\,
            in3 => \N__44376\,
            lcout => n1789,
            ltout => OPEN,
            carryin => n12588,
            carryout => n12589,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_15_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44372\,
            in2 => \N__53002\,
            in3 => \N__44343\,
            lcout => n1788,
            ltout => OPEN,
            carryin => n12589,
            carryout => n12590,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_16_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44579\,
            in2 => \N__53449\,
            in3 => \N__44553\,
            lcout => n1787,
            ltout => OPEN,
            carryin => n12590,
            carryout => n12591,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_17_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__52730\,
            in1 => \N__44543\,
            in2 => \N__47943\,
            in3 => \N__44526\,
            lcout => n1818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_2_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48223\,
            in3 => \N__44499\,
            lcout => n1601,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => n12550,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_3_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52721\,
            in2 => \N__45762\,
            in3 => \N__44496\,
            lcout => n1600,
            ltout => OPEN,
            carryin => n12550,
            carryout => n12551,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_4_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48168\,
            in3 => \N__44493\,
            lcout => n1599,
            ltout => OPEN,
            carryin => n12551,
            carryout => n12552,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_5_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52722\,
            in2 => \N__45557\,
            in3 => \N__44490\,
            lcout => n1598,
            ltout => OPEN,
            carryin => n12552,
            carryout => n12553,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_6_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50580\,
            in3 => \N__44487\,
            lcout => n1597,
            ltout => OPEN,
            carryin => n12553,
            carryout => n12554,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_7_lut_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50751\,
            in3 => \N__44484\,
            lcout => n1596,
            ltout => OPEN,
            carryin => n12554,
            carryout => n12555,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_8_lut_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52786\,
            in2 => \N__49987\,
            in3 => \N__44481\,
            lcout => n1595,
            ltout => OPEN,
            carryin => n12555,
            carryout => n12556,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_9_lut_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52723\,
            in2 => \N__50798\,
            in3 => \N__44649\,
            lcout => n1594,
            ltout => OPEN,
            carryin => n12556,
            carryout => n12557,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_10_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52711\,
            in2 => \N__50052\,
            in3 => \N__44646\,
            lcout => n1593,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => n12558,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_11_lut_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52713\,
            in2 => \N__48444\,
            in3 => \N__44643\,
            lcout => n1592,
            ltout => OPEN,
            carryin => n12558,
            carryout => n12559,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_12_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48416\,
            in2 => \N__53000\,
            in3 => \N__44634\,
            lcout => n1591,
            ltout => OPEN,
            carryin => n12559,
            carryout => n12560,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_13_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52717\,
            in2 => \N__47916\,
            in3 => \N__44631\,
            lcout => n1590,
            ltout => OPEN,
            carryin => n12560,
            carryout => n12561,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_14_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48263\,
            in2 => \N__53001\,
            in3 => \N__44628\,
            lcout => n1589,
            ltout => OPEN,
            carryin => n12561,
            carryout => n12562,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_15_lut_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__52712\,
            in1 => \N__45725\,
            in2 => \N__50820\,
            in3 => \N__44625\,
            lcout => n1620_adj_607,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i843_3_lut_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48606\,
            in2 => \N__48627\,
            in3 => \N__51590\,
            lcout => n1331,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i21_3_lut_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44622\,
            in1 => \N__46189\,
            in2 => \_gnd_net_\,
            in3 => \N__44610\,
            lcout => n299,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i7_3_lut_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46190\,
            in1 => \N__44904\,
            in2 => \_gnd_net_\,
            in3 => \N__44895\,
            lcout => n313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i23_3_lut_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44805\,
            in1 => \N__44817\,
            in2 => \_gnd_net_\,
            in3 => \N__46188\,
            lcout => n297,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44804\,
            lcout => n11_adj_632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i25_3_lut_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44730\,
            in1 => \N__44769\,
            in2 => \_gnd_net_\,
            in3 => \N__46187\,
            lcout => n295,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44729\,
            lcout => n9_adj_630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i640_3_lut_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__44691\,
            in1 => \_gnd_net_\,
            in2 => \N__44664\,
            in3 => \N__44956\,
            lcout => n1032,
            ltout => \n1032_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9947_3_lut_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__46266\,
            in1 => \_gnd_net_\,
            in2 => \N__44655\,
            in3 => \N__45934\,
            lcout => OPEN,
            ltout => \n11914_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_170_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__45133\,
            in1 => \N__45025\,
            in2 => \N__44652\,
            in3 => \N__45874\,
            lcout => OPEN,
            ltout => \n13716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12777_4_lut_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45107\,
            in1 => \N__45047\,
            in2 => \N__45000\,
            in3 => \N__45082\,
            lcout => n1059,
            ltout => \n1059_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i702_3_lut_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__45083\,
            in1 => \_gnd_net_\,
            in2 => \N__44997\,
            in3 => \N__45069\,
            lcout => n1126,
            ltout => \n1126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_171_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51787\,
            in2 => \N__44994\,
            in3 => \N__51748\,
            lcout => n14428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i704_3_lut_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45120\,
            in2 => \N__45140\,
            in3 => \N__46409\,
            lcout => n1128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i635_rep_55_3_lut_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__44991\,
            in1 => \_gnd_net_\,
            in2 => \N__44963\,
            in3 => \N__44925\,
            lcout => n1027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_2_lut_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46264\,
            in2 => \_gnd_net_\,
            in3 => \N__44919\,
            lcout => n1101,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => n12500,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_3_lut_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52557\,
            in2 => \N__45941\,
            in3 => \N__44916\,
            lcout => n1100,
            ltout => OPEN,
            carryin => n12500,
            carryout => n12501,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_4_lut_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45915\,
            in3 => \N__44913\,
            lcout => n1099,
            ltout => OPEN,
            carryin => n12501,
            carryout => n12502,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_5_lut_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52558\,
            in2 => \N__45875\,
            in3 => \N__44910\,
            lcout => n1098,
            ltout => OPEN,
            carryin => n12502,
            carryout => n12503,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_6_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45030\,
            in3 => \N__44907\,
            lcout => n1097,
            ltout => OPEN,
            carryin => n12503,
            carryout => n12504,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_7_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45141\,
            in3 => \N__45114\,
            lcout => n1096,
            ltout => OPEN,
            carryin => n12504,
            carryout => n12505,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_8_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52590\,
            in2 => \N__45111\,
            in3 => \N__45090\,
            lcout => n1095,
            ltout => OPEN,
            carryin => n12505,
            carryout => n12506,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_9_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52559\,
            in2 => \N__45087\,
            in3 => \N__45063\,
            lcout => n1094,
            ltout => OPEN,
            carryin => n12506,
            carryout => n12507,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_10_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52429\,
            in2 => \N__45057\,
            in3 => \N__45060\,
            lcout => n1093,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i701_3_lut_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45056\,
            in2 => \N__46424\,
            in3 => \N__45036\,
            lcout => n1125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i705_3_lut_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45029\,
            in2 => \N__45009\,
            in3 => \N__46414\,
            lcout => n1129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__49211\,
            in1 => \N__49388\,
            in2 => \N__49442\,
            in3 => \N__49340\,
            lcout => n23_adj_700,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.pwm_counter_661__i0_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45197\,
            in2 => \_gnd_net_\,
            in3 => \N__45183\,
            lcout => pwm_counter_0,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \PWM.n13056\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i1_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45179\,
            in2 => \_gnd_net_\,
            in3 => \N__45165\,
            lcout => pwm_counter_1,
            ltout => OPEN,
            carryin => \PWM.n13056\,
            carryout => \PWM.n13057\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i2_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46811\,
            in2 => \_gnd_net_\,
            in3 => \N__45162\,
            lcout => pwm_counter_2,
            ltout => OPEN,
            carryin => \PWM.n13057\,
            carryout => \PWM.n13058\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i3_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46793\,
            in2 => \_gnd_net_\,
            in3 => \N__45159\,
            lcout => pwm_counter_3,
            ltout => OPEN,
            carryin => \PWM.n13058\,
            carryout => \PWM.n13059\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i4_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47468\,
            in2 => \_gnd_net_\,
            in3 => \N__45156\,
            lcout => pwm_counter_4,
            ltout => OPEN,
            carryin => \PWM.n13059\,
            carryout => \PWM.n13060\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i5_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46772\,
            in2 => \_gnd_net_\,
            in3 => \N__45153\,
            lcout => pwm_counter_5,
            ltout => OPEN,
            carryin => \PWM.n13060\,
            carryout => \PWM.n13061\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i6_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46708\,
            in2 => \_gnd_net_\,
            in3 => \N__45150\,
            lcout => pwm_counter_6,
            ltout => OPEN,
            carryin => \PWM.n13061\,
            carryout => \PWM.n13062\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i7_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46741\,
            in2 => \_gnd_net_\,
            in3 => \N__45147\,
            lcout => pwm_counter_7,
            ltout => OPEN,
            carryin => \PWM.n13062\,
            carryout => \PWM.n13063\,
            clk => \N__55800\,
            ce => 'H',
            sr => \N__47118\
        );

    \PWM.pwm_counter_661__i8_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47338\,
            in2 => \_gnd_net_\,
            in3 => \N__45144\,
            lcout => pwm_counter_8,
            ltout => OPEN,
            carryin => \bfn_13_27_0_\,
            carryout => \PWM.n13064\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i9_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47269\,
            in2 => \_gnd_net_\,
            in3 => \N__45228\,
            lcout => pwm_counter_9,
            ltout => OPEN,
            carryin => \PWM.n13064\,
            carryout => \PWM.n13065\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i10_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46658\,
            in2 => \_gnd_net_\,
            in3 => \N__45225\,
            lcout => pwm_counter_10,
            ltout => OPEN,
            carryin => \PWM.n13065\,
            carryout => \PWM.n13066\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i11_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46679\,
            in2 => \_gnd_net_\,
            in3 => \N__45222\,
            lcout => pwm_counter_11,
            ltout => OPEN,
            carryin => \PWM.n13066\,
            carryout => \PWM.n13067\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i12_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47155\,
            in2 => \_gnd_net_\,
            in3 => \N__45219\,
            lcout => pwm_counter_12,
            ltout => OPEN,
            carryin => \PWM.n13067\,
            carryout => \PWM.n13068\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i13_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46537\,
            in2 => \_gnd_net_\,
            in3 => \N__45216\,
            lcout => pwm_counter_13,
            ltout => OPEN,
            carryin => \PWM.n13068\,
            carryout => \PWM.n13069\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i14_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46633\,
            in2 => \_gnd_net_\,
            in3 => \N__45213\,
            lcout => pwm_counter_14,
            ltout => OPEN,
            carryin => \PWM.n13069\,
            carryout => \PWM.n13070\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i15_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46444\,
            in2 => \_gnd_net_\,
            in3 => \N__45210\,
            lcout => pwm_counter_15,
            ltout => OPEN,
            carryin => \PWM.n13070\,
            carryout => \PWM.n13071\,
            clk => \N__55804\,
            ce => 'H',
            sr => \N__47110\
        );

    \PWM.pwm_counter_661__i16_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46590\,
            in2 => \_gnd_net_\,
            in3 => \N__45207\,
            lcout => pwm_counter_16,
            ltout => OPEN,
            carryin => \bfn_13_28_0_\,
            carryout => \PWM.n13072\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i17_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46560\,
            in2 => \_gnd_net_\,
            in3 => \N__45204\,
            lcout => pwm_counter_17,
            ltout => OPEN,
            carryin => \PWM.n13072\,
            carryout => \PWM.n13073\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i18_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46475\,
            in2 => \_gnd_net_\,
            in3 => \N__45255\,
            lcout => pwm_counter_18,
            ltout => OPEN,
            carryin => \PWM.n13073\,
            carryout => \PWM.n13074\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i19_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47087\,
            in2 => \_gnd_net_\,
            in3 => \N__45252\,
            lcout => pwm_counter_19,
            ltout => OPEN,
            carryin => \PWM.n13074\,
            carryout => \PWM.n13075\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i20_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46613\,
            in2 => \_gnd_net_\,
            in3 => \N__45249\,
            lcout => pwm_counter_20,
            ltout => OPEN,
            carryin => \PWM.n13075\,
            carryout => \PWM.n13076\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i21_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47179\,
            in2 => \_gnd_net_\,
            in3 => \N__45246\,
            lcout => pwm_counter_21,
            ltout => OPEN,
            carryin => \PWM.n13076\,
            carryout => \PWM.n13077\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i22_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46496\,
            in2 => \_gnd_net_\,
            in3 => \N__45243\,
            lcout => pwm_counter_22,
            ltout => OPEN,
            carryin => \PWM.n13077\,
            carryout => \PWM.n13078\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i23_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46514\,
            in2 => \_gnd_net_\,
            in3 => \N__45240\,
            lcout => pwm_counter_23,
            ltout => OPEN,
            carryin => \PWM.n13078\,
            carryout => \PWM.n13079\,
            clk => \N__55809\,
            ce => 'H',
            sr => \N__47109\
        );

    \PWM.pwm_counter_661__i24_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47052\,
            in2 => \_gnd_net_\,
            in3 => \N__45237\,
            lcout => pwm_counter_24,
            ltout => OPEN,
            carryin => \bfn_13_29_0_\,
            carryout => \PWM.n13080\,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \PWM.pwm_counter_661__i25_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46989\,
            in2 => \_gnd_net_\,
            in3 => \N__45234\,
            lcout => pwm_counter_25,
            ltout => OPEN,
            carryin => \PWM.n13080\,
            carryout => \PWM.n13081\,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \PWM.pwm_counter_661__i26_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47013\,
            in2 => \_gnd_net_\,
            in3 => \N__45231\,
            lcout => pwm_counter_26,
            ltout => OPEN,
            carryin => \PWM.n13081\,
            carryout => \PWM.n13082\,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \PWM.pwm_counter_661__i27_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47027\,
            in2 => \_gnd_net_\,
            in3 => \N__45333\,
            lcout => pwm_counter_27,
            ltout => OPEN,
            carryin => \PWM.n13082\,
            carryout => \PWM.n13083\,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \PWM.pwm_counter_661__i28_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46974\,
            in2 => \_gnd_net_\,
            in3 => \N__45330\,
            lcout => pwm_counter_28,
            ltout => OPEN,
            carryin => \PWM.n13083\,
            carryout => \PWM.n13084\,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \PWM.pwm_counter_661__i29_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47040\,
            in2 => \_gnd_net_\,
            in3 => \N__45327\,
            lcout => pwm_counter_29,
            ltout => OPEN,
            carryin => \PWM.n13084\,
            carryout => \PWM.n13085\,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \PWM.pwm_counter_661__i30_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47001\,
            in2 => \_gnd_net_\,
            in3 => \N__45324\,
            lcout => pwm_counter_30,
            ltout => OPEN,
            carryin => \PWM.n13085\,
            carryout => \PWM.n13086\,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \PWM.pwm_counter_661__i31_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46953\,
            in2 => \_gnd_net_\,
            in3 => \N__45321\,
            lcout => pwm_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55816\,
            ce => 'H',
            sr => \N__47111\
        );

    \commutation_state_i0_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__47637\,
            in1 => \N__47597\,
            in2 => \_gnd_net_\,
            in3 => \N__47690\,
            lcout => commutation_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55819\,
            ce => \N__45318\,
            sr => \N__47697\
        );

    \LessThan_299_i11_2_lut_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45302\,
            in2 => \_gnd_net_\,
            in3 => \N__46773\,
            lcout => n11_adj_660,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i13_2_lut_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45285\,
            in2 => \_gnd_net_\,
            in3 => \N__46709\,
            lcout => n13_adj_662,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i21_2_lut_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45269\,
            in2 => \_gnd_net_\,
            in3 => \N__46659\,
            lcout => n21_adj_667,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i23_2_lut_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46680\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45470\,
            lcout => n23_adj_668,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i25_2_lut_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45459\,
            in2 => \_gnd_net_\,
            in3 => \N__47157\,
            lcout => n25_adj_670,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i41_2_lut_LC_13_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45443\,
            in2 => \_gnd_net_\,
            in3 => \N__46614\,
            lcout => n41,
            ltout => \n41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12387_4_lut_LC_13_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__47757\,
            in1 => \N__45347\,
            in2 => \N__45426\,
            in3 => \N__45423\,
            lcout => n15112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.pwm_out_12_LC_13_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__46518\,
            in1 => \N__45408\,
            in2 => \_gnd_net_\,
            in3 => \N__45396\,
            lcout => pwm_out,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55824\,
            ce => 'H',
            sr => \N__46935\
        );

    \i12383_2_lut_4_lut_LC_13_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__47277\,
            in1 => \N__45381\,
            in2 => \N__47310\,
            in3 => \N__47190\,
            lcout => n15108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i43_2_lut_LC_13_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47189\,
            in2 => \_gnd_net_\,
            in3 => \N__45380\,
            lcout => n43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i39_2_lut_LC_13_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__45365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47088\,
            lcout => n39,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12878_1_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50170\,
            in3 => \_gnd_net_\,
            lcout => n15603,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1043_rep_35_3_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47802\,
            in2 => \N__49955\,
            in3 => \N__50144\,
            lcout => OPEN,
            ltout => \n14910_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12442_3_lut_4_lut_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__50145\,
            in1 => \N__49991\,
            in2 => \N__45540\,
            in3 => \N__50668\,
            lcout => n1726,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1107_3_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47787\,
            in1 => \_gnd_net_\,
            in2 => \N__47769\,
            in3 => \N__50146\,
            lcout => n1723,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1114_3_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__47841\,
            in1 => \_gnd_net_\,
            in2 => \N__50169\,
            in3 => \N__47861\,
            lcout => n1730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_76_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47786\,
            in1 => \N__45702\,
            in2 => \N__48125\,
            in3 => \N__50079\,
            lcout => OPEN,
            ltout => \n14514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12881_4_lut_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48026\,
            in1 => \N__48070\,
            in2 => \N__45510\,
            in3 => \N__47963\,
            lcout => n1653,
            ltout => \n1653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1117_3_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47511\,
            in2 => \N__45507\,
            in3 => \N__47544\,
            lcout => n1733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1046_3_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__45504\,
            in1 => \_gnd_net_\,
            in2 => \N__45558\,
            in3 => \N__50653\,
            lcout => n1630_adj_617,
            ltout => \n1630_adj_617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1113_3_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__50167\,
            in1 => \N__47817\,
            in2 => \N__45498\,
            in3 => \_gnd_net_\,
            lcout => n1729,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9935_3_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__47542\,
            in1 => \N__48181\,
            in2 => \_gnd_net_\,
            in3 => \N__47884\,
            lcout => OPEN,
            ltout => \n11902_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_75_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__47857\,
            in1 => \N__47828\,
            in2 => \N__45705\,
            in3 => \N__50554\,
            lcout => n13736,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1047_3_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45696\,
            in2 => \N__48167\,
            in3 => \N__50652\,
            lcout => n1631_adj_618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1115_3_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__50168\,
            in1 => \N__47871\,
            in2 => \N__47891\,
            in3 => \_gnd_net_\,
            lcout => n1731,
            ltout => \n1731_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10002_4_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__45658\,
            in1 => \N__45641\,
            in2 => \N__45612\,
            in3 => \N__45586\,
            lcout => n11970,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1116_3_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__50166\,
            in1 => \N__47499\,
            in2 => \N__48188\,
            in3 => \_gnd_net_\,
            lcout => n1732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1038_3_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47909\,
            in2 => \N__50662\,
            in3 => \N__45570\,
            lcout => n1622_adj_609,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i976_3_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51056\,
            in2 => \N__51400\,
            in3 => \N__51036\,
            lcout => n1528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1037_3_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45564\,
            in2 => \N__50661\,
            in3 => \N__48264\,
            lcout => n1621_adj_608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i979_3_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51387\,
            in1 => \N__50427\,
            in2 => \_gnd_net_\,
            in3 => \N__50453\,
            lcout => n1531,
            ltout => \n1531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10006_4_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__48224\,
            in1 => \N__45761\,
            in2 => \N__45774\,
            in3 => \N__48160\,
            lcout => n11974,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1040_3_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48440\,
            in2 => \N__45771\,
            in3 => \N__50633\,
            lcout => n1624_adj_611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i981_3_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50529\,
            in1 => \N__50502\,
            in2 => \_gnd_net_\,
            in3 => \N__51386\,
            lcout => n1533,
            ltout => \n1533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1048_3_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45747\,
            in2 => \N__45741\,
            in3 => \N__50632\,
            lcout => n1632_adj_619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i970_3_lut_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51391\,
            in1 => \_gnd_net_\,
            in2 => \N__50859\,
            in3 => \N__50879\,
            lcout => n1522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12857_1_lut_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50654\,
            lcout => n15582,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_72_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48436\,
            in1 => \N__48409\,
            in2 => \N__50051\,
            in3 => \N__45840\,
            lcout => OPEN,
            ltout => \n14294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_73_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__50575\,
            in1 => \N__50746\,
            in2 => \N__45714\,
            in3 => \N__45711\,
            lcout => n14296,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i975_3_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51016\,
            in2 => \N__51401\,
            in3 => \N__50994\,
            lcout => n1527,
            ltout => \n1527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_71_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45843\,
            in3 => \N__49977\,
            lcout => n14288,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i909_3_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48305\,
            in2 => \N__48285\,
            in3 => \N__51281\,
            lcout => n1429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i20_3_lut_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45816\,
            in1 => \N__45834\,
            in2 => \_gnd_net_\,
            in3 => \N__46191\,
            lcout => n300,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i842_3_lut_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48591\,
            in2 => \N__51601\,
            in3 => \N__51638\,
            lcout => n1330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i908_3_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__48725\,
            in1 => \_gnd_net_\,
            in2 => \N__51287\,
            in3 => \N__48273\,
            lcout => n1428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i910_3_lut_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48315\,
            in2 => \N__48341\,
            in3 => \N__51266\,
            lcout => n1430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i836_3_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__48855\,
            in1 => \_gnd_net_\,
            in2 => \N__51602\,
            in3 => \N__52200\,
            lcout => n1324,
            ltout => \n1324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i903_3_lut_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48522\,
            in2 => \N__45819\,
            in3 => \N__51270\,
            lcout => n1423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45815\,
            lcout => n14_adj_635,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i707_3_lut_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45914\,
            in2 => \N__45900\,
            in3 => \N__46410\,
            lcout => n1131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9941_3_lut_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__48391\,
            in1 => \_gnd_net_\,
            in2 => \N__48482\,
            in3 => \N__48703\,
            lcout => OPEN,
            ltout => \n11908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_176_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__48304\,
            in1 => \N__48334\,
            in2 => \N__45891\,
            in3 => \N__48721\,
            lcout => OPEN,
            ltout => \n13708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12822_4_lut_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48533\,
            in1 => \N__48839\,
            in2 => \N__45888\,
            in3 => \N__51075\,
            lcout => n1356,
            ltout => \n1356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i912_3_lut_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__48704\,
            in1 => \N__48363\,
            in2 => \N__45885\,
            in3 => \_gnd_net_\,
            lcout => n1432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12819_1_lut_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51277\,
            in3 => \_gnd_net_\,
            lcout => n15544,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i913_3_lut_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48392\,
            in2 => \N__48375\,
            in3 => \N__51248\,
            lcout => n1433,
            ltout => \n1433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9939_3_lut_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__50521\,
            in1 => \_gnd_net_\,
            in2 => \N__45882\,
            in3 => \N__50443\,
            lcout => n11906,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i706_3_lut_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45879\,
            in2 => \N__46420\,
            in3 => \N__45849\,
            lcout => n1130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i709_3_lut_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46265\,
            in2 => \N__46239\,
            in3 => \N__46404\,
            lcout => n1133,
            ltout => \n1133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10032_4_lut_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__51913\,
            in1 => \N__51463\,
            in2 => \N__46227\,
            in3 => \N__51953\,
            lcout => OPEN,
            ltout => \n12000_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12791_4_lut_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__52337\,
            in1 => \N__46224\,
            in2 => \N__46218\,
            in3 => \N__46341\,
            lcout => n1158,
            ltout => \n1158_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i777_3_lut_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__51441\,
            in1 => \N__51464\,
            in2 => \N__46215\,
            in3 => \_gnd_net_\,
            lcout => n1233,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i776_3_lut_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51969\,
            in2 => \N__51429\,
            in3 => \N__52239\,
            lcout => n1232,
            ltout => \n1232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9943_3_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48685\,
            in2 => \N__46212\,
            in3 => \N__48655\,
            lcout => n11910,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i22_3_lut_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46209\,
            in1 => \N__46194\,
            in2 => \_gnd_net_\,
            in3 => \N__46335\,
            lcout => n298,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i708_3_lut_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45954\,
            in2 => \N__45948\,
            in3 => \N__46418\,
            lcout => n1132,
            ltout => \n1132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i775_3_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52240\,
            in2 => \N__45918\,
            in3 => \N__51939\,
            lcout => n1231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12774_1_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46419\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n15499,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_53_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49249\,
            in1 => \N__54764\,
            in2 => \N__49589\,
            in3 => \N__49484\,
            lcout => n24_adj_561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_172_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51874\,
            in3 => \N__51824\,
            lcout => n14470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46327\,
            lcout => n12_adj_633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__49537\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49470\,
            lcout => OPEN,
            ltout => \n16_adj_701_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__49585\,
            in1 => \N__49289\,
            in2 => \N__46290\,
            in3 => \N__46872\,
            lcout => n25_adj_698,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48888\,
            in1 => \N__49008\,
            in2 => \N__49056\,
            in3 => \N__48972\,
            lcout => n10_adj_567,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i828_4_lut_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__46857\,
            in1 => \N__46287\,
            in2 => \N__54765\,
            in3 => \N__46278\,
            lcout => \direction_N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49156\,
            in1 => \N__48811\,
            in2 => \N__48784\,
            in3 => \N__48745\,
            lcout => OPEN,
            ltout => \n13932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49090\,
            in2 => \N__46269\,
            in3 => \N__49126\,
            lcout => OPEN,
            ltout => \n14110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_49_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__49242\,
            in1 => \N__48927\,
            in2 => \N__46881\,
            in3 => \N__46878\,
            lcout => n15_adj_702,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9888_2_lut_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49089\,
            in2 => \_gnd_net_\,
            in3 => \N__49125\,
            lcout => n11853,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_adj_54_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49194\,
            in1 => \N__49281\,
            in2 => \N__49333\,
            in3 => \N__54873\,
            lcout => n23_adj_562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12425_3_lut_4_lut_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__46848\,
            in1 => \N__46827\,
            in2 => \N__46812\,
            in3 => \N__46789\,
            lcout => n15150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i2_3_lut_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__46771\,
            in1 => \N__46740\,
            in2 => \_gnd_net_\,
            in3 => \N__46707\,
            lcout => \PWM.n13995\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i11_4_lut_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46678\,
            in1 => \N__46657\,
            in2 => \N__46638\,
            in3 => \N__46612\,
            lcout => \PWM.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i12_4_lut_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46589\,
            in1 => \N__46559\,
            in2 => \N__46542\,
            in3 => \N__46513\,
            lcout => \PWM.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i10_4_lut_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46495\,
            in1 => \N__46474\,
            in2 => \N__46455\,
            in3 => \N__47178\,
            lcout => OPEN,
            ltout => \PWM.n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i13_4_lut_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47156\,
            in1 => \N__47058\,
            in2 => \N__47136\,
            in3 => \N__46962\,
            lcout => OPEN,
            ltout => \PWM.n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i9624_4_lut_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__46952\,
            in1 => \N__47133\,
            in2 => \N__47127\,
            in3 => \N__47124\,
            lcout => \PWM.pwm_counter_31__N_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i1_4_lut_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__47086\,
            in1 => \N__47337\,
            in2 => \N__47067\,
            in3 => \N__47268\,
            lcout => \PWM.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47051\,
            in1 => \N__47039\,
            in2 => \N__47028\,
            in3 => \N__47012\,
            lcout => OPEN,
            ltout => \n12_adj_566_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47000\,
            in1 => \N__46988\,
            in2 => \N__46977\,
            in3 => \N__46973\,
            lcout => n5162,
            ltout => \n5162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46956\,
            in3 => \N__46951\,
            lcout => n5164,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i8_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55322\,
            in1 => \N__46923\,
            in2 => \_gnd_net_\,
            in3 => \N__46907\,
            lcout => pwm_setpoint_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55820\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i9_2_lut_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47490\,
            in2 => \_gnd_net_\,
            in3 => \N__47469\,
            lcout => n9_adj_658,
            ltout => \n9_adj_658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12480_4_lut_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__47454\,
            in1 => \N__47435\,
            in2 => \N__47424\,
            in3 => \N__47417\,
            lcout => n15205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12476_4_lut_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__47210\,
            in1 => \N__47228\,
            in2 => \N__47403\,
            in3 => \N__47388\,
            lcout => OPEN,
            ltout => \n15201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12536_4_lut_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47743\,
            in1 => \N__47722\,
            in2 => \N__47382\,
            in3 => \N__47246\,
            lcout => n15261,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i17_2_lut_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47357\,
            in2 => \_gnd_net_\,
            in3 => \N__47345\,
            lcout => n17_adj_665,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i19_2_lut_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47305\,
            in2 => \_gnd_net_\,
            in3 => \N__47276\,
            lcout => n19_adj_666,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12380_2_lut_4_lut_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000010"
        )
    port map (
            in0 => \N__49764\,
            in1 => \N__54693\,
            in2 => \N__54637\,
            in3 => \N__56100\,
            lcout => n15088,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12416_2_lut_4_lut_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000100000000"
        )
    port map (
            in0 => \N__56099\,
            in1 => \N__54624\,
            in2 => \N__54699\,
            in3 => \N__49610\,
            lcout => n15091,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12407_4_lut_LC_14_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__47247\,
            in1 => \N__47229\,
            in2 => \N__47217\,
            in3 => \N__47199\,
            lcout => OPEN,
            ltout => \n15132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12385_4_lut_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__47756\,
            in1 => \N__47745\,
            in2 => \N__47727\,
            in3 => \N__47724\,
            lcout => n15110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12420_2_lut_4_lut_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__54684\,
            in1 => \N__56101\,
            in2 => \N__54636\,
            in3 => \N__49735\,
            lcout => n15095,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i1_LC_14_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001100010000"
        )
    port map (
            in0 => \N__47635\,
            in1 => \N__47689\,
            in2 => \N__56029\,
            in3 => \N__47586\,
            lcout => commutation_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_14_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__47585\,
            in1 => \N__47685\,
            in2 => \_gnd_net_\,
            in3 => \N__47634\,
            lcout => \commutation_state_7__N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12419_2_lut_4_lut_LC_14_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__56118\,
            in1 => \N__54623\,
            in2 => \N__49703\,
            in3 => \N__54671\,
            lcout => n15094,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i2_LC_14_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001000110010"
        )
    port map (
            in0 => \N__47691\,
            in1 => \N__47636\,
            in2 => \N__55950\,
            in3 => \N__47596\,
            lcout => commutation_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55829\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_2_lut_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47543\,
            in2 => \_gnd_net_\,
            in3 => \N__47502\,
            lcout => n1701,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => n12563,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_3_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54188\,
            in2 => \N__48192\,
            in3 => \N__47493\,
            lcout => n1700,
            ltout => OPEN,
            carryin => n12563,
            carryout => n12564,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_4_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47895\,
            in3 => \N__47865\,
            lcout => n1699,
            ltout => OPEN,
            carryin => n12564,
            carryout => n12565,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_5_lut_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54189\,
            in2 => \N__47862\,
            in3 => \N__47835\,
            lcout => n1698,
            ltout => OPEN,
            carryin => n12565,
            carryout => n12566,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_6_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47832\,
            in3 => \N__47811\,
            lcout => n1697,
            ltout => OPEN,
            carryin => n12566,
            carryout => n12567,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_7_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50555\,
            in3 => \N__47808\,
            lcout => n1696,
            ltout => OPEN,
            carryin => n12567,
            carryout => n12568,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_8_lut_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54190\,
            in2 => \N__50711\,
            in3 => \N__47805\,
            lcout => n1695,
            ltout => OPEN,
            carryin => n12568,
            carryout => n12569,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_9_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49928\,
            in2 => \N__54359\,
            in3 => \N__47796\,
            lcout => n1694,
            ltout => OPEN,
            carryin => n12569,
            carryout => n12570,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_10_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53090\,
            in2 => \N__50769\,
            in3 => \N__47793\,
            lcout => n1693_adj_621,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => n12571,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_11_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53095\,
            in2 => \N__50012\,
            in3 => \N__47790\,
            lcout => n1692,
            ltout => OPEN,
            carryin => n12571,
            carryout => n12572,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_12_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47785\,
            in2 => \N__53451\,
            in3 => \N__47760\,
            lcout => n1691,
            ltout => OPEN,
            carryin => n12572,
            carryout => n12573,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_13_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53099\,
            in2 => \N__48126\,
            in3 => \N__48075\,
            lcout => n1690,
            ltout => OPEN,
            carryin => n12573,
            carryout => n12574,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_14_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53091\,
            in2 => \N__48071\,
            in3 => \N__48030\,
            lcout => n1689,
            ltout => OPEN,
            carryin => n12574,
            carryout => n12575,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_15_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48022\,
            in2 => \N__53450\,
            in3 => \N__47991\,
            lcout => n1688,
            ltout => OPEN,
            carryin => n12575,
            carryout => n12576,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_16_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53100\,
            in1 => \N__47981\,
            in2 => \N__47970\,
            in3 => \N__47946\,
            lcout => n1719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1108_3_lut_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47922\,
            in2 => \N__50013\,
            in3 => \N__50165\,
            lcout => n1724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i978_3_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50414\,
            in2 => \N__51398\,
            in3 => \N__50394\,
            lcout => n1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i911_3_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48354\,
            in2 => \N__48486\,
            in3 => \N__51282\,
            lcout => n1431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i971_3_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51212\,
            in2 => \N__51399\,
            in3 => \N__50895\,
            lcout => n1523,
            ltout => \n1523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12860_4_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50813\,
            in1 => \N__48262\,
            in2 => \N__48246\,
            in3 => \N__48243\,
            lcout => n1554,
            ltout => \n1554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1049_3_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__48237\,
            in1 => \_gnd_net_\,
            in2 => \N__48228\,
            in3 => \N__48225\,
            lcout => n1633_adj_620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i977_3_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50355\,
            in2 => \N__50385\,
            in3 => \N__51379\,
            lcout => n1529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i980_3_lut_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50466\,
            in2 => \N__50490\,
            in3 => \N__51375\,
            lcout => n1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_178_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__50410\,
            in1 => \N__51055\,
            in2 => \N__48141\,
            in3 => \N__50371\,
            lcout => n13727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i906_3_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51120\,
            in2 => \N__51295\,
            in3 => \N__48561\,
            lcout => n1426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i905_3_lut_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__48552\,
            in1 => \_gnd_net_\,
            in2 => \N__51099\,
            in3 => \N__51283\,
            lcout => n1425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_177_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51020\,
            in3 => \N__50978\,
            lcout => OPEN,
            ltout => \n14490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_179_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50920\,
            in1 => \N__50947\,
            in2 => \N__48129\,
            in3 => \N__51211\,
            lcout => OPEN,
            ltout => \n14496_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12841_4_lut_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__50875\,
            in1 => \N__48456\,
            in2 => \N__48450\,
            in3 => \N__50840\,
            lcout => n1455,
            ltout => \n1455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i973_3_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50948\,
            in2 => \N__48447\,
            in3 => \N__50934\,
            lcout => n1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i972_3_lut_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50921\,
            in2 => \N__50907\,
            in3 => \N__51392\,
            lcout => n1524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_2_lut_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48393\,
            in2 => \_gnd_net_\,
            in3 => \N__48366\,
            lcout => n1401,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => n12527,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_3_lut_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53196\,
            in2 => \N__48705\,
            in3 => \N__48357\,
            lcout => n1400,
            ltout => OPEN,
            carryin => n12527,
            carryout => n12528,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_4_lut_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48481\,
            in3 => \N__48345\,
            lcout => n1399,
            ltout => OPEN,
            carryin => n12528,
            carryout => n12529,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_5_lut_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53197\,
            in2 => \N__48342\,
            in3 => \N__48309\,
            lcout => n1398,
            ltout => OPEN,
            carryin => n12529,
            carryout => n12530,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_6_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48306\,
            in3 => \N__48276\,
            lcout => n1397,
            ltout => OPEN,
            carryin => n12530,
            carryout => n12531,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_7_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48726\,
            in3 => \N__48267\,
            lcout => n1396,
            ltout => OPEN,
            carryin => n12531,
            carryout => n12532,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_8_lut_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53198\,
            in2 => \N__51137\,
            in3 => \N__48564\,
            lcout => n1395,
            ltout => OPEN,
            carryin => n12532,
            carryout => n12533,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_9_lut_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51119\,
            in2 => \N__53576\,
            in3 => \N__48555\,
            lcout => n1394,
            ltout => OPEN,
            carryin => n12533,
            carryout => n12534,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_10_lut_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52898\,
            in2 => \N__51098\,
            in3 => \N__48543\,
            lcout => n1393,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => n12535,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_11_lut_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52979\,
            in2 => \N__51687\,
            in3 => \N__48540\,
            lcout => n1392,
            ltout => OPEN,
            carryin => n12535,
            carryout => n12536,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_12_lut_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52899\,
            in2 => \N__48537\,
            in3 => \N__48516\,
            lcout => n1391,
            ltout => OPEN,
            carryin => n12536,
            carryout => n12537,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_13_lut_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__52900\,
            in1 => \N__48840\,
            in2 => \N__48506\,
            in3 => \N__48489\,
            lcout => n1422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i771_3_lut_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52245\,
            in2 => \N__51803\,
            in3 => \N__51771\,
            lcout => n1227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i844_3_lut_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__48659\,
            in1 => \_gnd_net_\,
            in2 => \N__48639\,
            in3 => \N__51582\,
            lcout => n1332,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i841_3_lut_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48579\,
            in2 => \N__51597\,
            in3 => \N__51488\,
            lcout => n1329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i845_3_lut_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48669\,
            in1 => \N__48687\,
            in2 => \_gnd_net_\,
            in3 => \N__51581\,
            lcout => n1333,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_2_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48686\,
            in2 => \_gnd_net_\,
            in3 => \N__48663\,
            lcout => n1301,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => n12517,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_3_lut_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52973\,
            in2 => \N__48660\,
            in3 => \N__48630\,
            lcout => n1300,
            ltout => OPEN,
            carryin => n12517,
            carryout => n12518,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_4_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48623\,
            in3 => \N__48594\,
            lcout => n1299,
            ltout => OPEN,
            carryin => n12518,
            carryout => n12519,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_5_lut_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52974\,
            in2 => \N__51637\,
            in3 => \N__48582\,
            lcout => n1298,
            ltout => OPEN,
            carryin => n12519,
            carryout => n12520,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_6_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51489\,
            in3 => \N__48573\,
            lcout => n1297,
            ltout => OPEN,
            carryin => n12520,
            carryout => n12521,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_7_lut_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51669\,
            in3 => \N__48570\,
            lcout => n1296,
            ltout => OPEN,
            carryin => n12521,
            carryout => n12522,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_8_lut_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52975\,
            in2 => \N__51507\,
            in3 => \N__48567\,
            lcout => n1295,
            ltout => OPEN,
            carryin => n12522,
            carryout => n12523,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_9_lut_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51166\,
            in2 => \N__53339\,
            in3 => \N__48861\,
            lcout => n1294,
            ltout => OPEN,
            carryin => n12523,
            carryout => n12524,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_10_lut_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52891\,
            in2 => \N__51720\,
            in3 => \N__48858\,
            lcout => n1293,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => n12525,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_11_lut_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52971\,
            in2 => \N__52196\,
            in3 => \N__48846\,
            lcout => n1292,
            ltout => OPEN,
            carryin => n12525,
            carryout => n12526,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_12_lut_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__52972\,
            in1 => \N__51521\,
            in2 => \N__52323\,
            in3 => \N__48843\,
            lcout => n1323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12788_1_lut_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52241\,
            lcout => n15513,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_305_1_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52035\,
            in2 => \N__52082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => n12435,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i0_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48815\,
            in2 => \N__52146\,
            in3 => \N__48795\,
            lcout => encoder0_position_target_0,
            ltout => OPEN,
            carryin => n12435,
            carryout => n12436,
            clk => \N__55805\,
            ce => \N__55399\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i1_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52036\,
            in2 => \N__48788\,
            in3 => \N__48759\,
            lcout => encoder0_position_target_1,
            ltout => OPEN,
            carryin => n12436,
            carryout => n12437,
            clk => \N__55805\,
            ce => \N__55399\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i2_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52042\,
            in2 => \N__48755\,
            in3 => \N__48729\,
            lcout => encoder0_position_target_2,
            ltout => OPEN,
            carryin => n12437,
            carryout => n12438,
            clk => \N__55805\,
            ce => \N__55399\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i3_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52037\,
            in2 => \N__49166\,
            in3 => \N__49140\,
            lcout => encoder0_position_target_3,
            ltout => OPEN,
            carryin => n12438,
            carryout => n12439,
            clk => \N__55805\,
            ce => \N__55399\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i4_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52043\,
            in2 => \N__49136\,
            in3 => \N__49107\,
            lcout => encoder0_position_target_4,
            ltout => OPEN,
            carryin => n12439,
            carryout => n12440,
            clk => \N__55805\,
            ce => \N__55399\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i5_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52038\,
            in2 => \N__49100\,
            in3 => \N__49071\,
            lcout => encoder0_position_target_5,
            ltout => OPEN,
            carryin => n12440,
            carryout => n12441,
            clk => \N__55805\,
            ce => \N__55399\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i6_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52044\,
            in2 => \N__49057\,
            in3 => \N__49023\,
            lcout => encoder0_position_target_6,
            ltout => OPEN,
            carryin => n12441,
            carryout => n12442,
            clk => \N__55805\,
            ce => \N__55399\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i7_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52045\,
            in2 => \N__49018\,
            in3 => \N__48987\,
            lcout => encoder0_position_target_7,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => n12443,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i8_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48976\,
            in2 => \N__52083\,
            in3 => \N__48948\,
            lcout => encoder0_position_target_8,
            ltout => OPEN,
            carryin => n12443,
            carryout => n12444,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i9_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52049\,
            in2 => \N__48941\,
            in3 => \N__48903\,
            lcout => encoder0_position_target_9,
            ltout => OPEN,
            carryin => n12444,
            carryout => n12445,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i10_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48889\,
            in2 => \N__52084\,
            in3 => \N__48864\,
            lcout => encoder0_position_target_10,
            ltout => OPEN,
            carryin => n12445,
            carryout => n12446,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i11_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52053\,
            in2 => \N__49483\,
            in3 => \N__49446\,
            lcout => encoder0_position_target_11,
            ltout => OPEN,
            carryin => n12446,
            carryout => n12447,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i12_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49425\,
            in2 => \N__52085\,
            in3 => \N__49395\,
            lcout => encoder0_position_target_12,
            ltout => OPEN,
            carryin => n12447,
            carryout => n12448,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i13_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52057\,
            in2 => \N__49387\,
            in3 => \N__49347\,
            lcout => encoder0_position_target_13,
            ltout => OPEN,
            carryin => n12448,
            carryout => n12449,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i14_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49332\,
            in2 => \N__52086\,
            in3 => \N__49302\,
            lcout => encoder0_position_target_14,
            ltout => OPEN,
            carryin => n12449,
            carryout => n12450,
            clk => \N__55810\,
            ce => \N__55389\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i15_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52087\,
            in2 => \N__54882\,
            in3 => \N__49299\,
            lcout => encoder0_position_target_15,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => n12451,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i16_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49288\,
            in2 => \N__52106\,
            in3 => \N__49260\,
            lcout => encoder0_position_target_16,
            ltout => OPEN,
            carryin => n12451,
            carryout => n12452,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i17_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52091\,
            in2 => \N__49253\,
            in3 => \N__49218\,
            lcout => encoder0_position_target_17,
            ltout => OPEN,
            carryin => n12452,
            carryout => n12453,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i18_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49207\,
            in2 => \N__52107\,
            in3 => \N__49176\,
            lcout => encoder0_position_target_18,
            ltout => OPEN,
            carryin => n12453,
            carryout => n12454,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i19_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52095\,
            in2 => \N__54805\,
            in3 => \N__49173\,
            lcout => encoder0_position_target_19,
            ltout => OPEN,
            carryin => n12454,
            carryout => n12455,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i20_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49581\,
            in2 => \N__52108\,
            in3 => \N__49554\,
            lcout => encoder0_position_target_20,
            ltout => OPEN,
            carryin => n12455,
            carryout => n12456,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i21_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52099\,
            in2 => \N__54847\,
            in3 => \N__49551\,
            lcout => encoder0_position_target_21,
            ltout => OPEN,
            carryin => n12456,
            carryout => n12457,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i22_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49533\,
            in2 => \N__52109\,
            in3 => \N__49506\,
            lcout => encoder0_position_target_22,
            ltout => OPEN,
            carryin => n12457,
            carryout => n12458,
            clk => \N__55817\,
            ce => \N__55402\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i23_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52110\,
            in1 => \N__54755\,
            in2 => \_gnd_net_\,
            in3 => \N__49503\,
            lcout => encoder0_position_target_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55821\,
            ce => \N__55404\,
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_60_LC_15_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49699\,
            in2 => \_gnd_net_\,
            in3 => \N__49736\,
            lcout => n10_adj_719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12417_2_lut_4_lut_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000100"
        )
    port map (
            in0 => \N__56110\,
            in1 => \N__49639\,
            in2 => \N__54638\,
            in3 => \N__54688\,
            lcout => n15092,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_61_LC_15_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49609\,
            in1 => \N__49861\,
            in2 => \N__49643\,
            in3 => \N__49840\,
            lcout => OPEN,
            ltout => \n14_adj_718_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_15_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49666\,
            in1 => \N__49762\,
            in2 => \N__49500\,
            in3 => \N__49497\,
            lcout => n5119,
            ltout => \n5119_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9549_2_lut_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__55029\,
            in1 => \_gnd_net_\,
            in2 => \N__49491\,
            in3 => \_gnd_net_\,
            lcout => n11514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12422_2_lut_4_lut_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000010"
        )
    port map (
            in0 => \N__49862\,
            in1 => \N__56112\,
            in2 => \N__54698\,
            in3 => \N__54634\,
            lcout => n15089,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12418_2_lut_4_lut_LC_15_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000100"
        )
    port map (
            in0 => \N__56111\,
            in1 => \N__49667\,
            in2 => \N__54639\,
            in3 => \N__54689\,
            lcout => n15093,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i0_LC_15_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__49773\,
            in1 => \N__49763\,
            in2 => \N__54576\,
            in3 => \N__49746\,
            lcout => dti_counter_0,
            ltout => OPEN,
            carryin => \bfn_15_31_0_\,
            carryout => n12961,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i1_LC_15_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__49743\,
            in1 => \N__49737\,
            in2 => \N__49909\,
            in3 => \N__49713\,
            lcout => dti_counter_1,
            ltout => OPEN,
            carryin => n12961,
            carryout => n12962,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i2_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__49710\,
            in1 => \N__49899\,
            in2 => \N__49704\,
            in3 => \N__49677\,
            lcout => dti_counter_2,
            ltout => OPEN,
            carryin => n12962,
            carryout => n12963,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i3_LC_15_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__49674\,
            in1 => \N__49668\,
            in2 => \N__49910\,
            in3 => \N__49653\,
            lcout => dti_counter_3,
            ltout => OPEN,
            carryin => n12963,
            carryout => n12964,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i4_LC_15_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__49650\,
            in1 => \N__49903\,
            in2 => \N__49644\,
            in3 => \N__49620\,
            lcout => dti_counter_4,
            ltout => OPEN,
            carryin => n12964,
            carryout => n12965,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i5_LC_15_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__49617\,
            in1 => \N__49611\,
            in2 => \N__49911\,
            in3 => \N__49593\,
            lcout => dti_counter_5,
            ltout => OPEN,
            carryin => n12965,
            carryout => n12966,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i6_LC_15_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__49824\,
            in1 => \N__49907\,
            in2 => \N__49845\,
            in3 => \N__49914\,
            lcout => dti_counter_6,
            ltout => OPEN,
            carryin => n12966,
            carryout => n12967,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_659__i7_LC_15_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__49908\,
            in1 => \N__49878\,
            in2 => \N__49869\,
            in3 => \N__49872\,
            lcout => dti_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55830\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_62_LC_15_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__49812\,
            in1 => \N__55920\,
            in2 => \N__56017\,
            in3 => \N__49818\,
            lcout => n4_adj_716,
            ltout => \n4_adj_716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12404_2_lut_4_lut_LC_15_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__54670\,
            in1 => \N__56124\,
            in2 => \N__49848\,
            in3 => \N__49841\,
            lcout => n15090,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i0_LC_15_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => commutation_state_prev_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i1_LC_15_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => commutation_state_prev_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i2_LC_15_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__55921\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => commutation_state_prev_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55831\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1109_3_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50765\,
            in2 => \N__50186\,
            in3 => \N__49806\,
            lcout => n1725,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1111_3_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49800\,
            in2 => \N__50712\,
            in3 => \N__50175\,
            lcout => n1727,
            ltout => \n1727_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_77_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50092\,
            in2 => \N__50346\,
            in3 => \N__50338\,
            lcout => OPEN,
            ltout => \n14166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_78_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50299\,
            in1 => \N__50267\,
            in2 => \N__50256\,
            in3 => \N__50248\,
            lcout => n14172,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1112_3_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50208\,
            in2 => \N__50556\,
            in3 => \N__50171\,
            lcout => n1728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_74_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50764\,
            in1 => \N__50704\,
            in2 => \N__49929\,
            in3 => \N__50005\,
            lcout => n14508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i907_3_lut_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__51138\,
            in1 => \_gnd_net_\,
            in2 => \N__50070\,
            in3 => \N__51294\,
            lcout => n1427,
            ltout => \n1427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i974_3_lut_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50961\,
            in2 => \N__50055\,
            in3 => \N__51397\,
            lcout => n1526,
            ltout => \n1526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1041_3_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50648\,
            in2 => \N__50028\,
            in3 => \N__50025\,
            lcout => n1625_adj_612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1043_3_lut_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49992\,
            in2 => \N__49956\,
            in3 => \N__50647\,
            lcout => n1627_adj_614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1042_3_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50802\,
            in2 => \N__50667\,
            in3 => \N__50781\,
            lcout => n1626_adj_613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50747\,
            in2 => \N__50727\,
            in3 => \N__50646\,
            lcout => n1628_adj_615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1045_3_lut_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50688\,
            in2 => \N__50666\,
            in3 => \N__50576\,
            lcout => n1629_adj_616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_2_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50528\,
            in2 => \_gnd_net_\,
            in3 => \N__50493\,
            lcout => n1501,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => n12538,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_3_lut_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53609\,
            in2 => \N__50489\,
            in3 => \N__50460\,
            lcout => n1500,
            ltout => OPEN,
            carryin => n12538,
            carryout => n12539,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_4_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50457\,
            in3 => \N__50418\,
            lcout => n1499,
            ltout => OPEN,
            carryin => n12539,
            carryout => n12540,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_5_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53610\,
            in2 => \N__50415\,
            in3 => \N__50388\,
            lcout => n1498,
            ltout => OPEN,
            carryin => n12540,
            carryout => n12541,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_6_lut_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50384\,
            in3 => \N__50349\,
            lcout => n1497,
            ltout => OPEN,
            carryin => n12541,
            carryout => n12542,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_7_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51063\,
            in3 => \N__51027\,
            lcout => n1496,
            ltout => OPEN,
            carryin => n12542,
            carryout => n12543,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_8_lut_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53615\,
            in2 => \N__51024\,
            in3 => \N__50982\,
            lcout => n1495,
            ltout => OPEN,
            carryin => n12543,
            carryout => n12544,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_9_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53611\,
            in2 => \N__50979\,
            in3 => \N__50955\,
            lcout => n1494,
            ltout => OPEN,
            carryin => n12544,
            carryout => n12545,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_10_lut_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53607\,
            in2 => \N__50952\,
            in3 => \N__50928\,
            lcout => n1493,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => n12546,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_11_lut_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53612\,
            in2 => \N__50925\,
            in3 => \N__50898\,
            lcout => n1492,
            ltout => OPEN,
            carryin => n12546,
            carryout => n12547,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_12_lut_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53608\,
            in2 => \N__51213\,
            in3 => \N__50889\,
            lcout => n1491,
            ltout => OPEN,
            carryin => n12547,
            carryout => n12548,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_13_lut_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53613\,
            in2 => \N__50886\,
            in3 => \N__50847\,
            lcout => n1490,
            ltout => OPEN,
            carryin => n12548,
            carryout => n12549,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_14_lut_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53614\,
            in1 => \N__51317\,
            in2 => \N__50844\,
            in3 => \N__50823\,
            lcout => n1521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12837_1_lut_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51393\,
            lcout => n15562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i904_3_lut_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51306\,
            in1 => \N__51683\,
            in2 => \_gnd_net_\,
            in3 => \N__51296\,
            lcout => n1424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i838_3_lut_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51168\,
            in2 => \N__51589\,
            in3 => \N__51189\,
            lcout => n1326,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i839_3_lut_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__51506\,
            in1 => \_gnd_net_\,
            in2 => \N__51180\,
            in3 => \N__51569\,
            lcout => n1327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_173_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51167\,
            in2 => \N__51719\,
            in3 => \N__51505\,
            lcout => OPEN,
            ltout => \n14482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12806_4_lut_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__52322\,
            in1 => \N__52195\,
            in2 => \N__51153\,
            in3 => \N__51609\,
            lcout => n1257,
            ltout => \n1257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i840_3_lut_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51150\,
            in2 => \N__51141\,
            in3 => \N__51668\,
            lcout => n1328,
            ltout => \n1328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_175_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51118\,
            in1 => \N__51682\,
            in2 => \N__51102\,
            in3 => \N__51091\,
            lcout => n14282,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i770_3_lut_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51762\,
            in2 => \N__52278\,
            in3 => \N__51732\,
            lcout => n1226,
            ltout => \n1226_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i837_3_lut_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__51568\,
            in1 => \_gnd_net_\,
            in2 => \N__51699\,
            in3 => \N__51696\,
            lcout => n1325,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i773_3_lut_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__51852\,
            in1 => \N__51882\,
            in2 => \N__52276\,
            in3 => \_gnd_net_\,
            lcout => n1229,
            ltout => \n1229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_174_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__51654\,
            in1 => \N__51487\,
            in2 => \N__51642\,
            in3 => \N__51639\,
            lcout => n13711,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12803_1_lut_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51567\,
            lcout => n15528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i772_3_lut_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51843\,
            in2 => \N__52277\,
            in3 => \N__51813\,
            lcout => n1228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i774_3_lut_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51920\,
            in2 => \N__51894\,
            in3 => \N__52264\,
            lcout => n1230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_2_lut_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51468\,
            in3 => \N__51432\,
            lcout => n1201,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => n12508,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_3_lut_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52894\,
            in2 => \N__51428\,
            in3 => \N__51960\,
            lcout => n1200,
            ltout => OPEN,
            carryin => n12508,
            carryout => n12509,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_4_lut_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51957\,
            in2 => \_gnd_net_\,
            in3 => \N__51927\,
            lcout => n1199,
            ltout => OPEN,
            carryin => n12509,
            carryout => n12510,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_5_lut_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52895\,
            in2 => \N__51924\,
            in3 => \N__51885\,
            lcout => n1198,
            ltout => OPEN,
            carryin => n12510,
            carryout => n12511,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_6_lut_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51881\,
            in3 => \N__51846\,
            lcout => n1197,
            ltout => OPEN,
            carryin => n12511,
            carryout => n12512,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_7_lut_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51842\,
            in3 => \N__51807\,
            lcout => n1196,
            ltout => OPEN,
            carryin => n12512,
            carryout => n12513,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_8_lut_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52897\,
            in2 => \N__51804\,
            in3 => \N__51765\,
            lcout => n1195,
            ltout => OPEN,
            carryin => n12513,
            carryout => n12514,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_9_lut_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52896\,
            in2 => \N__51761\,
            in3 => \N__51726\,
            lcout => n1194,
            ltout => OPEN,
            carryin => n12514,
            carryout => n12515,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_10_lut_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52892\,
            in2 => \N__52305\,
            in3 => \N__51723\,
            lcout => n1193,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => n12516,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_11_lut_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__52893\,
            in1 => \N__52355\,
            in2 => \N__52344\,
            in3 => \N__52326\,
            lcout => n1224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i769_3_lut_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__52304\,
            in1 => \_gnd_net_\,
            in2 => \N__52287\,
            in3 => \N__52274\,
            lcout => n1225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9618_4_lut_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__52170\,
            in1 => \N__54714\,
            in2 => \N__52161\,
            in3 => \N__54762\,
            lcout => \direction_N_342\,
            ltout => \direction_N_342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_303_i1_3_lut_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52033\,
            in2 => \N__52149\,
            in3 => \N__52136\,
            lcout => n1693,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20_3_lut_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52137\,
            in1 => \N__52119\,
            in2 => \_gnd_net_\,
            in3 => \N__52034\,
            lcout => OPEN,
            ltout => \n13661_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \direction_167_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000010"
        )
    port map (
            in0 => \N__54894\,
            in1 => \N__54990\,
            in2 => \N__52113\,
            in3 => \N__52081\,
            lcout => direction_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55811\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12764_2_lut_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54893\,
            in2 => \_gnd_net_\,
            in3 => \N__54986\,
            lcout => n5197,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_adj_58_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__54944\,
            in1 => \N__55437\,
            in2 => \N__54930\,
            in3 => \N__55115\,
            lcout => OPEN,
            ltout => \n22_adj_705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_59_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__55145\,
            in1 => \N__54911\,
            in2 => \N__51972\,
            in3 => \N__54705\,
            lcout => n24_adj_704,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_56_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55466\,
            in2 => \_gnd_net_\,
            in3 => \N__55130\,
            lcout => OPEN,
            ltout => \n6_adj_582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_57_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__55052\,
            in1 => \N__55415\,
            in2 => \N__54897\,
            in3 => \N__55067\,
            lcout => n14108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__54874\,
            in1 => \N__54834\,
            in2 => \N__54801\,
            in3 => \N__54748\,
            lcout => n24_adj_699,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_LC_16_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55100\,
            in2 => \_gnd_net_\,
            in3 => \N__55451\,
            lcout => n16_adj_707,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_163_LC_16_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55030\,
            in2 => \_gnd_net_\,
            in3 => \N__54567\,
            lcout => dti,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55827\,
            ce => \N__54582\,
            sr => \_gnd_net_\
        );

    \i12594_2_lut_LC_16_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55028\,
            in2 => \_gnd_net_\,
            in3 => \N__54565\,
            lcout => OPEN,
            ltout => \dti_N_333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_16_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101101111"
        )
    port map (
            in0 => \N__54697\,
            in1 => \N__56126\,
            in2 => \N__54642\,
            in3 => \N__54635\,
            lcout => n5169,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9550_1_lut_2_lut_LC_16_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55027\,
            in2 => \_gnd_net_\,
            in3 => \N__54564\,
            lcout => n1377,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12554_4_lut_LC_16_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000111"
        )
    port map (
            in0 => \N__55951\,
            in1 => \N__56013\,
            in2 => \N__55035\,
            in3 => \N__54566\,
            lcout => n5183,
            ltout => \n5183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3262_2_lut_LC_16_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__55038\,
            in3 => \N__55034\,
            lcout => n5235,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_3_lut_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__54974\,
            in1 => \N__54959\,
            in2 => \_gnd_net_\,
            in3 => \N__55160\,
            lcout => OPEN,
            ltout => \n20_adj_706_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__55175\,
            in1 => \N__55086\,
            in2 => \N__54999\,
            in3 => \N__54996\,
            lcout => n13187,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sweep_counter_657_658__i1_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54975\,
            in2 => \_gnd_net_\,
            in3 => \N__54963\,
            lcout => sweep_counter_0,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => n12999,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i2_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54960\,
            in2 => \_gnd_net_\,
            in3 => \N__54948\,
            lcout => sweep_counter_1,
            ltout => OPEN,
            carryin => n12999,
            carryout => n13000,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i3_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54945\,
            in2 => \_gnd_net_\,
            in3 => \N__54933\,
            lcout => sweep_counter_2,
            ltout => OPEN,
            carryin => n13000,
            carryout => n13001,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i4_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54929\,
            in2 => \_gnd_net_\,
            in3 => \N__54915\,
            lcout => sweep_counter_3,
            ltout => OPEN,
            carryin => n13001,
            carryout => n13002,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i5_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54912\,
            in2 => \_gnd_net_\,
            in3 => \N__54900\,
            lcout => sweep_counter_4,
            ltout => OPEN,
            carryin => n13002,
            carryout => n13003,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i6_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55176\,
            in2 => \_gnd_net_\,
            in3 => \N__55164\,
            lcout => sweep_counter_5,
            ltout => OPEN,
            carryin => n13003,
            carryout => n13004,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i7_LC_17_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55161\,
            in2 => \_gnd_net_\,
            in3 => \N__55149\,
            lcout => sweep_counter_6,
            ltout => OPEN,
            carryin => n13004,
            carryout => n13005,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i8_LC_17_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55146\,
            in2 => \_gnd_net_\,
            in3 => \N__55134\,
            lcout => sweep_counter_7,
            ltout => OPEN,
            carryin => n13005,
            carryout => n13006,
            clk => \N__55822\,
            ce => 'H',
            sr => \N__55400\
        );

    \sweep_counter_657_658__i9_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55131\,
            in2 => \_gnd_net_\,
            in3 => \N__55119\,
            lcout => sweep_counter_8,
            ltout => OPEN,
            carryin => \bfn_17_27_0_\,
            carryout => n13007,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i10_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55116\,
            in2 => \_gnd_net_\,
            in3 => \N__55104\,
            lcout => sweep_counter_9,
            ltout => OPEN,
            carryin => n13007,
            carryout => n13008,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i11_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55101\,
            in2 => \_gnd_net_\,
            in3 => \N__55089\,
            lcout => sweep_counter_10,
            ltout => OPEN,
            carryin => n13008,
            carryout => n13009,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i12_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55085\,
            in2 => \_gnd_net_\,
            in3 => \N__55071\,
            lcout => sweep_counter_11,
            ltout => OPEN,
            carryin => n13009,
            carryout => n13010,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i13_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55068\,
            in2 => \_gnd_net_\,
            in3 => \N__55056\,
            lcout => sweep_counter_12,
            ltout => OPEN,
            carryin => n13010,
            carryout => n13011,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i14_LC_17_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55053\,
            in2 => \_gnd_net_\,
            in3 => \N__55041\,
            lcout => sweep_counter_13,
            ltout => OPEN,
            carryin => n13011,
            carryout => n13012,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i15_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55467\,
            in2 => \_gnd_net_\,
            in3 => \N__55455\,
            lcout => sweep_counter_14,
            ltout => OPEN,
            carryin => n13012,
            carryout => n13013,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i16_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55452\,
            in2 => \_gnd_net_\,
            in3 => \N__55440\,
            lcout => sweep_counter_15,
            ltout => OPEN,
            carryin => n13013,
            carryout => n13014,
            clk => \N__55825\,
            ce => 'H',
            sr => \N__55401\
        );

    \sweep_counter_657_658__i17_LC_17_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55436\,
            in2 => \_gnd_net_\,
            in3 => \N__55422\,
            lcout => sweep_counter_16,
            ltout => OPEN,
            carryin => \bfn_17_28_0_\,
            carryout => n13015,
            clk => \N__55828\,
            ce => 'H',
            sr => \N__55403\
        );

    \sweep_counter_657_658__i18_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55416\,
            in2 => \_gnd_net_\,
            in3 => \N__55419\,
            lcout => sweep_counter_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55828\,
            ce => 'H',
            sr => \N__55403\
        );

    \dir_160_LC_17_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55335\,
            lcout => dir,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55832\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GHB_172_LC_18_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000100001"
        )
    port map (
            in0 => \N__56147\,
            in1 => \N__56036\,
            in2 => \N__55968\,
            in3 => \N__55881\,
            lcout => \GHB\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55833\,
            ce => \N__55633\,
            sr => \N__55592\
        );

    \GHA_170_LC_18_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110011000"
        )
    port map (
            in0 => \N__56148\,
            in1 => \N__56030\,
            in2 => \N__55962\,
            in3 => \N__55872\,
            lcout => \GHA\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55834\,
            ce => \N__55638\,
            sr => \N__55590\
        );

    \GLB_173_LC_19_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100111110000"
        )
    port map (
            in0 => \N__56144\,
            in1 => \N__55964\,
            in2 => \N__56046\,
            in3 => \N__55890\,
            lcout => \INLB_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55835\,
            ce => \N__55629\,
            sr => \N__55596\
        );

    \GHC_174_LC_19_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001010010"
        )
    port map (
            in0 => \N__56143\,
            in1 => \N__55963\,
            in2 => \N__56045\,
            in3 => \N__55889\,
            lcout => \GHC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55835\,
            ce => \N__55629\,
            sr => \N__55596\
        );

    \GLA_171_LC_19_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100000000011"
        )
    port map (
            in0 => \N__56146\,
            in1 => \N__56043\,
            in2 => \N__55961\,
            in3 => \N__55882\,
            lcout => \INLA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55836\,
            ce => \N__55637\,
            sr => \N__55591\
        );

    \GLC_175_LC_19_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011011110000"
        )
    port map (
            in0 => \N__56145\,
            in1 => \N__56044\,
            in2 => \N__55960\,
            in3 => \N__55883\,
            lcout => \INLC_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55836\,
            ce => \N__55637\,
            sr => \N__55591\
        );

    \i9540_2_lut_LC_20_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55557\,
            lcout => \INHB_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9541_2_lut_LC_20_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55505\,
            lcout => \INHC_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9539_2_lut_LC_20_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55512\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55488\,
            lcout => \INHA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
