// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Oct  4 21:29:19 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    input PIN_3 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    output PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    output PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    output PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    output PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    output PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    inout PIN_20 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    inout PIN_21 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    inout PIN_22 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire GND_net, VCC_net, CLK_c, LED_c, PIN_6_c_0, PIN_7_c_1, PIN_8_c_2, 
        PIN_9_c_3, PIN_10_c_4, PIN_11_c_5, PIN_13_c, PIN_18_c_1, PIN_19_c_0, 
        PIN_23_c_1, PIN_24_c_0, tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(55[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(56[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(57[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(58[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(59[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(60[22:24])
    
    wire n48398;
    wire [23:0]Kd;   // verilog/TinyFPGA_B.v(61[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(62[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(63[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(64[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(65[22:30])
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(66[22:34])
    
    wire hall1, hall2, hall3;
    wire [23:0]pwm;   // verilog/TinyFPGA_B.v(74[10:13])
    wire [31:0]motor_state;   // verilog/TinyFPGA_B.v(134[22:33])
    
    wire PIN_13_N_26;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    
    wire rx_data_ready, n47035, n47012, n47008;
    wire [31:0]motor_state_23__N_27;
    wire [24:0]displacement_23__N_93;
    wire [23:0]displacement_23__N_1;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n48905, n49122;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(95[12:26])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n249, n248, n224, n6, n123, n124;
    wire [31:0]\FRAME_MATCHER.state_31__N_1861 ;
    
    wire n4, n48271, n2, n2281, n2280, n2279, n47858, n28462, 
        n740, n4_adj_4022, n48400, n2_adj_4023, n48445, n47816, 
        n22402, n22399, n22396, n46997, n43357, n48415, n22393, 
        n47798, n22390, n46987, n26846, n22387, n22384, n22381, 
        n49118, n2_adj_4024, n24099, n24098, n22378, n47773, n47771, 
        n24097, n22375, n24096, n22372, n24095, n28925, n24094, 
        n22369, n47761, n2278, n2277, n2103, n2250, n2249, n2248, 
        n2247, n2246, n2245, n2244, n2243, n2242, n2241, n2240, 
        n2239, n2238, n47759, n2857, n47755, n36229, n36228, n47753;
    wire [31:0]\FRAME_MATCHER.state_31__N_1989 ;
    
    wire n24093, n24092, n24091, n24090, n24089, n24088, n22366, 
        n24087, n24086, n24085, n24084, n24083, n24082, n36227, 
        n36226, n22363, n47747, n48453, n47745, n24081, n24080, 
        n48670, n28961, n3761, n36225, n47737, n47735, n47731, 
        n47729, n47725, n48197, n47721, n37005, n37004, n37003, 
        n37002, n37001, n37000, n36999, n36998, n36997, n36996, 
        n36995, n47707, n48205, n36994, n36993, n36992, n48447, 
        n47703, n36991, n47701, n36990, n48451, n22360, n36989, 
        n36988, n47698, n36987, n36986, n36985, n36984, n36983, 
        n36982, n36981, n36980, n36979, n36978, n25767, n36977, 
        n36976, n36975, n36974, n36973, n36972, n36971, n36970, 
        n36969, n36968, n36967, n36966, n36965, n36964, n36963, 
        n36962, n24079, n36961, n36960, n49114, n24078, n22357, 
        n49, n24077, n24076, n42425, n47681, n42559, n42424, n24075, 
        n23930, n23929, n23928, n23927, n23926, n23925, n23924, 
        n23923, n23914, n23913, n23912, n23911, n23910, n23909, 
        n23908, n23907, n23898, n23897, n23896, n23895, n23894, 
        n23893, n23892, n23891, n23882, n23881, n23880, n23879, 
        n23878, n23877, n23876, n23875, n23866, n23865, n23864, 
        n23863, n23862, n23861, n23860, n23859, n23858, n23857, 
        n23856, n23855, n23854, n23853, n23852, n23851, n23850, 
        n23849, n23848, n23847, n23846, n23844, n23843, n23834, 
        n23833, n23832, n23831, n23830, n23828, n23827, n23818, 
        n23817, n23816, n23815, n23814, n23813, n23812, n23811, 
        n23802, n23801, n23800, n23799, n23798, n23797, n23796, 
        n23795, n6832, n48578, n99, n98, n97, n96, n95, n94, 
        n93, n92, n91, n90, n89, n88, n87, n86, n85, n84, 
        n83, n82, n81, n80, n79, n78, n77, n75, n74, n73, 
        n72, n71, n70, n69, n68, n67, n66, n65, n64, n63, 
        n62, n61, n60, n59, n58, n57, n56, n55, n54, n53, 
        n25, n24, n23, n22, n21, n20, n19, n18, n17, n16, 
        n15, n14, n13, n12, n11, n10, n9, n8, n7, n6_adj_4025, 
        n5, n4_adj_4026, n3, n23786, n23785, n23784, n23783, n23782, 
        n23781, n23780, n23779, n23770, n23769, n23768, n23767, 
        n23766, n23765, n23764, n10_adj_4027, n36176, n36175, n36174, 
        n36173, n5_adj_4028, n36172, n36171, n7021, n6996, n6972, 
        n6949, n4010, n23763, n3813, n3812, n3811, n3810, n3809, 
        n3808, n3807, n3806, n3805, n3804, n3803, n3802, n3801, 
        n3800, n3799, n3798, n3797, n3796, n3795, n3794, n3793, 
        n3792, n3791, n3790, n2237, n2236, n2235, n2234, n2233, 
        n2_adj_4029, n4_adj_4030, n22354, n22351, n48247, n15_adj_4031, 
        n15_adj_4032, n2228, n2229, n89_adj_4033, n2227;
    wire [31:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(30[23:26])
    wire [31:0]\PID_CONTROLLER.err_prev ;   // verilog/motorControl.v(31[23:31])
    
    wire n36170;
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(32[23:29])
    wire [8:0]pwm_count;   // verilog/motorControl.v(62[13:22])
    
    wire n24074, n25_adj_4034, n24_adj_4035, n23_adj_4036, n22_adj_4037, 
        n21_adj_4038, n20_adj_4039, n19_adj_4040, n18_adj_4041, n17_adj_4042, 
        n16_adj_4043, n15_adj_4044, n14_adj_4045, n13_adj_4046, n12_adj_4047, 
        n11_adj_4048, n10_adj_4049, n9_adj_4050, n8_adj_4051, n7_adj_4052, 
        n6_adj_4053, n41786;
    wire [31:0]pwm_23__N_2960;
    
    wire pwm_23__N_2957, n387, n36169, n399, n400, n406, n407, 
        n413, n415, n448, n449, n452, n453, n454, n455, n456, 
        n459, n460, n461, n462, n463, n465, n467, n468, n469, 
        n470, n471, n36168, n4_adj_4054, n4_adj_4055, n2232, n2231, 
        n2230, n853, n855, n856, n857, n859, n860, n861, n862, 
        n863, n864, n865, n866, n867, n868, n869, n870, n871, 
        n872, n873, n874, n875, n4032, n36167, n22348, n22296, 
        n15_adj_4056, n6927, quadA_debounced, quadB_debounced, count_enable, 
        n47611, n36166, n36165, n36164, n36163, n36162, n48602, 
        n36161, quadA_debounced_adj_4057, quadB_debounced_adj_4058, count_enable_adj_4059, 
        n2300, n2299, n2298, n2297, n2296, n2295, n2294, n2293, 
        n2311, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n2292, n2291, n42418, n24073, n24072, n24071, n2290, 
        n36393, n36392;
    wire [2:0]r_SM_Main_adj_4476;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_4477;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_4478;   // verilog/uart_tx.v(33[16:27])
    
    wire n2289;
    wire [2:0]r_SM_Main_2__N_2753;
    
    wire o_Tx_Serial_N_2784, n313, n314, n315, n24070, n24069, n24068, 
        n22289, n316, n317, n318, n319, n320, n2288, n2287, 
        n2286, n2285, n2284;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n2283;
    wire [1:0]reg_B_adj_4485;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n36160, n2282, n44196, n36159, n6906, n36391, n36390, 
        n3346, n20420, n36389, n36388, n24066, n48664, n3_adj_4067, 
        n36158, n36893, n47549, n48269, n369, n370, n371, n372, 
        n373, n374, n375, n376, n377, n378, n379, n380, n381, 
        n382, n383, n384, n385, n386, n387_adj_4068, n388, n389, 
        n390, n391, n392, n393, n36892, n36891, n36890, n36889, 
        n36888, n36157, n36156, n36887, n36886, n36885, n36884, 
        n36155, n36154, n36883, n510, n533, n534, n36882, n36881, 
        n36880, n36879, n36878, n36877, n36876, n36875, n36874, 
        n558, n47539, n36873, n47537, n36872, n648, n649, n36871, 
        n36870, n36869, n671, n672, n36868, n36867, n36866, n36865, 
        n36864, n36863, n6849, n36862, n36861, n36860, n36859, 
        n20435, n783, n784, n785, n806, n807, n36858, n36857, 
        n36856, n36855, n36854, n36853, n48450, n36852, n36851, 
        n36850, n36849, n914, n915, n916, n917, n918, n938, 
        n939, n36848, n36847, n1043, n1044, n1045, n1046, n1047, 
        n1048, n1067, n1068, n36846, n36845, n23547, n1169, n1170, 
        n1171, n1172, n1173, n1174, n1175, n1193, n1194, n36844, 
        n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
        n23545, n1316, n1317, n36843, n36842, n6867, n1412, n1413, 
        n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1436, 
        n1437, n36841, n42413, n36840, n36839, n1529, n1530, n1531, 
        n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1553, 
        n1554, n47495, n36838, n36837, n48622, n36836, n6737, 
        n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, 
        n6746, n6747, n1643, n1644, n1645, n1646, n1647, n1648, 
        n1649, n1650, n1651, n1652, n1653, n1667, n1668, n36835, 
        n16810, n47484, n36834, n1754, n1755, n1756, n1757, n1758, 
        n1759, n1760, n1761, n1762, n1763, n1764, n1765, n47479, 
        n1778, n1779, n36833, n36832, n36831, n36830, n1862, n1863, 
        n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, 
        n1872, n1873, n1874, n1886, n1887, n36829, n36828, n20088, 
        n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, 
        n6843, n6844, n6845, n6846, n6847, n6848, n36827, n36826, 
        n36825, n20471, n1967, n1968, n1969, n1970, n1971, n1972, 
        n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
        n36824, n36823, n1991, n1992, n36822, n36821, n36820, 
        n36819, n6852, n6853, n6854, n6855, n6856, n6857, n6858, 
        n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, 
        n36818, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
        n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
        n36817, n2093, n2094, n48287, n36816, n36815, n6870, n6871, 
        n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, 
        n6880, n6881, n6882, n6883, n6884, n6885, n36814, n36813, 
        n36812, n36811, n2168, n2169, n2170, n2171, n2172, n2173, 
        n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, 
        n2182, n2183, n5820, n2192, n2193, n36810, n36809, n36808, 
        n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, 
        n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, 
        n6905, n36807, n36806, n2264, n2265, n2266, n2267, n2268, 
        n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
        n2277_adj_4069, n2278_adj_4070, n2279_adj_4071, n2280_adj_4072, 
        n2288_adj_4073, n2289_adj_4074, n20195, n6909, n6910, n6911, 
        n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, 
        n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6212, 
        n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, 
        n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
        n2373, n2374, n36805, n2381, n2382, n36804, n6930, n6931, 
        n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, 
        n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, 
        n6948, n2447, n2448, n2449, n2450, n2451, n2452, n2453, 
        n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, 
        n2462, n2463, n2464, n2465, n2471, n2472, n36803, n36802, 
        n48291, n36801, n6952, n6953, n6954, n6955, n6956, n6957, 
        n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
        n6966, n6967, n6968, n6969, n6970, n6971, n6573, n36800, 
        n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, 
        n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, 
        n2550, n2551, n2552, n2553, n2558, n2559, n36799, n36798, 
        n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, 
        n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, 
        n6991, n6992, n6993, n6994, n6995, n5821, n36797, n2618, 
        n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
        n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, 
        n2635, n2636, n2637, n2638, n2642, n2643, n6999, n7000, 
        n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, 
        n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, 
        n7017, n7018, n7019, n7020, n2699, n2700, n2701, n2702, 
        n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
        n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
        n2719, n2720, n36796, n2723, n2724, n2777, n2798, n2799, 
        n36795, n2801, n2802, n36794, n23732, n23731, n23730, 
        n23729, n23728, n23727, n23726, n23725, n23724, n23723, 
        n23722, n23721, n23720, n23719, n23718, n23717, n23716, 
        n36793, n36792, n36791, n6213, n23715, n36790, n36789, 
        n36788, n36787, n36786, n36785, n36784, n36783, n36782, 
        n36781, n36780, n36779, n36778, n48655, n48668, n6574, 
        n36777, n36776, n36775, n36774, n36773, n36772, n36771, 
        n36770, n6644, n5822, n36769, n36768, n36767, n36766, 
        n47413, n36765, n36764, n36763, n36762, n36761, n36760, 
        n63_adj_4075, n22277, n36759, n22309, n36758, n36757, n36756, 
        n36755, n36754, n36753, n36752, n36751, n36750, n36749, 
        n36748, n36747, n36746, n36745, n36744, n6214, n36743, 
        n7_adj_4076, n36742, n48608, n36741, n36740, n36739, n36738, 
        n36737, n36736, n36735, n36734, n6575, n36733, n36732, 
        n42406, n36731, n22345, n6684, n6645, n36730, n36729, 
        n36728, n5823, n36727, n36726, n36725, n36724, n47401, 
        n36723, n36722, n36721, n36720, n6215, n47397, n36719, 
        n36718, n36717, n36716, n36715, n36714, n36713, n36712, 
        n36711, n36710, n6576, n6724, n6685, n6646, n5824, n47395, 
        n36709, n36708, n36707, n36706, n36705, n36704, n23714, 
        n46881, n11_adj_4077, n15_adj_4078, n27, n29, n41, n43, 
        n11_adj_4079, n15_adj_4080, n27_adj_4081, n29_adj_4082, n41_adj_4083, 
        n43_adj_4084, n49982, n8_adj_4085, n11_adj_4086, n15_adj_4087, 
        n27_adj_4088, n29_adj_4089, n49095, n41_adj_4090, n43_adj_4091, 
        n23713, n23712, n23711, n23710, n6831, n36703, n42405, 
        n23709, n42422, n4_adj_4092, n6_adj_4093, n8_adj_4094, n9_adj_4095, 
        n11_adj_4096, n13_adj_4097, n14_adj_4098, n15_adj_4099, n23706, 
        n23705, n23704, n23703, n23702, n23701, n23700, n23699, 
        n23698, n8_adj_4100, n23697, n6_adj_4101, n23696, n4_adj_4102, 
        n23695, n23694, n23693, n23692, n23691, n23690, n2_adj_4103, 
        n23689, n23688, n23687, n23686, n23685, n23684, n23683, 
        n23680, n36702, n23650, n23649, n23648, n23647, n23646, 
        n23645, n23644, n23643, n23640, n23637, n23634, n23630, 
        n23629, n23627, n23624, n47387, n23621, n23618, n46865, 
        n23615, n23612, n46862, n23609, n36701, n6886, n47383, 
        n47381, n36700, n6216, n48309, n6577, n36699, n36698, 
        n6778, n36697, n6725, n6686, n36696, n6647, n36695, n36694, 
        n5825, n36693, n22303, n36692, n36691, n36690, n36689, 
        n47373, n6217, n36688, n36687, n36686, n36685, n6578, 
        n36684, n36683, n36682, n6819, n6779, n6726, n36681, n48452, 
        n6687, n6648, n23013, n36680, n36679, n47368, n36678, 
        n36677, n36676, n6218, n36675, n36674, n4_adj_4104, n6_adj_4105, 
        n8_adj_4106, n9_adj_4107, n16_adj_4108, n5017, n36673, n36672, 
        n6790, n6830, n48965, n36671, n36670, n36669, n36668, 
        n47366, n6579, n6820, n6780, n36667, n6727, n6688, n6649, 
        n36666, n36665, n36664, n2_adj_4109, n3_adj_4110, n4_adj_4111, 
        n5_adj_4112, n6_adj_4113, n7_adj_4114, n8_adj_4115, n9_adj_4116, 
        n10_adj_4117, n11_adj_4118, n12_adj_4119, n13_adj_4120, n14_adj_4121, 
        n15_adj_4122, n16_adj_4123, n17_adj_4124, n18_adj_4125, n19_adj_4126, 
        n20_adj_4127, n21_adj_4128, n22_adj_4129, n23_adj_4130, n24_adj_4131, 
        n25_adj_4132, n2_adj_4133, n3_adj_4134, n4_adj_4135, n5_adj_4136, 
        n6_adj_4137, n7_adj_4138, n8_adj_4139, n9_adj_4140, n10_adj_4141, 
        n11_adj_4142, n12_adj_4143, n13_adj_4144, n14_adj_4145, n15_adj_4146, 
        n16_adj_4147, n17_adj_4148, n18_adj_4149, n19_adj_4150, n20_adj_4151, 
        n21_adj_4152, n22_adj_4153, n23_adj_4154, n24_adj_4155, n25_adj_4156, 
        n36663, n6580, n36662, n6821, n6781, n6728, n6689, n6650, 
        n36661, n36660, n36659, n36658, n36657, n47354, n36656, 
        n36655, n36654, n36653, n36652, n6822, n6782, n6729, n6690, 
        n6651, n47352, n36651, n46, n36650, n36649, n48618, n36648, 
        n36647, n6823, n48963, n6783, n6730, n44, n48223, n36646, 
        n6691, n36645, n6652, n42421, n47348, n42, n48669, n46844, 
        n6824, n6784, n6731, n6692, n47343, n40, n42_adj_4157, 
        n44_adj_4158, n45, n38, n40_adj_4159, n42_adj_4160, n43_adj_4161, 
        n48227, n48667, n24258, n24257, n24256, n24255, n24254, 
        n24253, n24252, n24251, n6825, n6785, n6732, n6693, n24250, 
        n24249, n36, n38_adj_4162, n40_adj_4163, n41_adj_4164, n48966, 
        n24248, n24247, n24246, n24245, n24244, n24243, n24242, 
        n24241, n24240, n24239, n24238, n24237, n24236, n24235, 
        n34, n36_adj_4165, n38_adj_4166, n39, n41_adj_4167, n43_adj_4168, 
        n44_adj_4169, n45_adj_4170, n24231, n24227, n24225, n24224, 
        n24221, n24220, n24219, n24218, n24217, n6826, n6786, 
        n6733, n32, n34_adj_4171, n37, n39_adj_4172, n41_adj_4173, 
        n43_adj_4174, n24214, n24213, n24212, n24211, n24210, n24208, 
        n24206, n24205, n24204, n24203, n24202, n46834, n30, n31, 
        n32_adj_4175, n33, n34_adj_4176, n35, n37_adj_4177, n39_adj_4178, 
        n48449, n41_adj_4179, n42_adj_4180, n43_adj_4181, n45_adj_4182, 
        n24201, n24200, n24199, n24198, n24197, n24196, n24195, 
        n24194, n24193, n24192, n24191, n24190, n24189, n48663, 
        n24188, n6827, n24187, n6787, n28, n29_adj_4183, n30_adj_4184, 
        n31_adj_4185, n32_adj_4186, n33_adj_4187, n35_adj_4188, n37_adj_4189, 
        n39_adj_4190, n40_adj_4191, n41_adj_4192, n43_adj_4193, n48531, 
        n48861, n24186, n24185, n6734, n24184, n24183, n24182, 
        n24181, n26, n27_adj_4194, n28_adj_4195, n29_adj_4196, n30_adj_4197, 
        n31_adj_4198, n33_adj_4199, n35_adj_4200, n37_adj_4201, n38_adj_4202, 
        n39_adj_4203, n41_adj_4204, n24172, n24171, n24170, n24_adj_4205, 
        n25_adj_4206, n26_adj_4207, n27_adj_4208, n28_adj_4209, n29_adj_4210, 
        n30_adj_4211, n31_adj_4212, n32_adj_4213, n33_adj_4214, n35_adj_4215, 
        n36_adj_4216, n37_adj_4217, n39_adj_4218, n48533, n24063, 
        n23584, n23583, n23581, n43090, n23580, n22_adj_4219, n23_adj_4220, 
        n24_adj_4221, n25_adj_4222, n26_adj_4223, n27_adj_4224, n28_adj_4225, 
        n29_adj_4226, n30_adj_4227, n31_adj_4228, n33_adj_4229, n34_adj_4230, 
        n35_adj_4231, n37_adj_4232, n39_adj_4233, n48887, n41_adj_4234, 
        n43_adj_4235, n48859, n6828, n23579, n23578, n6788, n23577, 
        n23576, n23574, n20_adj_4236, n21_adj_4237, n22_adj_4238, 
        n23_adj_4239, n24_adj_4240, n25_adj_4241, n26_adj_4242, n27_adj_4243, 
        n28_adj_4244, n29_adj_4245, n31_adj_4246, n32_adj_4247, n33_adj_4248, 
        n35_adj_4249, n37_adj_4250, n39_adj_4251, n41_adj_4252, n48543, 
        n48968, n48927, n23463, n18_adj_4253, n19_adj_4254, n20_adj_4255, 
        n21_adj_4256, n22_adj_4257, n23_adj_4258, n24_adj_4259, n25_adj_4260, 
        n26_adj_4261, n27_adj_4262, n29_adj_4263, n30_adj_4264, n31_adj_4265, 
        n33_adj_4266, n35_adj_4267, n48891, n37_adj_4268, n39_adj_4269, 
        n41_adj_4270, n43_adj_4271, n45_adj_4272, n48545, n23457, 
        n43088, n43086, n16_adj_4273, n17_adj_4274, n18_adj_4275, 
        n19_adj_4276, n20_adj_4277, n21_adj_4278, n22_adj_4279, n23_adj_4280, 
        n25_adj_4281, n27_adj_4282, n28_adj_4283, n29_adj_4284, n31_adj_4285, 
        n33_adj_4286, n48893, n35_adj_4287, n37_adj_4288, n39_adj_4289, 
        n41_adj_4290, n43_adj_4291, n14_adj_4292, n16_adj_4293, n17_adj_4294, 
        n18_adj_4295, n19_adj_4296, n20_adj_4297, n21_adj_4298, n22_adj_4299, 
        n23_adj_4300, n25_adj_4301, n26_adj_4302, n27_adj_4303, n29_adj_4304, 
        n31_adj_4305, n48705, n33_adj_4306, n35_adj_4307, n37_adj_4308, 
        n39_adj_4309, n40_adj_4310, n41_adj_4311, n43_adj_4312, n45_adj_4313, 
        n48929, n23444, n12_adj_4314, n14_adj_4315, n15_adj_4316, 
        n16_adj_4317, n17_adj_4318, n18_adj_4319, n19_adj_4320, n20_adj_4321, 
        n21_adj_4322, n23_adj_4323, n24_adj_4324, n25_adj_4325, n27_adj_4326, 
        n29_adj_4327, n31_adj_4328, n33_adj_4329, n35_adj_4330, n37_adj_4331, 
        n38_adj_4332, n39_adj_4333, n41_adj_4334, n43_adj_4335, n48855, 
        n49125, n6829, n6789, n10_adj_4336, n12_adj_4337, n13_adj_4338, 
        n14_adj_4339, n15_adj_4340, n16_adj_4341, n17_adj_4342, n18_adj_4343, 
        n19_adj_4344, n21_adj_4345, n22_adj_4346, n23_adj_4347, n25_adj_4348, 
        n27_adj_4349, n48899, n29_adj_4350, n48409, n31_adj_4351, 
        n33_adj_4352, n35_adj_4353, n36_adj_4354, n37_adj_4355, n39_adj_4356, 
        n41_adj_4357, n49119, n6748, n8_adj_4358, n10_adj_4359, n11_adj_4360, 
        n12_adj_4361, n13_adj_4362, n14_adj_4363, n15_adj_4364, n16_adj_4365, 
        n17_adj_4366, n19_adj_4367, n20_adj_4368, n21_adj_4369, n23_adj_4370, 
        n25_adj_4371, n27_adj_4372, n29_adj_4373, n31_adj_4374, n33_adj_4375, 
        n34_adj_4376, n35_adj_4377, n37_adj_4378, n39_adj_4379, n48554, 
        n48970, n48556, n6_adj_4380, n8_adj_4381, n9_adj_4382, n10_adj_4383, 
        n11_adj_4384, n12_adj_4385, n13_adj_4386, n14_adj_4387, n15_adj_4388, 
        n17_adj_4389, n19_adj_4390, n21_adj_4391, n23_adj_4392, n48560, 
        n25_adj_4393, n48654, n27_adj_4394, n29_adj_4395, n48652, 
        n31_adj_4396, n32_adj_4397, n33_adj_4398, n35_adj_4399, n37_adj_4400, 
        n48648, n4_adj_4401, n6_adj_4402, n7_adj_4403, n8_adj_4404, 
        n9_adj_4405, n10_adj_4406, n11_adj_4407, n12_adj_4408, n13_adj_4409, 
        n15_adj_4410, n16_adj_4411, n17_adj_4412, n19_adj_4413, n21_adj_4414, 
        n48646, n23_adj_4415, n24_adj_4416, n25_adj_4417, n27_adj_4418, 
        n48644, n29_adj_4419, n30_adj_4420, n31_adj_4421, n33_adj_4422, 
        n35_adj_4423, n48576, n37_adj_4424, n39_adj_4425, n40_adj_4426, 
        n41_adj_4427, n43_adj_4428, n45_adj_4429, n48932, n47323, 
        n49981, n36614, n36613, n48624, n36612, n47321, n36611, 
        n36610, n6_adj_4430, n36609, n49980, n47317, n36608, n23570, 
        n47315, n47297, n47295, n47293, n47289, n48653, n47267, 
        n47265, n47261, n47259, n48448, n48630, n10_adj_4431, n47233, 
        n47231, n47225, n47221, n43935, n48446, n38879, n22538, 
        n22908, n46798, n24067, n22424, n22283, n22422, n49816, 
        n22411, n22405, n43884, n48647, n47185, n48952, n22589, 
        n47177, n47175, n42400, n22501, n30_adj_4432, n28_adj_4433, 
        n26_adj_4434, n47169, n25_adj_4435, n21_adj_4436, n47165, 
        n1, n46779, n46764, n46762, n22416, n46748, n46744, n46742, 
        n28374, n47149, n48645, n47141, n47137, n48428, n47131, 
        n47127, n48427, n48422, n48421, n47109, n48397, n47099, 
        n47097, n47093, n48151, n47089, n5_adj_4437, n46732, n6_adj_4438, 
        n46730, n44294, n48399, n48211, n49120, n49126, n49106, 
        n49105, n49100, n46671, n46670, n49121, n49060, n49056, 
        n49044, n49042, n49041, n49034, n49099, n49097, n49039, 
        n49043, n48999, n49055, n48983, n49057, n48979, n48978, 
        n49059, n48973, n48904, n48900, n48898, n48896, n48894, 
        n48892, n48890, n48888, n48866, n48864, n48860, n49116, 
        n42428, n48964, n48772, n48771, n48962, n42633, n7_adj_4439, 
        n48883, n48728, n48727, n48885, n48720, n48889, n48714, 
        n48712, n48710, n48895, n46620, n46619, n48704, n48897, 
        n48700, n10_adj_4440, n42621, n43181, n42614, n48698, n48901, 
        n48903, n48693, n48573, n48571, n48221, n48563, n48559, 
        n46724, n42896, n48548, n48546, n46722, n48660, n42920, 
        n43032, n48527, n48525, n50261, n50258, n48119, n48923, 
        n43011, n43035, n50246, n47976, n47974, n46707, n48416, 
        n48930, n48251, n48410, n48406, n47894, n47932, n48307, 
        n47940, n47944, n48590, n48405;
    
    VCC i2 (.Y(VCC_net));
    SB_CARRY div_11_unary_minus_4_add_3_12 (.CI(n36969), .I0(GND_net), .I1(n15_adj_4122), 
            .CO(n36970));
    SB_IO hall1_input (.PACKAGE_PIN(PIN_20), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4123), .I3(n36968), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_IO hall2_input (.PACKAGE_PIN(PIN_21), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_22), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_93[21]), 
            .I2(n3_adj_4067), .I3(n36174), .O(displacement_23__N_1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY div_11_unary_minus_4_add_3_11 (.CI(n36968), .I0(GND_net), .I1(n16_adj_4123), 
            .CO(n36969));
    SB_LUT4 div_11_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4124), .I3(n36967), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    motorControl control (.GND_net(GND_net), .deadband({deadband}), .\PID_CONTROLLER.result[13] (\PID_CONTROLLER.result [13]), 
            .n459(n459), .n460(n460), .\PID_CONTROLLER.err[9] (\PID_CONTROLLER.err [9]), 
            .n461(n461), .\PID_CONTROLLER.err[8] (\PID_CONTROLLER.err [8]), 
            .\PID_CONTROLLER.err[7] (\PID_CONTROLLER.err [7]), .n462(n462), 
            .\PID_CONTROLLER.err[6] (\PID_CONTROLLER.err [6]), .n463(n463), 
            .\PID_CONTROLLER.err[5] (\PID_CONTROLLER.err [5]), .\PID_CONTROLLER.result[7] (\PID_CONTROLLER.result [7]), 
            .n465(n465), .\PID_CONTROLLER.err[4] (\PID_CONTROLLER.err [4]), 
            .\PID_CONTROLLER.err[3] (\PID_CONTROLLER.err [3]), .\PID_CONTROLLER.err[2] (\PID_CONTROLLER.err [2]), 
            .\PID_CONTROLLER.err[1] (\PID_CONTROLLER.err [1]), .\PID_CONTROLLER.err[0] (\PID_CONTROLLER.err [0]), 
            .pwm_count({pwm_count}), .\pwm_23__N_2960[13] (pwm_23__N_2960[13]), 
            .VCC_net(VCC_net), .\PID_CONTROLLER.result[5] (\PID_CONTROLLER.result [5]), 
            .\pwm_23__N_2960[14] (pwm_23__N_2960[14]), .\PID_CONTROLLER.result[14] (\PID_CONTROLLER.result [14]), 
            .n467(n467), .n468(n468), .n469(n469), .n470(n470), .n50246(n50246), 
            .\PID_CONTROLLER.result[21] (\PID_CONTROLLER.result [21]), .\pwm_23__N_2960[20] (pwm_23__N_2960[20]), 
            .\PID_CONTROLLER.result[20] (\PID_CONTROLLER.result [20]), .n27(n27), 
            .n29(n29), .n471(n471), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .\motor_state[18] (motor_state[18]), .\motor_state[17] (motor_state[17]), 
            .n41(n41), .pwm_23__N_2957(pwm_23__N_2957), .\motor_state[16] (motor_state[16]), 
            .n399(n399), .n24225(n24225), .pwm({pwm}), .clk32MHz(clk32MHz), 
            .n24224(n24224), .n24221(n24221), .n24220(n24220), .n24219(n24219), 
            .n24218(n24218), .n24217(n24217), .n24214(n24214), .n24213(n24213), 
            .n24212(n24212), .n24211(n24211), .n24210(n24210), .n24208(n24208), 
            .n24206(n24206), .n24205(n24205), .n24204(n24204), .n24203(n24203), 
            .n24172(n24172), .n400(n400), .\motor_state[15] (motor_state[15]), 
            .PIN_7_c_1(PIN_7_c_1), .\motor_state[14] (motor_state[14]), 
            .PIN_6_c_0(PIN_6_c_0), .\motor_state[13] (motor_state[13]), 
            .\motor_state[12] (motor_state[12]), .\motor_state[11] (motor_state[11]), 
            .\motor_state[10] (motor_state[10]), .\motor_state[9] (motor_state[9]), 
            .\motor_state[8] (motor_state[8]), .\motor_state[7] (motor_state[7]), 
            .\motor_state[6] (motor_state[6]), .\motor_state[5] (motor_state[5]), 
            .\motor_state[4] (motor_state[4]), .\motor_state[3] (motor_state[3]), 
            .\motor_state[2] (motor_state[2]), .n406(n406), .\motor_state[1] (motor_state[1]), 
            .n407(n407), .\motor_state[0] (motor_state[0]), .\PID_CONTROLLER.err_prev[31] (\PID_CONTROLLER.err_prev [31]), 
            .\PID_CONTROLLER.err_prev[23] (\PID_CONTROLLER.err_prev [23]), 
            .\PID_CONTROLLER.err_prev[22] (\PID_CONTROLLER.err_prev [22]), 
            .\PID_CONTROLLER.err_prev[21] (\PID_CONTROLLER.err_prev [21]), 
            .\PID_CONTROLLER.err_prev[20] (\PID_CONTROLLER.err_prev [20]), 
            .\PID_CONTROLLER.err_prev[19] (\PID_CONTROLLER.err_prev [19]), 
            .\PID_CONTROLLER.err_prev[18] (\PID_CONTROLLER.err_prev [18]), 
            .\PID_CONTROLLER.err_prev[17] (\PID_CONTROLLER.err_prev [17]), 
            .\PID_CONTROLLER.err_prev[16] (\PID_CONTROLLER.err_prev [16]), 
            .n413(n413), .\PID_CONTROLLER.err_prev[15] (\PID_CONTROLLER.err_prev [15]), 
            .\PID_CONTROLLER.err_prev[14] (\PID_CONTROLLER.err_prev [14]), 
            .\PID_CONTROLLER.err_prev[13] (\PID_CONTROLLER.err_prev [13]), 
            .\PID_CONTROLLER.err_prev[12] (\PID_CONTROLLER.err_prev [12]), 
            .\PID_CONTROLLER.err_prev[11] (\PID_CONTROLLER.err_prev [11]), 
            .\Kd[4] (Kd[4]), .\Kp[7] (Kp[7]), .\PID_CONTROLLER.err[17] (\PID_CONTROLLER.err [17]), 
            .n415(n415), .\PID_CONTROLLER.err_prev[10] (\PID_CONTROLLER.err_prev [10]), 
            .\PID_CONTROLLER.err_prev[9] (\PID_CONTROLLER.err_prev [9]), .\PID_CONTROLLER.err_prev[8] (\PID_CONTROLLER.err_prev [8]), 
            .\PID_CONTROLLER.err_prev[7] (\PID_CONTROLLER.err_prev [7]), .\PID_CONTROLLER.err[31] (\PID_CONTROLLER.err [31]), 
            .\PID_CONTROLLER.err_prev[6] (\PID_CONTROLLER.err_prev [6]), .\Kp[1] (Kp[1]), 
            .\PID_CONTROLLER.err[20] (\PID_CONTROLLER.err [20]), .\Kp[0] (Kp[0]), 
            .\PID_CONTROLLER.err[21] (\PID_CONTROLLER.err [21]), .\PID_CONTROLLER.err_prev[5] (\PID_CONTROLLER.err_prev [5]), 
            .\Kd[0] (Kd[0]), .\Kd[1] (Kd[1]), .\Kd[2] (Kd[2]), .\PID_CONTROLLER.err_prev[4] (\PID_CONTROLLER.err_prev [4]), 
            .\PID_CONTROLLER.err_prev[3] (\PID_CONTROLLER.err_prev [3]), .\Kp[2] (Kp[2]), 
            .\Kd[5] (Kd[5]), .\Kp[3] (Kp[3]), .hall1(hall1), .hall2(hall2), 
            .\Kp[4] (Kp[4]), .\PID_CONTROLLER.err[10] (\PID_CONTROLLER.err [10]), 
            .\Kp[5] (Kp[5]), .\PID_CONTROLLER.err_prev[2] (\PID_CONTROLLER.err_prev [2]), 
            .\PID_CONTROLLER.err_prev[1] (\PID_CONTROLLER.err_prev [1]), .\PID_CONTROLLER.err_prev[0] (\PID_CONTROLLER.err_prev [0]), 
            .\Kp[6] (Kp[6]), .\PID_CONTROLLER.err[11] (\PID_CONTROLLER.err [11]), 
            .n853(n853), .n21(n21_adj_4436), .n855(n855), .n856(n856), 
            .n857(n857), .n859(n859), .n860(n860), .n861(n861), .n862(n862), 
            .n863(n863), .n864(n864), .n865(n865), .n866(n866), .\PID_CONTROLLER.err[12] (\PID_CONTROLLER.err [12]), 
            .PWMLimit({PWMLimit}), .setpoint({setpoint}), .\Kd[6] (Kd[6]), 
            .\PID_CONTROLLER.err[16] (\PID_CONTROLLER.err [16]), .n867(n867), 
            .\PID_CONTROLLER.err[13] (\PID_CONTROLLER.err [13]), .n868(n868), 
            .n869(n869), .\Ki[3] (Ki[3]), .\Kd[7] (Kd[7]), .\Ki[7] (Ki[7]), 
            .\Kd[3] (Kd[3]), .n870(n870), .n871(n871), .n872(n872), 
            .n873(n873), .n874(n874), .n875(n875), .\PID_CONTROLLER.err[15] (\PID_CONTROLLER.err [15]), 
            .n46619(n46619), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\PID_CONTROLLER.err[14] (\PID_CONTROLLER.err [14]), .\Ki[1] (Ki[1]), 
            .\Ki[0] (Ki[0]), .\PID_CONTROLLER.err[18] (\PID_CONTROLLER.err [18]), 
            .\PID_CONTROLLER.err[19] (\PID_CONTROLLER.err [19]), .\Ki[2] (Ki[2]), 
            .\PID_CONTROLLER.err[22] (\PID_CONTROLLER.err [22]), .n448(n448), 
            .n449(n449), .\PID_CONTROLLER.err[23] (\PID_CONTROLLER.err [23]), 
            .n23732(n23732), .n23731(n23731), .n23730(n23730), .n23729(n23729), 
            .n23728(n23728), .n23727(n23727), .n23726(n23726), .n23725(n23725), 
            .n23724(n23724), .n23723(n23723), .n23722(n23722), .n23721(n23721), 
            .n23720(n23720), .n23719(n23719), .n23718(n23718), .n23717(n23717), 
            .n23716(n23716), .n23715(n23715), .n23714(n23714), .n23713(n23713), 
            .n23712(n23712), .n23711(n23711), .n23710(n23710), .n23709(n23709), 
            .n452(n452), .PIN_8_c_2(PIN_8_c_2), .PIN_9_c_3(PIN_9_c_3), 
            .PIN_10_c_4(PIN_10_c_4), .PIN_11_c_5(PIN_11_c_5), .n453(n453), 
            .n454(n454), .n455(n455), .n456(n456), .n23574(n23574), 
            .hall3(hall3), .n48211(n48211), .n25(n25_adj_4435), .n30(n30_adj_4432), 
            .n26(n26_adj_4434), .n27_adj_13(n27_adj_4088), .n15(n15_adj_4087), 
            .n11(n11_adj_4086), .n29_adj_14(n29_adj_4089), .n43(n43_adj_4091), 
            .n41_adj_15(n41_adj_4090), .n387(n387), .n27_adj_16(n27_adj_4081), 
            .n15_adj_17(n15_adj_4080), .n11_adj_18(n11_adj_4079), .n29_adj_19(n29_adj_4082), 
            .n43_adj_20(n43_adj_4084), .n41_adj_21(n41_adj_4083), .n43_adj_22(n43), 
            .n50261(n50261), .n16(n16_adj_4108), .n50258(n50258), .n15_adj_23(n15_adj_4078), 
            .n11_adj_24(n11_adj_4077), .n43357(n43357), .IntegralLimit({IntegralLimit})) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(143[16] 159[4])
    SB_CARRY div_11_unary_minus_4_add_3_10 (.CI(n36967), .I0(GND_net), .I1(n17_adj_4124), 
            .CO(n36968));
    SB_LUT4 div_11_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4125), .I3(n36966), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_10_pad (.PACKAGE_PIN(PIN_10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_10_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_10_pad.PIN_TYPE = 6'b011001;
    defparam PIN_10_pad.PULLUP = 1'b0;
    defparam PIN_10_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY div_11_unary_minus_4_add_3_9 (.CI(n36966), .I0(GND_net), .I1(n18_adj_4125), 
            .CO(n36967));
    SB_LUT4 div_11_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4126), .I3(n36965), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_8 (.CI(n36965), .I0(GND_net), .I1(n19_adj_4126), 
            .CO(n36966));
    SB_LUT4 add_2996_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n36746), 
            .O(n6876)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_12 (.CI(n36746), .I0(n2174), .I1(n90), .CO(n36747));
    SB_LUT4 add_2996_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n36745), 
            .O(n6877)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n36174), .I0(displacement_23__N_93[21]), 
            .I1(n3_adj_4067), .CO(n36175));
    SB_LUT4 div_11_i1597_3_lut_3_lut (.I0(n2381), .I1(n6923), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4127), .I3(n36964), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_11 (.CI(n36745), .I0(n2175), .I1(n91), .CO(n36746));
    SB_LUT4 i33143_3_lut (.I0(n48896), .I1(n89), .I2(n33_adj_4306), .I3(GND_net), 
            .O(n48704));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33143_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_93[20]), 
            .I2(n3_adj_4067), .I3(n36173), .O(displacement_23__N_1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33047_4_lut (.I0(n43_adj_4312), .I1(n41_adj_4311), .I2(n39_adj_4309), 
            .I3(n47177), .O(n48608));
    defparam i33047_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2996_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n36744), 
            .O(n6878)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1598_3_lut_3_lut (.I0(n2381), .I1(n6924), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_11_unary_minus_4_add_3_7 (.CI(n36964), .I0(GND_net), .I1(n20_adj_4127), 
            .CO(n36965));
    SB_LUT4 i33366_4_lut (.I0(n47747), .I1(n48548), .I2(n45_adj_4313), 
            .I3(n47169), .O(n48927));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33366_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_11_i1594_3_lut_3_lut (.I0(n2381), .I1(n6920), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2996_10 (.CI(n36744), .I0(n2176), .I1(n92), .CO(n36745));
    SB_LUT4 div_11_i1593_3_lut_3_lut (.I0(n2381), .I1(n6919), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2996_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n36743), 
            .O(n6879)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4128), .I3(n36963), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n36173), .I0(displacement_23__N_93[20]), 
            .I1(n3_adj_4067), .CO(n36174));
    SB_CARRY div_11_unary_minus_4_add_3_6 (.CI(n36963), .I0(GND_net), .I1(n21_adj_4128), 
            .CO(n36964));
    SB_CARRY add_2996_9 (.CI(n36743), .I0(n2177), .I1(n93), .CO(n36744));
    SB_LUT4 div_11_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4129), .I3(n36962), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_93[19]), 
            .I2(n6_adj_4053), .I3(n36172), .O(displacement_23__N_1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_5 (.CI(n36962), .I0(GND_net), .I1(n22_adj_4129), 
            .CO(n36963));
    SB_LUT4 div_11_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4130), .I3(n36961), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1592_3_lut_3_lut (.I0(n2381), .I1(n6918), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32184_3_lut (.I0(n48704), .I1(n88), .I2(n35_adj_4307), .I3(GND_net), 
            .O(n47745));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32184_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_11_unary_minus_4_add_3_4 (.CI(n36961), .I0(GND_net), .I1(n23_adj_4130), 
            .CO(n36962));
    SB_LUT4 add_2996_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n36742), 
            .O(n6880)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n36172), .I0(displacement_23__N_93[19]), 
            .I1(n6_adj_4053), .CO(n36173));
    SB_CARRY add_2996_8 (.CI(n36742), .I0(n2178), .I1(n94), .CO(n36743));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_93[18]), 
            .I2(n7_adj_4052), .I3(n36171), .O(displacement_23__N_1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n36741), 
            .O(n6881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4131), .I3(n36960), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_7 (.CI(n36741), .I0(n2179), .I1(n95), .CO(n36742));
    SB_CARRY div_11_unary_minus_4_add_3_3 (.CI(n36960), .I0(GND_net), .I1(n24_adj_4131), 
            .CO(n36961));
    SB_LUT4 add_2996_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n36740), 
            .O(n6882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4132), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_6 (.CI(n36740), .I0(n2180), .I1(n96), .CO(n36741));
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n36171), .I0(displacement_23__N_93[18]), 
            .I1(n7_adj_4052), .CO(n36172));
    SB_LUT4 i33368_4_lut (.I0(n47745), .I1(n48927), .I2(n45_adj_4313), 
            .I3(n48608), .O(n48929));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33368_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut (.I0(n48929), .I1(n22396), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 add_2996_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n36739), 
            .O(n6883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_5 (.CI(n36739), .I0(n2181), .I1(n97), .CO(n36740));
    SB_CARRY div_11_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4132), 
            .CO(n36960));
    SB_LUT4 add_2996_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n36738), 
            .O(n6884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_93[17]), 
            .I2(n8_adj_4051), .I3(n36170), .O(displacement_23__N_1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_4 (.CI(n36738), .I0(n2182), .I1(n98), .CO(n36739));
    SB_LUT4 div_11_i1591_3_lut_3_lut (.I0(n2381), .I1(n6917), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n36170), .I0(displacement_23__N_93[17]), 
            .I1(n8_adj_4051), .CO(n36171));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_93[16]), 
            .I2(n9_adj_4050), .I3(n36169), .O(displacement_23__N_1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32964_3_lut (.I0(n34_adj_4171), .I1(n96), .I2(n37), .I3(GND_net), 
            .O(n48525));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32964_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2996_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n36737), 
            .O(n6885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_3 (.CI(n36737), .I0(n2183), .I1(n99), .CO(n36738));
    SB_LUT4 add_2996_2_lut (.I0(GND_net), .I1(n384), .I2(n558), .I3(VCC_net), 
            .O(n6886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_2 (.CI(VCC_net), .I0(n384), .I1(n558), .CO(n36737));
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n36169), .I0(displacement_23__N_93[16]), 
            .I1(n9_adj_4050), .CO(n36170));
    SB_LUT4 add_2995_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n36736), 
            .O(n6852)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2995_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n36735), 
            .O(n6853)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_16 (.CI(n36735), .I0(n2070), .I1(n86), .CO(n36736));
    SB_LUT4 add_2995_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n36734), 
            .O(n6854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_15 (.CI(n36734), .I0(n2071), .I1(n87), .CO(n36735));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_93[15]), 
            .I2(n10_adj_4049), .I3(n36168), .O(displacement_23__N_1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2995_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n36733), 
            .O(n6855)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n36168), .I0(displacement_23__N_93[15]), 
            .I1(n10_adj_4049), .CO(n36169));
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_93[14]), 
            .I2(n11_adj_4048), .I3(n36167), .O(displacement_23__N_1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n36167), .I0(displacement_23__N_93[14]), 
            .I1(n11_adj_4048), .CO(n36168));
    SB_CARRY add_2995_14 (.CI(n36733), .I0(n2072), .I1(n88), .CO(n36734));
    SB_LUT4 add_2995_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n36732), 
            .O(n6856)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_93[13]), 
            .I2(n12_adj_4047), .I3(n36166), .O(displacement_23__N_1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n36166), .I0(displacement_23__N_93[13]), 
            .I1(n12_adj_4047), .CO(n36167));
    SB_LUT4 div_11_i1590_3_lut_3_lut (.I0(n2381), .I1(n6916), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1596_3_lut_3_lut (.I0(n2381), .I1(n6922), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4288));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1399 (.I0(n48227), .I1(n22366), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1399.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1589_3_lut_3_lut (.I0(n2381), .I1(n6915), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4291));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2995_13 (.CI(n36732), .I0(n2073), .I1(n89), .CO(n36733));
    SB_LUT4 add_2995_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n36731), 
            .O(n6857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_12 (.CI(n36731), .I0(n2074), .I1(n90), .CO(n36732));
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_93[12]), 
            .I2(n13_adj_4046), .I3(n36165), .O(displacement_23__N_1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2995_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n36730), 
            .O(n6858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_11 (.CI(n36730), .I0(n2075), .I1(n91), .CO(n36731));
    SB_LUT4 add_2995_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n36729), 
            .O(n6859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n36165), .I0(displacement_23__N_93[12]), 
            .I1(n13_adj_4046), .CO(n36166));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_93[11]), 
            .I2(n14_adj_4045), .I3(n36164), .O(displacement_23__N_1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_10 (.CI(n36729), .I0(n2076), .I1(n92), .CO(n36730));
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n36164), .I0(displacement_23__N_93[11]), 
            .I1(n14_adj_4045), .CO(n36165));
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_93[10]), 
            .I2(n15_adj_4044), .I3(n36163), .O(displacement_23__N_1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4290));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2995_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n36728), 
            .O(n6860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_9 (.CI(n36728), .I0(n2077), .I1(n93), .CO(n36729));
    SB_LUT4 add_2995_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n36727), 
            .O(n6861)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n36163), .I0(displacement_23__N_93[10]), 
            .I1(n15_adj_4044), .CO(n36164));
    SB_CARRY add_2995_8 (.CI(n36727), .I0(n2078), .I1(n94), .CO(n36728));
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_93[9]), 
            .I2(n16_adj_4043), .I3(n36162), .O(displacement_23__N_1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2995_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n36726), 
            .O(n6862)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_7 (.CI(n36726), .I0(n2079), .I1(n95), .CO(n36727));
    SB_LUT4 add_2995_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n36725), 
            .O(n6863)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n36162), .I0(displacement_23__N_93[9]), 
            .I1(n16_adj_4043), .CO(n36163));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_93[8]), 
            .I2(n17_adj_4042), .I3(n36161), .O(displacement_23__N_1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_6 (.CI(n36725), .I0(n2080), .I1(n96), .CO(n36726));
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n36161), .I0(displacement_23__N_93[8]), 
            .I1(n17_adj_4042), .CO(n36162));
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_93[7]), 
            .I2(n18_adj_4041), .I3(n36160), .O(displacement_23__N_1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1600_3_lut_3_lut (.I0(n2381), .I1(n6926), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1599_3_lut_3_lut (.I0(n2381), .I1(n6925), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2995_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n36724), 
            .O(n6864)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_5 (.CI(n36724), .I0(n2081), .I1(n97), .CO(n36725));
    SB_LUT4 add_2995_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n36723), 
            .O(n6865)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n36160), .I0(displacement_23__N_93[7]), 
            .I1(n18_adj_4041), .CO(n36161));
    SB_CARRY add_2995_4 (.CI(n36723), .I0(n2082), .I1(n98), .CO(n36724));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_93[6]), 
            .I2(n19_adj_4040), .I3(n36159), .O(displacement_23__N_1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4289));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2995_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n36722), 
            .O(n6866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_3 (.CI(n36722), .I0(n2083), .I1(n99), .CO(n36723));
    SB_LUT4 add_2995_2_lut (.I0(GND_net), .I1(n383), .I2(n558), .I3(VCC_net), 
            .O(n6867)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2995_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n36159), .I0(displacement_23__N_93[6]), 
            .I1(n19_adj_4040), .CO(n36160));
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_93[5]), 
            .I2(n20_adj_4039), .I3(n36158), .O(displacement_23__N_1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2995_2 (.CI(VCC_net), .I0(n383), .I1(n558), .CO(n36722));
    SB_LUT4 div_11_i1659_3_lut_3_lut (.I0(n2471), .I1(n6947), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n36158), .I0(displacement_23__N_93[5]), 
            .I1(n20_adj_4039), .CO(n36159));
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_93[4]), 
            .I2(n21_adj_4038), .I3(n36157), .O(displacement_23__N_1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2994_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n36721), 
            .O(n6835)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2994_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n36720), 
            .O(n6836)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_15 (.CI(n36720), .I0(n1968), .I1(n87), .CO(n36721));
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n36157), .I0(displacement_23__N_93[4]), 
            .I1(n21_adj_4038), .CO(n36158));
    SB_LUT4 add_2994_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n36719), 
            .O(n6837)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_93[3]), 
            .I2(n22_adj_4037), .I3(n36156), .O(displacement_23__N_1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_14 (.CI(n36719), .I0(n1969), .I1(n88), .CO(n36720));
    SB_LUT4 add_2994_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n36718), 
            .O(n6838)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_13 (.CI(n36718), .I0(n1970), .I1(n89), .CO(n36719));
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n36156), .I0(displacement_23__N_93[3]), 
            .I1(n22_adj_4037), .CO(n36157));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_93[2]), 
            .I2(n23_adj_4036), .I3(n36155), .O(displacement_23__N_1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n385));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1642_3_lut_3_lut (.I0(n2471), .I1(n6930), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1643_3_lut_3_lut (.I0(n2471), .I1(n6931), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1644_3_lut_3_lut (.I0(n2471), .I1(n6932), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n36155), .I0(displacement_23__N_93[2]), 
            .I1(n23_adj_4036), .CO(n36156));
    SB_LUT4 div_11_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4285));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4286));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2994_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n36717), 
            .O(n6839)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_12 (.CI(n36717), .I0(n1971), .I1(n90), .CO(n36718));
    SB_LUT4 add_2994_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n36716), 
            .O(n6840)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_93[1]), 
            .I2(n24_adj_4035), .I3(n36154), .O(displacement_23__N_1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_11 (.CI(n36716), .I0(n1972), .I1(n91), .CO(n36717));
    SB_LUT4 add_2994_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n36715), 
            .O(n6841)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_10 (.CI(n36715), .I0(n1973), .I1(n92), .CO(n36716));
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n36154), .I0(displacement_23__N_93[1]), 
            .I1(n24_adj_4035), .CO(n36155));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_93[0]), 
            .I2(n25_adj_4034), .I3(VCC_net), .O(displacement_23__N_1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2994_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n36714), 
            .O(n6842)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_93[0]), 
            .I1(n25_adj_4034), .CO(n36154));
    SB_CARRY add_2994_9 (.CI(n36714), .I0(n1974), .I1(n93), .CO(n36715));
    SB_LUT4 add_2994_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n36713), 
            .O(n6843)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_8 (.CI(n36713), .I0(n1975), .I1(n94), .CO(n36714));
    SB_LUT4 add_2994_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n36712), 
            .O(n6844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_7 (.CI(n36712), .I0(n1976), .I1(n95), .CO(n36713));
    SB_LUT4 add_2994_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n36711), 
            .O(n6845)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_6 (.CI(n36711), .I0(n1977), .I1(n96), .CO(n36712));
    SB_LUT4 add_2994_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n36710), 
            .O(n6846)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_5 (.CI(n36710), .I0(n1978), .I1(n97), .CO(n36711));
    SB_LUT4 add_2994_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n36709), 
            .O(n6847)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_4 (.CI(n36709), .I0(n1979), .I1(n98), .CO(n36710));
    SB_LUT4 add_2969_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n36393), 
            .O(n6212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2969_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2969_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n36392), 
            .O(n6213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2969_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2994_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n36708), 
            .O(n6848)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2969_7 (.CI(n36392), .I0(n1044), .I1(n95), .CO(n36393));
    SB_LUT4 add_2969_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n36391), 
            .O(n6214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2969_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_3 (.CI(n36708), .I0(n1980), .I1(n99), .CO(n36709));
    SB_CARRY add_2969_6 (.CI(n36391), .I0(n1045), .I1(n96), .CO(n36392));
    SB_LUT4 add_2994_2_lut (.I0(GND_net), .I1(n382), .I2(n558), .I3(VCC_net), 
            .O(n6849)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2994_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4287));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2969_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n36390), 
            .O(n6215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2969_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2994_2 (.CI(VCC_net), .I0(n382), .I1(n558), .CO(n36708));
    SB_CARRY add_2969_5 (.CI(n36390), .I0(n1046), .I1(n97), .CO(n36391));
    SB_LUT4 add_2969_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n36389), 
            .O(n6216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2969_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n36707), 
            .O(n6819)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2969_4 (.CI(n36389), .I0(n1047), .I1(n98), .CO(n36390));
    SB_LUT4 add_2969_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n36388), 
            .O(n6217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2969_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n36706), 
            .O(n6820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2969_3 (.CI(n36388), .I0(n1048), .I1(n99), .CO(n36389));
    SB_CARRY add_2993_14 (.CI(n36706), .I0(n1863), .I1(n88), .CO(n36707));
    SB_LUT4 add_2969_2_lut (.I0(GND_net), .I1(n374), .I2(n558), .I3(VCC_net), 
            .O(n6218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2969_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2993_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n36705), 
            .O(n6821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2969_2 (.CI(VCC_net), .I0(n374), .I1(n558), .CO(n36388));
    SB_CARRY add_2993_13 (.CI(n36705), .I0(n1864), .I1(n89), .CO(n36706));
    SB_LUT4 div_11_i1647_3_lut_3_lut (.I0(n2471), .I1(n6935), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2993_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n36704), 
            .O(n6822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_12 (.CI(n36704), .I0(n1865), .I1(n90), .CO(n36705));
    SB_LUT4 add_2993_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n36703), 
            .O(n6823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1645_3_lut_3_lut (.I0(n2471), .I1(n6933), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1648_3_lut_3_lut (.I0(n2471), .I1(n6936), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1661_3_lut_3_lut (.I0(n2471), .I1(n6949), .I2(n387_adj_4068), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4282));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4284));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i19_2_lut (.I0(n2278_adj_4070), .I1(n97), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4276));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i21_2_lut (.I0(n2277_adj_4069), .I1(n96), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4278));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4280));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4281));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1484_1_lut (.I0(n2288_adj_4073), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289_adj_4074));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_1482_i17_2_lut (.I0(n2279_adj_4071), .I1(n98), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4274));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1646_3_lut_3_lut (.I0(n2471), .I1(n6934), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i807_3_lut (.I0(n1174), .I1(n6578), .I2(n1193), .I3(GND_net), 
            .O(n1297));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1650_3_lut_3_lut (.I0(n2471), .I1(n6938), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31672_4_lut (.I0(n23_adj_4280), .I1(n21_adj_4278), .I2(n19_adj_4276), 
            .I3(n17_adj_4274), .O(n47233));
    defparam i31672_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_i1651_3_lut_3_lut (.I0(n2471), .I1(n6939), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31664_4_lut (.I0(n29_adj_4284), .I1(n27_adj_4282), .I2(n25_adj_4281), 
            .I3(n47233), .O(n47225));
    defparam i31664_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33057_4_lut (.I0(n35_adj_4287), .I1(n33_adj_4286), .I2(n31_adj_4285), 
            .I3(n47225), .O(n48618));
    defparam i33057_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_11_LessThan_1482_i16_4_lut (.I0(n385), .I1(n99), .I2(n2280_adj_4072), 
            .I3(n558), .O(n16_adj_4273));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32860_3_lut (.I0(n16_adj_4273), .I1(n87), .I2(n39_adj_4289), 
            .I3(GND_net), .O(n48421));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32860_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1660_3_lut_3_lut (.I0(n2471), .I1(n6948), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32861_3_lut (.I0(n48421), .I1(n86), .I2(n41_adj_4290), .I3(GND_net), 
            .O(n48422));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32861_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32379_4_lut (.I0(n41_adj_4290), .I1(n39_adj_4289), .I2(n27_adj_4282), 
            .I3(n47231), .O(n47940));
    defparam i32379_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_11_i1655_3_lut_3_lut (.I0(n2471), .I1(n6943), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32985_3_lut (.I0(n22_adj_4279), .I1(n93), .I2(n27_adj_4282), 
            .I3(GND_net), .O(n48546));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32985_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32176_3_lut (.I0(n48422), .I1(n85), .I2(n43_adj_4291), .I3(GND_net), 
            .O(n47737));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32176_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1649_3_lut_3_lut (.I0(n2471), .I1(n6937), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1653_3_lut_3_lut (.I0(n2471), .I1(n6941), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1482_i28_3_lut (.I0(n20_adj_4277), .I1(n91), 
            .I2(n31_adj_4285), .I3(GND_net), .O(n28_adj_4283));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33332_4_lut (.I0(n28_adj_4283), .I1(n18_adj_4275), .I2(n31_adj_4285), 
            .I3(n47221), .O(n48893));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33332_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_11_i1654_3_lut_3_lut (.I0(n2471), .I1(n6942), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1652_3_lut_3_lut (.I0(n2471), .I1(n6940), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33333_3_lut (.I0(n48893), .I1(n90), .I2(n33_adj_4286), .I3(GND_net), 
            .O(n48894));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33333_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1658_3_lut_3_lut (.I0(n2471), .I1(n6946), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33149_3_lut (.I0(n48894), .I1(n89), .I2(n35_adj_4287), .I3(GND_net), 
            .O(n48710));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33149_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32383_4_lut (.I0(n41_adj_4290), .I1(n39_adj_4289), .I2(n37_adj_4288), 
            .I3(n48618), .O(n47944));
    defparam i32383_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_2993_11 (.CI(n36703), .I0(n1866), .I1(n91), .CO(n36704));
    SB_LUT4 i33144_4_lut (.I0(n47737), .I1(n48546), .I2(n43_adj_4291), 
            .I3(n47940), .O(n48705));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33144_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_11_i1657_3_lut_3_lut (.I0(n2471), .I1(n6945), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32174_3_lut (.I0(n48710), .I1(n88), .I2(n37_adj_4288), .I3(GND_net), 
            .O(n47735));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32174_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1656_3_lut_3_lut (.I0(n2471), .I1(n6944), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33417_4_lut (.I0(n47735), .I1(n48705), .I2(n43_adj_4291), 
            .I3(n47944), .O(n48978));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33417_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33418_3_lut (.I0(n48978), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n48979));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33418_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_11_i1713_3_lut_3_lut (.I0(n2558), .I1(n6966), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1400 (.I0(n48979), .I1(n22393), .I2(n83), .I3(n2264), 
            .O(n2288_adj_4073));
    defparam i1_4_lut_adj_1400.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_906_i32_4_lut (.I0(n377), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_i1699_3_lut_3_lut (.I0(n2558), .I1(n6952), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32890_3_lut (.I0(n32), .I1(n95), .I2(n39_adj_4172), .I3(GND_net), 
            .O(n48451));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32890_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1700_3_lut_3_lut (.I0(n2558), .I1(n6953), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1701_3_lut_3_lut (.I0(n2558), .I1(n6954), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1702_3_lut_3_lut (.I0(n2558), .I1(n6955), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2993_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n36702), 
            .O(n6824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_10 (.CI(n36702), .I0(n1867), .I1(n92), .CO(n36703));
    SB_LUT4 add_2993_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n36701), 
            .O(n6825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_9_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_18_pad (.PACKAGE_PIN(PIN_18), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_18_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_18_pad.PIN_TYPE = 6'b000001;
    defparam PIN_18_pad.PULLUP = 1'b0;
    defparam PIN_18_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_i1705_3_lut_3_lut (.I0(n2558), .I1(n6958), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32891_3_lut (.I0(n48451), .I1(n94), .I2(n41_adj_4173), .I3(GND_net), 
            .O(n48452));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32891_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2993_9 (.CI(n36701), .I0(n1868), .I1(n93), .CO(n36702));
    SB_LUT4 add_2993_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n36700), 
            .O(n6826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32137_3_lut (.I0(n48452), .I1(n93), .I2(n43_adj_4174), .I3(GND_net), 
            .O(n47698));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32137_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2993_8 (.CI(n36700), .I0(n1869), .I1(n94), .CO(n36701));
    SB_LUT4 add_2993_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n36699), 
            .O(n6827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1703_3_lut_3_lut (.I0(n2558), .I1(n6956), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2993_7 (.CI(n36699), .I0(n1870), .I1(n95), .CO(n36700));
    SB_LUT4 add_2993_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n36698), 
            .O(n6828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4269));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2993_6 (.CI(n36698), .I0(n1871), .I1(n96), .CO(n36699));
    SB_LUT4 div_11_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4272));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2993_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n36697), 
            .O(n6829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_5 (.CI(n36697), .I0(n1872), .I1(n97), .CO(n36698));
    SB_LUT4 div_11_i1706_3_lut_3_lut (.I0(n2558), .I1(n6959), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2993_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n36696), 
            .O(n6830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4270));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4271));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2993_4 (.CI(n36696), .I0(n1873), .I1(n98), .CO(n36697));
    SB_LUT4 add_2993_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n36695), 
            .O(n6831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_3 (.CI(n36695), .I0(n1874), .I1(n99), .CO(n36696));
    SB_LUT4 add_2993_2_lut (.I0(GND_net), .I1(n381), .I2(n558), .I3(VCC_net), 
            .O(n6832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2993_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2993_2 (.CI(VCC_net), .I0(n381), .I1(n558), .CO(n36695));
    SB_LUT4 add_2991_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n36694), 
            .O(n6778)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2991_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n36693), 
            .O(n6779)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_13 (.CI(n36693), .I0(n1755), .I1(n89), .CO(n36694));
    SB_LUT4 add_2991_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n36692), 
            .O(n6780)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4266));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2991_12 (.CI(n36692), .I0(n1756), .I1(n90), .CO(n36693));
    SB_LUT4 add_2991_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n36691), 
            .O(n6781)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_11 (.CI(n36691), .I0(n1757), .I1(n91), .CO(n36692));
    SB_LUT4 add_2991_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n36690), 
            .O(n6782)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_10 (.CI(n36690), .I0(n1758), .I1(n92), .CO(n36691));
    SB_LUT4 add_2991_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n36689), 
            .O(n6783)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_9 (.CI(n36689), .I0(n1759), .I1(n93), .CO(n36690));
    SB_LUT4 add_2991_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n36688), 
            .O(n6784)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1719_3_lut_3_lut (.I0(n2558), .I1(n6972), .I2(n388), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2991_8 (.CI(n36688), .I0(n1760), .I1(n94), .CO(n36689));
    SB_LUT4 add_2991_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n36687), 
            .O(n6785)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_7 (.CI(n36687), .I0(n1761), .I1(n95), .CO(n36688));
    SB_LUT4 add_2991_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n36686), 
            .O(n6786)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_6 (.CI(n36686), .I0(n1762), .I1(n96), .CO(n36687));
    SB_LUT4 add_2991_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n36685), 
            .O(n6787)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_5 (.CI(n36685), .I0(n1763), .I1(n97), .CO(n36686));
    SB_LUT4 add_2991_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n36684), 
            .O(n6788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_4 (.CI(n36684), .I0(n1764), .I1(n98), .CO(n36685));
    SB_LUT4 add_2991_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n36683), 
            .O(n6789)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4267));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2991_3 (.CI(n36683), .I0(n1765), .I1(n99), .CO(n36684));
    SB_LUT4 div_11_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4268));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4263));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4265));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1708_3_lut_3_lut (.I0(n2558), .I1(n6961), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2991_2_lut (.I0(GND_net), .I1(n380), .I2(n558), .I3(VCC_net), 
            .O(n6790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2991_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2991_2 (.CI(VCC_net), .I0(n380), .I1(n558), .CO(n36683));
    SB_LUT4 add_2989_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n36682), 
            .O(n6737)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4256));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1709_3_lut_3_lut (.I0(n2558), .I1(n6962), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1704_3_lut_3_lut (.I0(n2558), .I1(n6957), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4258));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1710_3_lut_3_lut (.I0(n2558), .I1(n6963), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4260));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2989_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n36681), 
            .O(n6738)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1711_3_lut_3_lut (.I0(n2558), .I1(n6964), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4262));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2989_12 (.CI(n36681), .I0(n1644), .I1(n90), .CO(n36682));
    SB_LUT4 div_11_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2989_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n36680), 
            .O(n6739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2989_11 (.CI(n36680), .I0(n1645), .I1(n91), .CO(n36681));
    SB_LUT4 div_11_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4254));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2989_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n36679), 
            .O(n6740)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2989_10 (.CI(n36679), .I0(n1646), .I1(n92), .CO(n36680));
    SB_LUT4 div_11_i1715_3_lut_3_lut (.I0(n2558), .I1(n6968), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31706_4_lut (.I0(n25_adj_4260), .I1(n23_adj_4258), .I2(n21_adj_4256), 
            .I3(n19_adj_4254), .O(n47267));
    defparam i31706_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2989_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n36678), 
            .O(n6741)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1712_3_lut_3_lut (.I0(n2558), .I1(n6965), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2989_9 (.CI(n36678), .I0(n1647), .I1(n93), .CO(n36679));
    SB_LUT4 add_2989_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n36677), 
            .O(n6742)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10811_4_lut (.I0(pwm_23__N_2957), .I1(n448), .I2(PWMLimit[23]), 
            .I3(n387), .O(n24225));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10811_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i31700_4_lut (.I0(n31_adj_4265), .I1(n29_adj_4263), .I2(n27_adj_4262), 
            .I3(n47267), .O(n47261));
    defparam i31700_4_lut.LUT_INIT = 16'haaab;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_1[0]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_LUT4 div_11_i1716_3_lut_3_lut (.I0(n2558), .I1(n6969), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2989_8 (.CI(n36677), .I0(n1648), .I1(n94), .CO(n36678));
    SB_LUT4 add_2989_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n36676), 
            .O(n6743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1718_3_lut_3_lut (.I0(n2558), .I1(n6971), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_i1717_3_lut_3_lut (.I0(n2558), .I1(n6970), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33061_4_lut (.I0(n37_adj_4268), .I1(n35_adj_4267), .I2(n33_adj_4266), 
            .I3(n47261), .O(n48622));
    defparam i33061_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2989_7 (.CI(n36676), .I0(n1649), .I1(n95), .CO(n36677));
    SB_LUT4 add_2989_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n36675), 
            .O(n6744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2989_6 (.CI(n36675), .I0(n1650), .I1(n96), .CO(n36676));
    SB_LUT4 i10813_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n44196), 
            .I3(GND_net), .O(n24227));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10813_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2989_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n36674), 
            .O(n6745)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1417_i18_4_lut (.I0(n384), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4253));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32866_3_lut (.I0(n18_adj_4253), .I1(n87), .I2(n41_adj_4270), 
            .I3(GND_net), .O(n48427));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32866_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2989_5 (.CI(n36674), .I0(n1651), .I1(n97), .CO(n36675));
    SB_LUT4 i32867_3_lut (.I0(n48427), .I1(n86), .I2(n43_adj_4271), .I3(GND_net), 
            .O(n48428));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32867_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34246_4_lut (.I0(r_SM_Main[2]), .I1(n46670), .I2(n46671), 
            .I3(r_SM_Main[1]), .O(n28961));
    defparam i34246_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 add_2989_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n36673), 
            .O(n6746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32558_4_lut (.I0(n41_adj_4173), .I1(n39_adj_4172), .I2(n37), 
            .I3(n47413), .O(n48119));
    defparam i32558_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_3003_25_lut (.I0(n249), .I1(n49816), .I2(n248), .I3(n36893), 
            .O(displacement_23__N_93[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3003_24_lut (.I0(n393), .I1(n49816), .I2(n392), .I3(n36892), 
            .O(displacement_23__N_93[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3003_24 (.CI(n36892), .I0(n49816), .I1(n392), .CO(n36893));
    SB_LUT4 add_3003_23_lut (.I0(n534), .I1(n49816), .I2(n533), .I3(n36891), 
            .O(displacement_23__N_93[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2989_4 (.CI(n36673), .I0(n1652), .I1(n98), .CO(n36674));
    SB_LUT4 add_2989_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n36672), 
            .O(n6747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2989_3 (.CI(n36672), .I0(n1653), .I1(n99), .CO(n36673));
    SB_LUT4 add_2989_2_lut (.I0(GND_net), .I1(n379), .I2(n558), .I3(VCC_net), 
            .O(n6748)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2989_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2989_2 (.CI(VCC_net), .I0(n379), .I1(n558), .CO(n36672));
    SB_LUT4 add_2988_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n36671), 
            .O(n6724)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2988_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n36670), 
            .O(n6725)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_11 (.CI(n36670), .I0(n1530), .I1(n91), .CO(n36671));
    SB_LUT4 add_2988_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n36669), 
            .O(n6726)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_10 (.CI(n36669), .I0(n1531), .I1(n92), .CO(n36670));
    SB_LUT4 add_2988_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n36668), 
            .O(n6727)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_9 (.CI(n36668), .I0(n1532), .I1(n93), .CO(n36669));
    SB_LUT4 add_2988_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n36667), 
            .O(n6728)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_8 (.CI(n36667), .I0(n1533), .I1(n94), .CO(n36668));
    SB_LUT4 add_2988_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n36666), 
            .O(n6729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_7 (.CI(n36666), .I0(n1534), .I1(n95), .CO(n36667));
    SB_LUT4 add_2988_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n36665), 
            .O(n6730)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_6 (.CI(n36665), .I0(n1535), .I1(n96), .CO(n36666));
    SB_LUT4 add_2988_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n36664), 
            .O(n6731)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_5 (.CI(n36664), .I0(n1536), .I1(n97), .CO(n36665));
    SB_LUT4 add_2988_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n36663), 
            .O(n6732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_4 (.CI(n36663), .I0(n1537), .I1(n98), .CO(n36664));
    SB_LUT4 add_2988_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n36662), 
            .O(n6733)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1714_3_lut_3_lut (.I0(n2558), .I1(n6967), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2988_3 (.CI(n36662), .I0(n1538), .I1(n99), .CO(n36663));
    SB_LUT4 i32413_4_lut (.I0(n43_adj_4271), .I1(n41_adj_4270), .I2(n29_adj_4263), 
            .I3(n47265), .O(n47974));
    defparam i32413_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2988_2_lut (.I0(GND_net), .I1(n378), .I2(n558), .I3(VCC_net), 
            .O(n6734)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2988_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2988_2 (.CI(VCC_net), .I0(n378), .I1(n558), .CO(n36662));
    SB_LUT4 div_11_LessThan_1417_i26_3_lut (.I0(n24_adj_4259), .I1(n93), 
            .I2(n29_adj_4263), .I3(GND_net), .O(n26_adj_4261));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32170_3_lut (.I0(n48428), .I1(n85), .I2(n45_adj_4272), .I3(GND_net), 
            .O(n47731));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32170_3_lut.LUT_INIT = 16'h3a3a;
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_11_pad (.PACKAGE_PIN(PIN_11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_11_c_5)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_11_pad.PIN_TYPE = 6'b011001;
    defparam PIN_11_pad.PULLUP = 1'b0;
    defparam PIN_11_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_23_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b000001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i10817_3_lut (.I0(quadA_debounced_adj_4057), .I1(reg_B_adj_4485[1]), 
            .I2(n43884), .I3(GND_net), .O(n24231));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10817_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1707_3_lut_3_lut (.I0(n2558), .I1(n6960), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1769_3_lut_3_lut (.I0(n2642), .I1(n6990), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1754_3_lut_3_lut (.I0(n2642), .I1(n6975), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2986_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n36661), 
            .O(n6684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1417_i30_3_lut (.I0(n22_adj_4257), .I1(n91), 
            .I2(n33_adj_4266), .I3(GND_net), .O(n30_adj_4264));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1755_3_lut_3_lut (.I0(n2642), .I1(n6976), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3003_23 (.CI(n36891), .I0(n49816), .I1(n533), .CO(n36892));
    SB_LUT4 add_3003_22_lut (.I0(n672), .I1(n49816), .I2(n671), .I3(n36890), 
            .O(displacement_23__N_93[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2986_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n36660), 
            .O(n6685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1756_3_lut_3_lut (.I0(n2642), .I1(n6977), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33330_4_lut (.I0(n30_adj_4264), .I1(n20_adj_4255), .I2(n33_adj_4266), 
            .I3(n47259), .O(n48891));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33330_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3003_22 (.CI(n36890), .I0(n49816), .I1(n671), .CO(n36891));
    SB_CARRY add_2986_10 (.CI(n36660), .I0(n1413), .I1(n92), .CO(n36661));
    SB_LUT4 add_2986_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n36659), 
            .O(n6686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_9 (.CI(n36659), .I0(n1414), .I1(n93), .CO(n36660));
    SB_LUT4 add_3003_21_lut (.I0(n807), .I1(n49816), .I2(n806), .I3(n36889), 
            .O(displacement_23__N_93[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1531_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6898), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1757_3_lut_3_lut (.I0(n2642), .I1(n6978), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2986_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n36658), 
            .O(n6687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1758_3_lut_3_lut (.I0(n2642), .I1(n6979), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33331_3_lut (.I0(n48891), .I1(n90), .I2(n35_adj_4267), .I3(GND_net), 
            .O(n48892));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33331_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33151_3_lut (.I0(n48892), .I1(n89), .I2(n37_adj_4268), .I3(GND_net), 
            .O(n48712));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33151_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2986_8 (.CI(n36658), .I0(n1415), .I1(n94), .CO(n36659));
    SB_LUT4 add_2986_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n36657), 
            .O(n6688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_7 (.CI(n36657), .I0(n1416), .I1(n95), .CO(n36658));
    SB_CARRY add_3003_21 (.CI(n36889), .I0(n49816), .I1(n806), .CO(n36890));
    SB_LUT4 add_2986_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n36656), 
            .O(n6689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32415_4_lut (.I0(n43_adj_4271), .I1(n41_adj_4270), .I2(n39_adj_4269), 
            .I3(n48622), .O(n47976));
    defparam i32415_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33166_4_lut (.I0(n47698), .I1(n48525), .I2(n43_adj_4174), 
            .I3(n48119), .O(n48727));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33166_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2986_6 (.CI(n36656), .I0(n1417), .I1(n96), .CO(n36657));
    SB_LUT4 add_3003_20_lut (.I0(n939), .I1(n49816), .I2(n938), .I3(n36888), 
            .O(displacement_23__N_93[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2986_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n36655), 
            .O(n6690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33167_3_lut (.I0(n48727), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n48728));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33167_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i10822_3_lut (.I0(setpoint[1]), .I1(n3791), .I2(n43935), .I3(GND_net), 
            .O(n24236));   // verilog/coms.v(126[12] 289[6])
    defparam i10822_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_20 (.CI(n36888), .I0(n49816), .I1(n938), .CO(n36889));
    SB_CARRY add_2986_5 (.CI(n36655), .I0(n1418), .I1(n97), .CO(n36656));
    SB_LUT4 div_11_i1761_3_lut_3_lut (.I0(n2642), .I1(n6982), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10823_3_lut (.I0(setpoint[2]), .I1(n3792), .I2(n43935), .I3(GND_net), 
            .O(n24237));   // verilog/coms.v(126[12] 289[6])
    defparam i10823_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10824_3_lut (.I0(setpoint[3]), .I1(n3793), .I2(n43935), .I3(GND_net), 
            .O(n24238));   // verilog/coms.v(126[12] 289[6])
    defparam i10824_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10825_3_lut (.I0(setpoint[4]), .I1(n3794), .I2(n43935), .I3(GND_net), 
            .O(n24239));   // verilog/coms.v(126[12] 289[6])
    defparam i10825_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_19_lut (.I0(n1068), .I1(n49816), .I2(n1067), .I3(n36887), 
            .O(displacement_23__N_93[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1759_3_lut_3_lut (.I0(n2642), .I1(n6980), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2986_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n36654), 
            .O(n6691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10826_3_lut (.I0(setpoint[5]), .I1(n3795), .I2(n43935), .I3(GND_net), 
            .O(n24240));   // verilog/coms.v(126[12] 289[6])
    defparam i10826_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32982_4_lut (.I0(n47731), .I1(n26_adj_4261), .I2(n45_adj_4272), 
            .I3(n47974), .O(n48543));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32982_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2986_4 (.CI(n36654), .I0(n1419), .I1(n98), .CO(n36655));
    SB_LUT4 i32168_3_lut (.I0(n48712), .I1(n88), .I2(n39_adj_4269), .I3(GND_net), 
            .O(n47729));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32168_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1762_3_lut_3_lut (.I0(n2642), .I1(n6983), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32984_4_lut (.I0(n47729), .I1(n48543), .I2(n45_adj_4272), 
            .I3(n47976), .O(n48545));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32984_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1401 (.I0(n48545), .I1(n22390), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1401.LUT_INIT = 16'hceef;
    SB_LUT4 add_2986_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n36653), 
            .O(n6692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1760_3_lut_3_lut (.I0(n2642), .I1(n6981), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3003_19 (.CI(n36887), .I0(n49816), .I1(n1067), .CO(n36888));
    SB_LUT4 i10827_3_lut (.I0(setpoint[6]), .I1(n3796), .I2(n43935), .I3(GND_net), 
            .O(n24241));   // verilog/coms.v(126[12] 289[6])
    defparam i10827_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2986_3 (.CI(n36653), .I0(n1420), .I1(n99), .CO(n36654));
    SB_LUT4 i10828_3_lut (.I0(setpoint[7]), .I1(n3797), .I2(n43935), .I3(GND_net), 
            .O(n24242));   // verilog/coms.v(126[12] 289[6])
    defparam i10828_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2986_2_lut (.I0(GND_net), .I1(n377), .I2(n558), .I3(VCC_net), 
            .O(n6693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_2_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_9_pad (.PACKAGE_PIN(PIN_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_9_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_9_pad.PIN_TYPE = 6'b011001;
    defparam PIN_9_pad.PULLUP = 1'b0;
    defparam PIN_9_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c_2)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_i1775_3_lut_3_lut (.I0(n2642), .I1(n6996), .I2(n389), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10829_3_lut (.I0(setpoint[8]), .I1(n3798), .I2(n43935), .I3(GND_net), 
            .O(n24243));   // verilog/coms.v(126[12] 289[6])
    defparam i10829_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10830_3_lut (.I0(setpoint[9]), .I1(n3799), .I2(n43935), .I3(GND_net), 
            .O(n24244));   // verilog/coms.v(126[12] 289[6])
    defparam i10830_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_18_lut (.I0(n1194), .I1(n49816), .I2(n1193), .I3(n36886), 
            .O(displacement_23__N_93[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2986_2 (.CI(VCC_net), .I0(n377), .I1(n558), .CO(n36653));
    SB_CARRY add_3003_18 (.CI(n36886), .I0(n49816), .I1(n1193), .CO(n36887));
    SB_LUT4 i10831_3_lut (.I0(setpoint[10]), .I1(n3800), .I2(n43935), 
            .I3(GND_net), .O(n24245));   // verilog/coms.v(126[12] 289[6])
    defparam i10831_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2984_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n36652), 
            .O(n6644)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2984_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n36651), 
            .O(n6645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10832_3_lut (.I0(setpoint[11]), .I1(n3801), .I2(n43935), 
            .I3(GND_net), .O(n24246));   // verilog/coms.v(126[12] 289[6])
    defparam i10832_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_17_lut (.I0(n1317), .I1(n49816), .I2(n1316), .I3(n36885), 
            .O(displacement_23__N_93[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1764_3_lut_3_lut (.I0(n2642), .I1(n6985), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3003_17 (.CI(n36885), .I0(n49816), .I1(n1316), .CO(n36886));
    SB_CARRY add_2984_9 (.CI(n36651), .I0(n1293), .I1(n93), .CO(n36652));
    SB_LUT4 add_2984_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n36650), 
            .O(n6646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2984_8 (.CI(n36650), .I0(n1294), .I1(n94), .CO(n36651));
    SB_LUT4 i10833_3_lut (.I0(setpoint[12]), .I1(n3802), .I2(n43935), 
            .I3(GND_net), .O(n24247));   // verilog/coms.v(126[12] 289[6])
    defparam i10833_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1765_3_lut_3_lut (.I0(n2642), .I1(n6986), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3003_16_lut (.I0(n1437), .I1(n49816), .I2(n1436), .I3(n36884), 
            .O(displacement_23__N_93[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2984_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n36649), 
            .O(n6647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1766_3_lut_3_lut (.I0(n2642), .I1(n6987), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2984_7 (.CI(n36649), .I0(n1295), .I1(n95), .CO(n36650));
    SB_CARRY add_3003_16 (.CI(n36884), .I0(n49816), .I1(n1436), .CO(n36885));
    SB_LUT4 div_11_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2984_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n36648), 
            .O(n6648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2984_6 (.CI(n36648), .I0(n1296), .I1(n96), .CO(n36649));
    SB_LUT4 add_3003_15_lut (.I0(n1554), .I1(n49816), .I2(n1553), .I3(n36883), 
            .O(displacement_23__N_93[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2984_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n36647), 
            .O(n6649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2984_5 (.CI(n36647), .I0(n1297), .I1(n97), .CO(n36648));
    SB_LUT4 i10834_3_lut (.I0(setpoint[13]), .I1(n3803), .I2(n43935), 
            .I3(GND_net), .O(n24248));   // verilog/coms.v(126[12] 289[6])
    defparam i10834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1767_3_lut_3_lut (.I0(n2642), .I1(n6988), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10835_3_lut (.I0(setpoint[14]), .I1(n3804), .I2(n43935), 
            .I3(GND_net), .O(n24249));   // verilog/coms.v(126[12] 289[6])
    defparam i10835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2984_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n36646), 
            .O(n6650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2984_4 (.CI(n36646), .I0(n1298), .I1(n98), .CO(n36647));
    SB_CARRY add_3003_15 (.CI(n36883), .I0(n49816), .I1(n1553), .CO(n36884));
    SB_LUT4 add_2984_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n36645), 
            .O(n6651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3003_14_lut (.I0(n1668), .I1(n49816), .I2(n1667), .I3(n36882), 
            .O(displacement_23__N_93[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3003_14 (.CI(n36882), .I0(n49816), .I1(n1667), .CO(n36883));
    SB_LUT4 add_3003_13_lut (.I0(n1779), .I1(n49816), .I2(n1778), .I3(n36881), 
            .O(displacement_23__N_93[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2984_3 (.CI(n36645), .I0(n1299), .I1(n99), .CO(n36646));
    SB_LUT4 add_2984_2_lut (.I0(GND_net), .I1(n376), .I2(n558), .I3(VCC_net), 
            .O(n6652)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2984_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2984_2 (.CI(VCC_net), .I0(n376), .I1(n558), .CO(n36645));
    SB_CARRY add_3003_13 (.CI(n36881), .I0(n49816), .I1(n1778), .CO(n36882));
    SB_LUT4 i10836_3_lut (.I0(setpoint[15]), .I1(n3805), .I2(n43935), 
            .I3(GND_net), .O(n24250));   // verilog/coms.v(126[12] 289[6])
    defparam i10836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_12_lut (.I0(n1887), .I1(n49816), .I2(n1886), .I3(n36880), 
            .O(displacement_23__N_93[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i10837_3_lut (.I0(setpoint[16]), .I1(n3806), .I2(n43935), 
            .I3(GND_net), .O(n24251));   // verilog/coms.v(126[12] 289[6])
    defparam i10837_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_12 (.CI(n36880), .I0(n49816), .I1(n1886), .CO(n36881));
    SB_LUT4 div_11_i1773_3_lut_3_lut (.I0(n2642), .I1(n6994), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3003_11_lut (.I0(n1992), .I1(n49816), .I2(n1991), .I3(n36879), 
            .O(displacement_23__N_93[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i10838_3_lut (.I0(setpoint[17]), .I1(n3807), .I2(n43935), 
            .I3(GND_net), .O(n24252));   // verilog/coms.v(126[12] 289[6])
    defparam i10838_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_11 (.CI(n36879), .I0(n49816), .I1(n1991), .CO(n36880));
    SB_LUT4 add_3003_10_lut (.I0(n2094), .I1(n49816), .I2(n2093), .I3(n36878), 
            .O(displacement_23__N_93[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3003_10 (.CI(n36878), .I0(n49816), .I1(n2093), .CO(n36879));
    SB_LUT4 div_11_i1774_3_lut_3_lut (.I0(n2642), .I1(n6995), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3003_9_lut (.I0(n2193), .I1(n49816), .I2(n2192), .I3(n36877), 
            .O(displacement_23__N_93[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i10839_3_lut (.I0(setpoint[18]), .I1(n3808), .I2(n43935), 
            .I3(GND_net), .O(n24253));   // verilog/coms.v(126[12] 289[6])
    defparam i10839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1770_3_lut_3_lut (.I0(n2642), .I1(n6991), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10840_3_lut (.I0(setpoint[19]), .I1(n3809), .I2(n43935), 
            .I3(GND_net), .O(n24254));   // verilog/coms.v(126[12] 289[6])
    defparam i10840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10461_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n20471), 
            .I3(GND_net), .O(n23875));   // verilog/coms.v(126[12] 289[6])
    defparam i10461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10462_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n20471), 
            .I3(GND_net), .O(n23876));   // verilog/coms.v(126[12] 289[6])
    defparam i10462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10841_3_lut (.I0(setpoint[20]), .I1(n3810), .I2(n43935), 
            .I3(GND_net), .O(n24255));   // verilog/coms.v(126[12] 289[6])
    defparam i10841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1763_3_lut_3_lut (.I0(n2642), .I1(n6984), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10842_3_lut (.I0(setpoint[21]), .I1(n3811), .I2(n43935), 
            .I3(GND_net), .O(n24256));   // verilog/coms.v(126[12] 289[6])
    defparam i10842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1768_3_lut_3_lut (.I0(n2642), .I1(n6989), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1402 (.I0(n48728), .I1(n22369), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1402.LUT_INIT = 16'hceef;
    SB_LUT4 i10843_3_lut (.I0(setpoint[22]), .I1(n3812), .I2(n43935), 
            .I3(GND_net), .O(n24257));   // verilog/coms.v(126[12] 289[6])
    defparam i10843_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_9 (.CI(n36877), .I0(n49816), .I1(n2192), .CO(n36878));
    SB_LUT4 add_3003_8_lut (.I0(n2289_adj_4074), .I1(n49816), .I2(n2288_adj_4073), 
            .I3(n36876), .O(displacement_23__N_93[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1772_3_lut_3_lut (.I0(n2642), .I1(n6993), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3003_8 (.CI(n36876), .I0(n49816), .I1(n2288_adj_4073), 
            .CO(n36877));
    SB_LUT4 add_3003_7_lut (.I0(n2382), .I1(n49816), .I2(n2381), .I3(n36875), 
            .O(displacement_23__N_93[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3003_7 (.CI(n36875), .I0(n49816), .I1(n2381), .CO(n36876));
    SB_LUT4 div_11_i1771_3_lut_3_lut (.I0(n2642), .I1(n6992), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i888_3_lut (.I0(n1297), .I1(n6649), .I2(n1316), .I3(GND_net), 
            .O(n1417));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_6_lut (.I0(n2472), .I1(n49816), .I2(n2471), .I3(n36874), 
            .O(displacement_23__N_93[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13443_3_lut (.I0(n20471), .I1(rx_data[5]), .I2(\data_in_frame[7] [5]), 
            .I3(GND_net), .O(n23877));   // verilog/coms.v(89[13:20])
    defparam i13443_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10844_3_lut (.I0(setpoint[23]), .I1(n3813), .I2(n43935), 
            .I3(GND_net), .O(n24258));   // verilog/coms.v(126[12] 289[6])
    defparam i10844_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3003_6 (.CI(n36874), .I0(n49816), .I1(n2471), .CO(n36875));
    SB_LUT4 i10229_4_lut (.I0(n23545), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n23457), .O(n23643));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10229_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 add_3003_5_lut (.I0(n2559), .I1(n49816), .I2(n2558), .I3(n36873), 
            .O(displacement_23__N_93[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3003_5 (.CI(n36873), .I0(n49816), .I1(n2558), .CO(n36874));
    SB_LUT4 add_3003_4_lut (.I0(n2643), .I1(n49816), .I2(n2642), .I3(n36872), 
            .O(displacement_23__N_93[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3003_4 (.CI(n36872), .I0(n49816), .I1(n2642), .CO(n36873));
    SB_LUT4 div_11_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1530_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6897), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31840_4_lut (.I0(n37_adj_4177), .I1(n35), .I2(n33), .I3(n31), 
            .O(n47401));
    defparam i31840_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10464_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n20471), 
            .I3(GND_net), .O(n23878));   // verilog/coms.v(126[12] 289[6])
    defparam i10464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10465_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n20471), 
            .I3(GND_net), .O(n23879));   // verilog/coms.v(126[12] 289[6])
    defparam i10465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3003_3_lut (.I0(n2724), .I1(n49816), .I2(n2723), .I3(n36871), 
            .O(displacement_23__N_93[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_11_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i987_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3003_3 (.CI(n36871), .I0(n49816), .I1(n2723), .CO(n36872));
    SB_LUT4 div_11_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3003_2_lut (.I0(n2802), .I1(n49816), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_93[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3003_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3003_2 (.CI(VCC_net), .I0(n49816), .I1(n2801), .CO(n36871));
    SB_LUT4 div_11_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3002_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n36870), 
            .O(n6999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3002_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n36869), 
            .O(n7000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_24 (.CI(n36869), .I0(n2700), .I1(n79), .CO(n36870));
    SB_LUT4 add_3002_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n36868), 
            .O(n7001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_23 (.CI(n36868), .I0(n2701), .I1(n80), .CO(n36869));
    SB_LUT4 add_3002_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n36867), 
            .O(n7002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_22 (.CI(n36867), .I0(n2702), .I1(n81), .CO(n36868));
    SB_LUT4 add_3002_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n36866), 
            .O(n7003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_21 (.CI(n36866), .I0(n2703), .I1(n82), .CO(n36867));
    SB_LUT4 add_3002_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n36865), 
            .O(n7004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_20 (.CI(n36865), .I0(n2704), .I1(n83), .CO(n36866));
    SB_LUT4 add_3002_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n36864), 
            .O(n7005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_19 (.CI(n36864), .I0(n2705), .I1(n84), .CO(n36865));
    SB_LUT4 add_3002_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n36863), 
            .O(n7006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_18 (.CI(n36863), .I0(n2706), .I1(n85), .CO(n36864));
    SB_LUT4 div_11_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3002_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n36862), 
            .O(n7007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_17 (.CI(n36862), .I0(n2707), .I1(n86), .CO(n36863));
    SB_LUT4 add_3002_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n36861), 
            .O(n7008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_16 (.CI(n36861), .I0(n2708), .I1(n87), .CO(n36862));
    SB_LUT4 add_3002_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n36860), 
            .O(n7009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_15 (.CI(n36860), .I0(n2709), .I1(n88), .CO(n36861));
    SB_LUT4 i10466_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n20471), 
            .I3(GND_net), .O(n23880));   // verilog/coms.v(126[12] 289[6])
    defparam i10466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3002_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n36859), 
            .O(n7010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_14 (.CI(n36859), .I0(n2710), .I1(n89), .CO(n36860));
    SB_LUT4 add_3002_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n36858), 
            .O(n7011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_13 (.CI(n36858), .I0(n2711), .I1(n90), .CO(n36859));
    SB_LUT4 add_3002_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n36857), 
            .O(n7012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_12 (.CI(n36857), .I0(n2712), .I1(n91), .CO(n36858));
    SB_LUT4 add_3002_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n36856), 
            .O(n7013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_11 (.CI(n36856), .I0(n2713), .I1(n92), .CO(n36857));
    SB_LUT4 add_3002_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n36855), 
            .O(n7014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_10 (.CI(n36855), .I0(n2714), .I1(n93), .CO(n36856));
    SB_LUT4 add_3002_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n36854), 
            .O(n7015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_9 (.CI(n36854), .I0(n2715), .I1(n94), .CO(n36855));
    SB_LUT4 add_3002_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n36853), 
            .O(n7016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_8 (.CI(n36853), .I0(n2716), .I1(n95), .CO(n36854));
    SB_LUT4 add_3002_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n36852), 
            .O(n7017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_7 (.CI(n36852), .I0(n2717), .I1(n96), .CO(n36853));
    SB_LUT4 add_3002_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n36851), 
            .O(n7018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3002_6 (.CI(n36851), .I0(n2718), .I1(n97), .CO(n36852));
    SB_LUT4 add_3002_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n36850), 
            .O(n7019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2981_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n36614), 
            .O(n6573)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2981_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n36613), 
            .O(n6574)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2981_8 (.CI(n36613), .I0(n1170), .I1(n94), .CO(n36614));
    SB_CARRY add_3002_5 (.CI(n36850), .I0(n2719), .I1(n98), .CO(n36851));
    SB_LUT4 add_2981_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n36612), 
            .O(n6575)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2981_7 (.CI(n36612), .I0(n1171), .I1(n95), .CO(n36613));
    SB_LUT4 i10226_4_lut (.I0(n23545), .I1(r_Bit_Index[2]), .I2(n4010), 
            .I3(n23457), .O(n23640));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10226_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 add_2981_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n36611), 
            .O(n6576)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3002_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n36849), 
            .O(n7020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2981_6 (.CI(n36611), .I0(n1172), .I1(n96), .CO(n36612));
    SB_LUT4 add_2981_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n36610), 
            .O(n6577)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2981_5 (.CI(n36610), .I0(n1173), .I1(n97), .CO(n36611));
    SB_LUT4 add_2981_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n36609), 
            .O(n6578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2981_4 (.CI(n36609), .I0(n1174), .I1(n98), .CO(n36610));
    SB_LUT4 add_2981_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n36608), 
            .O(n6579)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2981_3 (.CI(n36608), .I0(n1175), .I1(n99), .CO(n36609));
    SB_CARRY add_3002_4 (.CI(n36849), .I0(n2720), .I1(n99), .CO(n36850));
    SB_LUT4 add_2981_2_lut (.I0(GND_net), .I1(n375), .I2(n558), .I3(VCC_net), 
            .O(n6580)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2981_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2981_2 (.CI(VCC_net), .I0(n375), .I1(n558), .CO(n36608));
    SB_LUT4 i10223_4_lut (.I0(n23547), .I1(r_Bit_Index_adj_4478[1]), .I2(r_Bit_Index_adj_4478[0]), 
            .I3(n23463), .O(n23637));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10223_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i10467_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n20471), 
            .I3(GND_net), .O(n23881));   // verilog/coms.v(126[12] 289[6])
    defparam i10467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3002_3_lut (.I0(GND_net), .I1(n390), .I2(n558), .I3(n36848), 
            .O(n7021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3002_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10468_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n20471), 
            .I3(GND_net), .O(n23882));   // verilog/coms.v(126[12] 289[6])
    defparam i10468_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3002_3 (.CI(n36848), .I0(n390), .I1(n558), .CO(n36849));
    SB_LUT4 i10220_4_lut (.I0(n23547), .I1(r_Bit_Index_adj_4478[2]), .I2(n4032), 
            .I3(n23463), .O(n23634));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10220_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i10216_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[1]), .I2(n320), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23630));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10216_4_lut.LUT_INIT = 16'h88a0;
    SB_CARRY add_3002_2 (.CI(VCC_net), .I0(n391), .I1(VCC_net), .CO(n36848));
    SB_LUT4 i10213_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[2]), .I2(n319), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23627));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10213_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 add_3001_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n36847), 
            .O(n6975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10210_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[3]), .I2(n318), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23624));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10210_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10207_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[4]), .I2(n317), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23621));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10207_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10204_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[5]), .I2(n316), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23618));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10204_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10201_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[6]), .I2(n315), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23615));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10201_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i10198_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[7]), .I2(n314), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23612));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10198_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_11_LessThan_985_i42_3_lut (.I0(n34_adj_4176), .I1(n91), 
            .I2(n45_adj_4182), .I3(GND_net), .O(n42_adj_4180));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_985_i30_4_lut (.I0(n378), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32888_3_lut (.I0(n30), .I1(n95), .I2(n37_adj_4177), .I3(GND_net), 
            .O(n48449));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32888_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32889_3_lut (.I0(n48449), .I1(n94), .I2(n39_adj_4178), .I3(GND_net), 
            .O(n48450));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32889_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31836_4_lut (.I0(n43_adj_4181), .I1(n41_adj_4179), .I2(n39_adj_4178), 
            .I3(n47401), .O(n47397));
    defparam i31836_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32966_4_lut (.I0(n42_adj_4180), .I1(n32_adj_4175), .I2(n45_adj_4182), 
            .I3(n47395), .O(n48527));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32966_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32140_3_lut (.I0(n48450), .I1(n93), .I2(n41_adj_4179), .I3(GND_net), 
            .O(n47701));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32140_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33362_4_lut (.I0(n47701), .I1(n48527), .I2(n45_adj_4182), 
            .I3(n47397), .O(n48923));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33362_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1403 (.I0(n48923), .I1(n22372), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1403.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i967_3_lut (.I0(n1417), .I1(n6689), .I2(n1436), .I3(GND_net), 
            .O(n1534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4183));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31826_4_lut (.I0(n35_adj_4188), .I1(n33_adj_4187), .I2(n31_adj_4185), 
            .I3(n29_adj_4183), .O(n47387));
    defparam i31826_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1062_i40_3_lut (.I0(n32_adj_4186), .I1(n91), 
            .I2(n43_adj_4193), .I3(GND_net), .O(n40_adj_4191));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1062_i28_4_lut (.I0(n379), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32886_3_lut (.I0(n28), .I1(n95), .I2(n35_adj_4188), .I3(GND_net), 
            .O(n48447));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32886_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32887_3_lut (.I0(n48447), .I1(n94), .I2(n37_adj_4189), .I3(GND_net), 
            .O(n48448));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32887_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31822_4_lut (.I0(n41_adj_4192), .I1(n39_adj_4190), .I2(n37_adj_4189), 
            .I3(n47387), .O(n47383));
    defparam i31822_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i659_1_lut.LUT_INIT = 16'h5555;
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_7_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b011001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i33300_4_lut (.I0(n40_adj_4191), .I1(n30_adj_4184), .I2(n43_adj_4193), 
            .I3(n47381), .O(n48861));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33300_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32142_3_lut (.I0(n48448), .I1(n93), .I2(n39_adj_4190), .I3(GND_net), 
            .O(n47703));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32142_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33480_4_lut (.I0(n47703), .I1(n48861), .I2(n43_adj_4193), 
            .I3(n47383), .O(n49041));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33480_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33481_3_lut (.I0(n49041), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n49042));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33481_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1404 (.I0(n49042), .I1(n22375), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1404.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1044_3_lut (.I0(n1534), .I1(n6729), .I2(n1553), .I3(GND_net), 
            .O(n1648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4194));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31812_4_lut (.I0(n33_adj_4199), .I1(n31_adj_4198), .I2(n29_adj_4196), 
            .I3(n27_adj_4194), .O(n47373));
    defparam i31812_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1137_i38_3_lut (.I0(n30_adj_4197), .I1(n91), 
            .I2(n41_adj_4204), .I3(GND_net), .O(n38_adj_4202));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1137_i26_4_lut (.I0(n380), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32884_3_lut (.I0(n26), .I1(n95), .I2(n33_adj_4199), .I3(GND_net), 
            .O(n48445));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32884_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32885_3_lut (.I0(n48445), .I1(n94), .I2(n35_adj_4200), .I3(GND_net), 
            .O(n48446));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32885_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31807_4_lut (.I0(n39_adj_4203), .I1(n37_adj_4201), .I2(n35_adj_4200), 
            .I3(n47373), .O(n47368));
    defparam i31807_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33322_4_lut (.I0(n38_adj_4202), .I1(n28_adj_4195), .I2(n41_adj_4204), 
            .I3(n47366), .O(n48883));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33322_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32146_3_lut (.I0(n48446), .I1(n93), .I2(n37_adj_4201), .I3(GND_net), 
            .O(n47707));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32146_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33494_4_lut (.I0(n47707), .I1(n48883), .I2(n41_adj_4204), 
            .I3(n47368), .O(n49055));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33494_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33495_3_lut (.I0(n49055), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n49056));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33495_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33422_3_lut (.I0(n49056), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n48983));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33422_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1405 (.I0(n48983), .I1(n22378), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1405.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1119_3_lut (.I0(n1648), .I1(n6742), .I2(n1667), .I3(GND_net), 
            .O(n1759));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10195_4_lut (.I0(n23629), .I1(r_Clock_Count_adj_4477[8]), .I2(n313), 
            .I3(r_SM_Main_adj_4476[2]), .O(n23609));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10195_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 add_3001_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n36846), 
            .O(n6976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_22 (.CI(n36846), .I0(n2619), .I1(n80), .CO(n36847));
    SB_LUT4 add_3001_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n36845), 
            .O(n6977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_21 (.CI(n36845), .I0(n2620), .I1(n81), .CO(n36846));
    SB_LUT4 add_3001_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n36844), 
            .O(n6978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4206));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31793_4_lut (.I0(n31_adj_4212), .I1(n29_adj_4210), .I2(n27_adj_4208), 
            .I3(n25_adj_4206), .O(n47354));
    defparam i31793_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_22_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[16]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_27[16]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[17]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_3001_20 (.CI(n36844), .I0(n2621), .I1(n82), .CO(n36845));
    SB_LUT4 mux_21_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_27[17]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3001_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n36843), 
            .O(n6979)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_19 (.CI(n36843), .I0(n2622), .I1(n83), .CO(n36844));
    SB_LUT4 add_3001_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n36842), 
            .O(n6980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_18 (.CI(n36842), .I0(n2623), .I1(n84), .CO(n36843));
    SB_LUT4 add_3001_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n36841), 
            .O(n6981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_17 (.CI(n36841), .I0(n2624), .I1(n85), .CO(n36842));
    SB_LUT4 add_3001_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n36840), 
            .O(n6982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_16 (.CI(n36840), .I0(n2625), .I1(n86), .CO(n36841));
    SB_LUT4 add_3001_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n36839), 
            .O(n6983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_15 (.CI(n36839), .I0(n2626), .I1(n87), .CO(n36840));
    SB_LUT4 mux_22_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[18]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3001_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n36838), 
            .O(n6984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_14 (.CI(n36838), .I0(n2627), .I1(n88), .CO(n36839));
    SB_LUT4 mux_21_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_27[18]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3001_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n36837), 
            .O(n6985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_13 (.CI(n36837), .I0(n2628), .I1(n89), .CO(n36838));
    SB_LUT4 i10477_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n20195), 
            .I3(GND_net), .O(n23891));   // verilog/coms.v(126[12] 289[6])
    defparam i10477_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3001_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n36836), 
            .O(n6986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_22_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[19]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10478_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n20195), 
            .I3(GND_net), .O(n23892));   // verilog/coms.v(126[12] 289[6])
    defparam i10478_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3001_12 (.CI(n36836), .I0(n2629), .I1(n90), .CO(n36837));
    SB_LUT4 add_3001_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n36835), 
            .O(n6987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_21_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_27[19]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3001_11 (.CI(n36835), .I0(n2630), .I1(n91), .CO(n36836));
    SB_LUT4 mux_22_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[20]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_3001_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n36834), 
            .O(n6988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_10 (.CI(n36834), .I0(n2631), .I1(n92), .CO(n36835));
    SB_LUT4 add_3001_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n36833), 
            .O(n6989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_9 (.CI(n36833), .I0(n2632), .I1(n93), .CO(n36834));
    SB_LUT4 mux_21_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_27[20]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14978_3_lut (.I0(n20195), .I1(rx_data[5]), .I2(\data_in_frame[5] [5]), 
            .I3(GND_net), .O(n23893));   // verilog/coms.v(89[13:20])
    defparam i14978_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3001_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n36832), 
            .O(n6990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_8 (.CI(n36832), .I0(n2633), .I1(n94), .CO(n36833));
    SB_LUT4 add_3001_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n36831), 
            .O(n6991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_7 (.CI(n36831), .I0(n2634), .I1(n95), .CO(n36832));
    SB_LUT4 add_3001_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n36830), 
            .O(n6992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_6 (.CI(n36830), .I0(n2635), .I1(n96), .CO(n36831));
    SB_LUT4 add_3001_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n36829), 
            .O(n6993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_LessThan_1210_i36_3_lut (.I0(n28_adj_4209), .I1(n91), 
            .I2(n39_adj_4218), .I3(GND_net), .O(n36_adj_4216));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1210_i24_4_lut (.I0(n381), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4205));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_1210_i32_3_lut (.I0(n30_adj_4211), .I1(n93), 
            .I2(n35_adj_4215), .I3(GND_net), .O(n32_adj_4213));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31787_4_lut (.I0(n37_adj_4217), .I1(n35_adj_4215), .I2(n33_adj_4214), 
            .I3(n47354), .O(n47348));
    defparam i31787_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33324_4_lut (.I0(n36_adj_4216), .I1(n26_adj_4207), .I2(n39_adj_4218), 
            .I3(n47343), .O(n48885));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33324_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32970_4_lut (.I0(n32_adj_4213), .I1(n24_adj_4205), .I2(n35_adj_4215), 
            .I3(n47352), .O(n48531));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32970_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33498_4_lut (.I0(n48531), .I1(n48885), .I2(n39_adj_4218), 
            .I3(n47348), .O(n49059));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33498_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33499_3_lut (.I0(n49059), .I1(n90), .I2(n1865), .I3(GND_net), 
            .O(n49060));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33499_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33412_3_lut (.I0(n49060), .I1(n89), .I2(n1864), .I3(GND_net), 
            .O(n48973));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33412_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i32972_3_lut (.I0(n48973), .I1(n88), .I2(n1863), .I3(GND_net), 
            .O(n48533));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32972_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1406 (.I0(n48533), .I1(n22381), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1406.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1192_3_lut (.I0(n1759), .I1(n6783), .I2(n1778), .I3(GND_net), 
            .O(n1867));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1263_3_lut (.I0(n1867), .I1(n6824), .I2(n1886), .I3(GND_net), 
            .O(n1972));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4232));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4222));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4220));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31762_4_lut (.I0(n29_adj_4226), .I1(n27_adj_4224), .I2(n25_adj_4222), 
            .I3(n23_adj_4220), .O(n47323));
    defparam i31762_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31756_4_lut (.I0(n35_adj_4231), .I1(n33_adj_4229), .I2(n31_adj_4228), 
            .I3(n47323), .O(n47317));
    defparam i31756_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3001_5 (.CI(n36829), .I0(n2636), .I1(n97), .CO(n36830));
    SB_LUT4 mux_22_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[21]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_27[21]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10663_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24077));   // verilog/coms.v(126[12] 289[6])
    defparam i10663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[22]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_27[22]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3001_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n36828), 
            .O(n6994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n22283), 
            .I3(GND_net), .O(n15_adj_4056));   // verilog/TinyFPGA_B.v(138[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i4_4_lut (.I0(control_mode[3]), .I1(control_mode[5]), .I2(control_mode[4]), 
            .I3(control_mode[7]), .O(n10_adj_4431));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3001_4 (.CI(n36828), .I0(n2637), .I1(n98), .CO(n36829));
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4431), .I2(control_mode[2]), 
            .I3(GND_net), .O(n22283));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_22_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[23]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_27[23]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4034));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4035));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3001_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n36827), 
            .O(n6995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10480_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n20195), 
            .I3(GND_net), .O(n23894));   // verilog/coms.v(126[12] 289[6])
    defparam i10480_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3001_3 (.CI(n36827), .I0(n2638), .I1(n99), .CO(n36828));
    SB_LUT4 add_3001_2_lut (.I0(GND_net), .I1(n389), .I2(n558), .I3(VCC_net), 
            .O(n6996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3001_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3001_2 (.CI(VCC_net), .I0(n389), .I1(n558), .CO(n36827));
    SB_LUT4 add_3000_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n36826), 
            .O(n6952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3000_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n36825), 
            .O(n6953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_21 (.CI(n36825), .I0(n2535), .I1(n81), .CO(n36826));
    SB_LUT4 add_3000_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n36824), 
            .O(n6954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_20 (.CI(n36824), .I0(n2536), .I1(n82), .CO(n36825));
    SB_LUT4 add_3000_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n36823), 
            .O(n6955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_1[23]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_CARRY add_3000_19 (.CI(n36823), .I0(n2537), .I1(n83), .CO(n36824));
    SB_LUT4 add_3000_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n36822), 
            .O(n6956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_18 (.CI(n36822), .I0(n2538), .I1(n84), .CO(n36823));
    SB_LUT4 add_3000_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n36821), 
            .O(n6957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_17 (.CI(n36821), .I0(n2539), .I1(n85), .CO(n36822));
    SB_LUT4 add_3000_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n36820), 
            .O(n6958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_16 (.CI(n36820), .I0(n2540), .I1(n86), .CO(n36821));
    SB_LUT4 add_3000_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n36819), 
            .O(n6959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_15 (.CI(n36819), .I0(n2541), .I1(n87), .CO(n36820));
    SB_LUT4 add_3000_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n36818), 
            .O(n6960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_14 (.CI(n36818), .I0(n2542), .I1(n88), .CO(n36819));
    SB_LUT4 add_3000_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n36817), 
            .O(n6961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10664_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24078));   // verilog/coms.v(126[12] 289[6])
    defparam i10664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10665_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24079));   // verilog/coms.v(126[12] 289[6])
    defparam i10665_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3000_13 (.CI(n36817), .I0(n2543), .I1(n89), .CO(n36818));
    SB_LUT4 add_3000_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n36816), 
            .O(n6962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10481_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n20195), 
            .I3(GND_net), .O(n23895));   // verilog/coms.v(126[12] 289[6])
    defparam i10481_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10666_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24080));   // verilog/coms.v(126[12] 289[6])
    defparam i10666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10667_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24081));   // verilog/coms.v(126[12] 289[6])
    defparam i10667_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3000_12 (.CI(n36816), .I0(n2544), .I1(n90), .CO(n36817));
    SB_LUT4 add_3000_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n36815), 
            .O(n6963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_11 (.CI(n36815), .I0(n2545), .I1(n91), .CO(n36816));
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_1[22]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_LUT4 add_3000_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n36814), 
            .O(n6964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_10 (.CI(n36814), .I0(n2546), .I1(n92), .CO(n36815));
    SB_LUT4 add_3000_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n36813), 
            .O(n6965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_9 (.CI(n36813), .I0(n2547), .I1(n93), .CO(n36814));
    SB_LUT4 add_3000_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n36812), 
            .O(n6966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_8 (.CI(n36812), .I0(n2548), .I1(n94), .CO(n36813));
    SB_LUT4 add_3000_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n36811), 
            .O(n6967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_7 (.CI(n36811), .I0(n2549), .I1(n95), .CO(n36812));
    SB_LUT4 add_3000_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n36810), 
            .O(n6968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_6 (.CI(n36810), .I0(n2550), .I1(n96), .CO(n36811));
    SB_LUT4 add_3000_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n36809), 
            .O(n6969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_5 (.CI(n36809), .I0(n2551), .I1(n97), .CO(n36810));
    SB_LUT4 add_3000_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n36808), 
            .O(n6970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_4 (.CI(n36808), .I0(n2552), .I1(n98), .CO(n36809));
    SB_LUT4 add_3000_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n36807), 
            .O(n6971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3000_3 (.CI(n36807), .I0(n2553), .I1(n99), .CO(n36808));
    SB_LUT4 add_3000_2_lut (.I0(GND_net), .I1(n388), .I2(n558), .I3(VCC_net), 
            .O(n6972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3000_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_1[21]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_1[20]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_1[19]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_1[18]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_1[17]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_1[16]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_1[15]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_1[14]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_1[13]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_1[12]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_1[11]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_1[10]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_1[9]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_1[8]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_1[7]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_1[6]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_1[5]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_1[4]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_1[3]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_1[2]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_1[1]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_LUT4 i10668_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24082));   // verilog/coms.v(126[12] 289[6])
    defparam i10668_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3000_2 (.CI(VCC_net), .I0(n388), .I1(n558), .CO(n36807));
    SB_LUT4 add_2999_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n36806), 
            .O(n6930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1400_3_lut (.I0(n2075), .I1(n6858), .I2(n2093), .I3(GND_net), 
            .O(n2174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10669_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24083));   // verilog/coms.v(126[12] 289[6])
    defparam i10669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i22_4_lut (.I0(n382), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4219));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_1281_i30_3_lut (.I0(n28_adj_4225), .I1(n93), 
            .I2(n33_adj_4229), .I3(GND_net), .O(n30_adj_4227));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10670_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24084));   // verilog/coms.v(126[12] 289[6])
    defparam i10670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i34_3_lut (.I0(n26_adj_4223), .I1(n91), 
            .I2(n37_adj_4232), .I3(GND_net), .O(n34_adj_4230));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10671_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24085));   // verilog/coms.v(126[12] 289[6])
    defparam i10671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33326_4_lut (.I0(n34_adj_4230), .I1(n24_adj_4221), .I2(n37_adj_4232), 
            .I3(n47315), .O(n48887));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33326_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33327_3_lut (.I0(n48887), .I1(n90), .I2(n39_adj_4233), .I3(GND_net), 
            .O(n48888));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33327_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33159_3_lut (.I0(n48888), .I1(n89), .I2(n41_adj_4234), .I3(GND_net), 
            .O(n48720));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33159_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33069_4_lut (.I0(n41_adj_4234), .I1(n39_adj_4233), .I2(n37_adj_4232), 
            .I3(n47317), .O(n48630));
    defparam i33069_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10482_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n20195), 
            .I3(GND_net), .O(n23896));   // verilog/coms.v(126[12] 289[6])
    defparam i10482_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2999_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n36805), 
            .O(n6931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10672_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24086));   // verilog/coms.v(126[12] 289[6])
    defparam i10672_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2999_20 (.CI(n36805), .I0(n2448), .I1(n82), .CO(n36806));
    SB_LUT4 i10673_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24087));   // verilog/coms.v(126[12] 289[6])
    defparam i10673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10674_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24088));   // verilog/coms.v(126[12] 289[6])
    defparam i10674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2999_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n36804), 
            .O(n6932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_19 (.CI(n36804), .I0(n2449), .I1(n83), .CO(n36805));
    SB_LUT4 add_2999_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n36803), 
            .O(n6933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10483_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n20195), 
            .I3(GND_net), .O(n23897));   // verilog/coms.v(126[12] 289[6])
    defparam i10483_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33099_4_lut (.I0(n30_adj_4227), .I1(n22_adj_4219), .I2(n33_adj_4229), 
            .I3(n47321), .O(n48660));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33099_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10484_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n20195), 
            .I3(GND_net), .O(n23898));   // verilog/coms.v(126[12] 289[6])
    defparam i10484_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2999_18 (.CI(n36803), .I0(n2450), .I1(n84), .CO(n36804));
    SB_LUT4 i10675_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24089));   // verilog/coms.v(126[12] 289[6])
    defparam i10675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2999_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n36802), 
            .O(n6934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_17 (.CI(n36802), .I0(n2451), .I1(n85), .CO(n36803));
    SB_LUT4 i10676_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24090));   // verilog/coms.v(126[12] 289[6])
    defparam i10676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10677_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24091));   // verilog/coms.v(126[12] 289[6])
    defparam i10677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10678_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24092));   // verilog/coms.v(126[12] 289[6])
    defparam i10678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4133), .I3(n37005), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_11_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4134), .I3(n37004), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_24 (.CI(n37004), .I0(GND_net), .I1(n3_adj_4134), 
            .CO(n37005));
    SB_LUT4 add_2999_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n36801), 
            .O(n6935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_16 (.CI(n36801), .I0(n2452), .I1(n86), .CO(n36802));
    SB_LUT4 div_11_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4135), .I3(n37003), .O(n4_adj_4026)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n36800), 
            .O(n6936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_15 (.CI(n36800), .I0(n2453), .I1(n87), .CO(n36801));
    SB_CARRY div_11_unary_minus_2_add_3_23 (.CI(n37003), .I0(GND_net), .I1(n4_adj_4135), 
            .CO(n37004));
    SB_LUT4 div_11_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4136), .I3(n37002), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n36799), 
            .O(n6937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_22 (.CI(n37002), .I0(GND_net), .I1(n5_adj_4136), 
            .CO(n37003));
    SB_CARRY add_2999_14 (.CI(n36799), .I0(n2454), .I1(n88), .CO(n36800));
    SB_LUT4 add_2956_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n36229), 
            .O(n5820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2956_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n36798), 
            .O(n6938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4137), .I3(n37001), .O(n6_adj_4025)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10679_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24093));   // verilog/coms.v(126[12] 289[6])
    defparam i10679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2956_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n36228), 
            .O(n5821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2956_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10680_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24094));   // verilog/coms.v(126[12] 289[6])
    defparam i10680_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2956_6 (.CI(n36228), .I0(n915), .I1(n96), .CO(n36229));
    SB_LUT4 add_2956_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n36227), 
            .O(n5822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2956_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4036));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2956_5 (.CI(n36227), .I0(n916), .I1(n97), .CO(n36228));
    SB_LUT4 add_2956_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n36226), 
            .O(n5823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2956_4_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_6_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b011001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_24_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b000001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4037));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_11_unary_minus_2_add_3_21 (.CI(n37001), .I0(GND_net), .I1(n6_adj_4137), 
            .CO(n37002));
    SB_CARRY add_2999_13 (.CI(n36798), .I0(n2455), .I1(n89), .CO(n36799));
    SB_LUT4 div_11_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4138), .I3(n37000), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2956_4 (.CI(n36226), .I0(n917), .I1(n98), .CO(n36227));
    SB_LUT4 add_2999_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n36797), 
            .O(n6939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_12 (.CI(n36797), .I0(n2456), .I1(n90), .CO(n36798));
    SB_CARRY div_11_unary_minus_2_add_3_20 (.CI(n37000), .I0(GND_net), .I1(n7_adj_4138), 
            .CO(n37001));
    SB_LUT4 div_11_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4139), .I3(n36999), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n36796), 
            .O(n6940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_11 (.CI(n36796), .I0(n2457), .I1(n91), .CO(n36797));
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4038));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_11_unary_minus_2_add_3_19 (.CI(n36999), .I0(GND_net), .I1(n8_adj_4139), 
            .CO(n37000));
    SB_LUT4 add_2999_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n36795), 
            .O(n6941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2956_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n36225), 
            .O(n5824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2956_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_10 (.CI(n36795), .I0(n2458), .I1(n92), .CO(n36796));
    SB_CARRY add_2956_3 (.CI(n36225), .I0(n918), .I1(n99), .CO(n36226));
    SB_LUT4 div_11_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4140), .I3(n36998), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n36794), 
            .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2956_2_lut (.I0(GND_net), .I1(n373), .I2(n558), .I3(VCC_net), 
            .O(n5825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2956_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_9 (.CI(n36794), .I0(n2459), .I1(n93), .CO(n36795));
    SB_CARRY add_2956_2 (.CI(VCC_net), .I0(n373), .I1(n558), .CO(n36225));
    SB_CARRY div_11_unary_minus_2_add_3_18 (.CI(n36998), .I0(GND_net), .I1(n9_adj_4140), 
            .CO(n36999));
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4039));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4141), .I3(n36997), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_17 (.CI(n36997), .I0(GND_net), .I1(n10_adj_4141), 
            .CO(n36998));
    SB_LUT4 add_2999_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n36793), 
            .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_8 (.CI(n36793), .I0(n2460), .I1(n94), .CO(n36794));
    SB_LUT4 div_11_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4142), .I3(n36996), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n36792), 
            .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_16 (.CI(n36996), .I0(GND_net), .I1(n11_adj_4142), 
            .CO(n36997));
    SB_CARRY add_2999_7 (.CI(n36792), .I0(n2461), .I1(n95), .CO(n36793));
    SB_LUT4 add_2999_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n36791), 
            .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_6 (.CI(n36791), .I0(n2462), .I1(n96), .CO(n36792));
    SB_LUT4 add_2999_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n36790), 
            .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4143), .I3(n36995), .O(n12)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_5 (.CI(n36790), .I0(n2463), .I1(n97), .CO(n36791));
    SB_LUT4 add_2999_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n36789), 
            .O(n6947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_15 (.CI(n36995), .I0(GND_net), .I1(n12_adj_4143), 
            .CO(n36996));
    SB_CARRY add_2999_4 (.CI(n36789), .I0(n2464), .I1(n98), .CO(n36790));
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4040));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2999_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n36788), 
            .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4144), .I3(n36994), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_14 (.CI(n36994), .I0(GND_net), .I1(n13_adj_4144), 
            .CO(n36995));
    SB_CARRY add_2999_3 (.CI(n36788), .I0(n2465), .I1(n99), .CO(n36789));
    SB_LUT4 div_11_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4145), .I3(n36993), .O(n14)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_2_lut (.I0(GND_net), .I1(n387_adj_4068), .I2(n558), 
            .I3(VCC_net), .O(n6949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_2 (.CI(VCC_net), .I0(n387_adj_4068), .I1(n558), 
            .CO(n36788));
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4041));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10681_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24095));   // verilog/coms.v(126[12] 289[6])
    defparam i10681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2998_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n36787), 
            .O(n6909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_13 (.CI(n36993), .I0(GND_net), .I1(n14_adj_4145), 
            .CO(n36994));
    SB_LUT4 add_2998_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n36786), 
            .O(n6910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_19 (.CI(n36786), .I0(n2358), .I1(n83), .CO(n36787));
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4042));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2998_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n36785), 
            .O(n6911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4146), .I3(n36992), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_12 (.CI(n36992), .I0(GND_net), .I1(n15_adj_4146), 
            .CO(n36993));
    SB_CARRY add_2998_18 (.CI(n36785), .I0(n2359), .I1(n84), .CO(n36786));
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4043));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2998_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n36784), 
            .O(n6912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_17 (.CI(n36784), .I0(n2360), .I1(n85), .CO(n36785));
    SB_LUT4 div_11_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4147), .I3(n36991), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_11 (.CI(n36991), .I0(GND_net), .I1(n16_adj_4147), 
            .CO(n36992));
    SB_LUT4 div_11_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4148), .I3(n36990), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4044));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_11_unary_minus_2_add_3_10 (.CI(n36990), .I0(GND_net), .I1(n17_adj_4148), 
            .CO(n36991));
    SB_LUT4 add_2998_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n36783), 
            .O(n6913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_16 (.CI(n36783), .I0(n2361), .I1(n86), .CO(n36784));
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4045));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10682_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24096));   // verilog/coms.v(126[12] 289[6])
    defparam i10682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4149), .I3(n36989), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2998_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n36782), 
            .O(n6914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_9 (.CI(n36989), .I0(GND_net), .I1(n18_adj_4149), 
            .CO(n36990));
    SB_CARRY add_2998_15 (.CI(n36782), .I0(n2362), .I1(n87), .CO(n36783));
    SB_LUT4 add_2998_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n36781), 
            .O(n6915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4046));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4150), .I3(n36988), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_8 (.CI(n36988), .I0(GND_net), .I1(n19_adj_4150), 
            .CO(n36989));
    SB_CARRY add_2998_14 (.CI(n36781), .I0(n2363), .I1(n88), .CO(n36782));
    SB_LUT4 add_2998_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n36780), 
            .O(n6916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_13 (.CI(n36780), .I0(n2364), .I1(n89), .CO(n36781));
    SB_LUT4 div_11_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4151), .I3(n36987), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2998_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n36779), 
            .O(n6917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_7 (.CI(n36987), .I0(GND_net), .I1(n20_adj_4151), 
            .CO(n36988));
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4047));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32160_3_lut (.I0(n48720), .I1(n88), .I2(n43_adj_4235), .I3(GND_net), 
            .O(n47721));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32160_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2998_12 (.CI(n36779), .I0(n2365), .I1(n90), .CO(n36780));
    SB_LUT4 div_11_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4152), .I3(n36986), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_6 (.CI(n36986), .I0(GND_net), .I1(n21_adj_4152), 
            .CO(n36987));
    SB_LUT4 add_2998_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n36778), 
            .O(n6918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_11_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_19_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b000001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_11_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4153), .I3(n36985), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4048));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2998_11 (.CI(n36778), .I0(n2366), .I1(n91), .CO(n36779));
    SB_LUT4 div_11_i1529_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6896), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2998_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n36777), 
            .O(n6919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_5 (.CI(n36985), .I0(GND_net), .I1(n22_adj_4153), 
            .CO(n36986));
    SB_LUT4 div_11_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4154), .I3(n36984), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_10 (.CI(n36777), .I0(n2367), .I1(n92), .CO(n36778));
    SB_LUT4 add_2998_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n36776), 
            .O(n6920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_2_add_3_4 (.CI(n36984), .I0(GND_net), .I1(n23_adj_4154), 
            .CO(n36985));
    SB_LUT4 div_11_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4155), .I3(n36983), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_9 (.CI(n36776), .I0(n2368), .I1(n93), .CO(n36777));
    SB_LUT4 add_2998_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n36775), 
            .O(n6921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33298_4_lut (.I0(n47721), .I1(n48660), .I2(n43_adj_4235), 
            .I3(n48630), .O(n48859));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33298_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2998_8 (.CI(n36775), .I0(n2369), .I1(n94), .CO(n36776));
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4049));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_11_unary_minus_2_add_3_3 (.CI(n36983), .I0(GND_net), .I1(n24_adj_4155), 
            .CO(n36984));
    SB_LUT4 add_2998_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n36774), 
            .O(n6922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n384));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2998_7 (.CI(n36774), .I0(n2370), .I1(n95), .CO(n36775));
    SB_LUT4 add_2998_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n36773), 
            .O(n6923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_6 (.CI(n36773), .I0(n2371), .I1(n96), .CO(n36774));
    SB_LUT4 div_11_i1409_3_lut (.I0(n383), .I1(n6867), .I2(n2093), .I3(GND_net), 
            .O(n2183));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4156), .I3(VCC_net), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10683_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24097));   // verilog/coms.v(126[12] 289[6])
    defparam i10683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2998_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n36772), 
            .O(n6924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10684_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24098));   // verilog/coms.v(126[12] 289[6])
    defparam i10684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4050));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2998_5 (.CI(n36772), .I0(n2372), .I1(n97), .CO(n36773));
    SB_LUT4 i10685_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24099));   // verilog/coms.v(126[12] 289[6])
    defparam i10685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22345), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4051));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_11_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4156), 
            .CO(n36983));
    SB_LUT4 div_11_i1408_3_lut (.I0(n2083), .I1(n6866), .I2(n2093), .I3(GND_net), 
            .O(n2182));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2998_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n36771), 
            .O(n6925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34257_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n49816));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i34257_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2998_4 (.CI(n36771), .I0(n2373), .I1(n98), .CO(n36772));
    SB_LUT4 add_2998_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n36770), 
            .O(n6926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4109), .I3(n36982), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i33299_3_lut (.I0(n48859), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n48860));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33299_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_11_i1407_3_lut (.I0(n2082), .I1(n6865), .I2(n2093), .I3(GND_net), 
            .O(n2181));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10493_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n42406), 
            .I3(GND_net), .O(n23907));   // verilog/coms.v(126[12] 289[6])
    defparam i10493_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2_adj_4024), 
            .I3(n5_adj_4437), .O(n43086));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_CARRY add_2998_3 (.CI(n36770), .I0(n2374), .I1(n99), .CO(n36771));
    SB_LUT4 i10494_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n42406), 
            .I3(GND_net), .O(n23908));   // verilog/coms.v(126[12] 289[6])
    defparam i10494_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2998_2_lut (.I0(GND_net), .I1(n386), .I2(n558), .I3(VCC_net), 
            .O(n6927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2998_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4110), .I3(n36981), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2998_2 (.CI(VCC_net), .I0(n386), .I1(n558), .CO(n36770));
    SB_LUT4 add_2997_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n36769), 
            .O(n6889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_24 (.CI(n36981), .I0(GND_net), .I1(n3_adj_4110), 
            .CO(n36982));
    SB_LUT4 add_2997_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n36768), 
            .O(n6890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_18 (.CI(n36768), .I0(n2265), .I1(n84), .CO(n36769));
    SB_LUT4 div_11_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4111), .I3(n36980), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n36767), 
            .O(n6891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_17 (.CI(n36767), .I0(n2266), .I1(n85), .CO(n36768));
    SB_CARRY div_11_unary_minus_4_add_3_23 (.CI(n36980), .I0(GND_net), .I1(n4_adj_4111), 
            .CO(n36981));
    SB_LUT4 add_2997_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n36766), 
            .O(n6892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_16 (.CI(n36766), .I0(n2267), .I1(n86), .CO(n36767));
    SB_LUT4 div_11_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4112), .I3(n36979), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n36765), 
            .O(n6893)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_15 (.CI(n36765), .I0(n2268), .I1(n87), .CO(n36766));
    SB_CARRY div_11_unary_minus_4_add_3_22 (.CI(n36979), .I0(GND_net), .I1(n5_adj_4112), 
            .CO(n36980));
    SB_LUT4 add_2997_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n36764), 
            .O(n6894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_14 (.CI(n36764), .I0(n2269), .I1(n88), .CO(n36765));
    SB_LUT4 i10495_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n42406), 
            .I3(GND_net), .O(n23909));   // verilog/coms.v(126[12] 289[6])
    defparam i10495_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4113), .I3(n36978), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n36763), 
            .O(n6895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_13 (.CI(n36763), .I0(n2270), .I1(n89), .CO(n36764));
    SB_LUT4 add_2997_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n36762), 
            .O(n6896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_21 (.CI(n36978), .I0(GND_net), .I1(n6_adj_4113), 
            .CO(n36979));
    SB_LUT4 div_11_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4114), .I3(n36977), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_12 (.CI(n36762), .I0(n2271), .I1(n90), .CO(n36763));
    SB_LUT4 add_2997_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n36761), 
            .O(n6897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_11 (.CI(n36761), .I0(n2272), .I1(n91), .CO(n36762));
    SB_CARRY div_11_unary_minus_4_add_3_20 (.CI(n36977), .I0(GND_net), .I1(n7_adj_4114), 
            .CO(n36978));
    SB_LUT4 add_2997_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n36760), 
            .O(n6898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4115), .I3(n36976), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_10 (.CI(n36760), .I0(n2273), .I1(n92), .CO(n36761));
    SB_LUT4 add_2997_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n36759), 
            .O(n6899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10496_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n42406), 
            .I3(GND_net), .O(n23910));   // verilog/coms.v(126[12] 289[6])
    defparam i10496_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2997_9 (.CI(n36759), .I0(n2274), .I1(n93), .CO(n36760));
    SB_CARRY div_11_unary_minus_4_add_3_19 (.CI(n36976), .I0(GND_net), .I1(n8_adj_4115), 
            .CO(n36977));
    SB_LUT4 add_2997_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n36758), 
            .O(n6900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1407 (.I0(n48860), .I1(n22384), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1407.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1268_3_lut (.I0(n1872), .I1(n6829), .I2(n1886), .I3(GND_net), 
            .O(n1977));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1337_3_lut (.I0(n1977), .I1(n6845), .I2(n1991), .I3(GND_net), 
            .O(n2079));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1337_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2997_8 (.CI(n36758), .I0(n2275), .I1(n94), .CO(n36759));
    SB_LUT4 div_11_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4116), .I3(n36975), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n36757), 
            .O(n6901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10497_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n42406), 
            .I3(GND_net), .O(n23911));   // verilog/coms.v(126[12] 289[6])
    defparam i10497_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2997_7 (.CI(n36757), .I0(n2276), .I1(n95), .CO(n36758));
    SB_LUT4 div_11_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY div_11_unary_minus_4_add_3_18 (.CI(n36975), .I0(GND_net), .I1(n9_adj_4116), 
            .CO(n36976));
    SB_LUT4 add_2997_6_lut (.I0(GND_net), .I1(n2277_adj_4069), .I2(n96), 
            .I3(n36756), .O(n6902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_6 (.CI(n36756), .I0(n2277_adj_4069), .I1(n96), .CO(n36757));
    SB_LUT4 div_11_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4117), .I3(n36974), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_17 (.CI(n36974), .I0(GND_net), .I1(n10_adj_4117), 
            .CO(n36975));
    SB_LUT4 add_2997_5_lut (.I0(GND_net), .I1(n2278_adj_4070), .I2(n97), 
            .I3(n36755), .O(n6903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_5 (.CI(n36755), .I0(n2278_adj_4070), .I1(n97), .CO(n36756));
    SB_LUT4 i10498_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n42406), 
            .I3(GND_net), .O(n23912));   // verilog/coms.v(126[12] 289[6])
    defparam i10498_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2997_4_lut (.I0(GND_net), .I1(n2279_adj_4071), .I2(n98), 
            .I3(n36754), .O(n6904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1339_3_lut (.I0(n1979), .I1(n6847), .I2(n1991), .I3(GND_net), 
            .O(n2081));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1339_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10499_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n42406), 
            .I3(GND_net), .O(n23913));   // verilog/coms.v(126[12] 289[6])
    defparam i10499_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2997_4 (.CI(n36754), .I0(n2279_adj_4071), .I1(n98), .CO(n36755));
    SB_LUT4 div_11_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4118), .I3(n36973), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2997_3_lut (.I0(GND_net), .I1(n2280_adj_4072), .I2(n99), 
            .I3(n36753), .O(n6905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2997_3 (.CI(n36753), .I0(n2280_adj_4072), .I1(n99), .CO(n36754));
    GND i1 (.Y(GND_net));
    SB_LUT4 i10500_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n42406), 
            .I3(GND_net), .O(n23914));   // verilog/coms.v(126[12] 289[6])
    defparam i10500_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[7] [6]), .I1(n22501), .I2(GND_net), 
            .I3(GND_net), .O(n43011));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1408 (.I0(n42896), .I1(n23013), .I2(\data_in_frame[7] [5]), 
            .I3(n43011), .O(n10_adj_4440));   // verilog/coms.v(94[12:25])
    defparam i4_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1409 (.I0(n42621), .I1(n10_adj_4440), .I2(\data_in_frame[9] [7]), 
            .I3(GND_net), .O(n38879));   // verilog/coms.v(94[12:25])
    defparam i5_3_lut_adj_1409.LUT_INIT = 16'h9696;
    SB_LUT4 div_11_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4126));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4125));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4124));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_11_unary_minus_4_add_3_16 (.CI(n36973), .I0(GND_net), .I1(n11_adj_4118), 
            .CO(n36974));
    SB_LUT4 add_2997_2_lut (.I0(GND_net), .I1(n385), .I2(n558), .I3(VCC_net), 
            .O(n6906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2997_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_i1528_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6895), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4239));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10509_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n42405), 
            .I3(GND_net), .O(n23923));   // verilog/coms.v(126[12] 289[6])
    defparam i10509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10510_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n42405), 
            .I3(GND_net), .O(n23924));   // verilog/coms.v(126[12] 289[6])
    defparam i10510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4241));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4243));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1410 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42896));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1410.LUT_INIT = 16'h6666;
    SB_CARRY add_2997_2 (.CI(VCC_net), .I0(n385), .I1(n558), .CO(n36753));
    SB_LUT4 div_11_i1340_3_lut (.I0(n1980), .I1(n6848), .I2(n1991), .I3(GND_net), 
            .O(n2082));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1340_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4119), .I3(n36972), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n36752), 
            .O(n6870)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_11_unary_minus_4_add_3_15 (.CI(n36972), .I0(GND_net), .I1(n12_adj_4119), 
            .CO(n36973));
    SB_LUT4 i10511_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n42405), 
            .I3(GND_net), .O(n23925));   // verilog/coms.v(126[12] 289[6])
    defparam i10511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4237));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4120), .I3(n36971), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10512_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n42405), 
            .I3(GND_net), .O(n23926));   // verilog/coms.v(126[12] 289[6])
    defparam i10512_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_11_unary_minus_4_add_3_14 (.CI(n36971), .I0(GND_net), .I1(n13_adj_4120), 
            .CO(n36972));
    SB_LUT4 add_2996_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n36751), 
            .O(n6871)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_11_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4121), .I3(n36970), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_17 (.CI(n36751), .I0(n2169), .I1(n85), .CO(n36752));
    SB_LUT4 add_2996_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n36750), 
            .O(n6872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_16 (.CI(n36750), .I0(n2170), .I1(n86), .CO(n36751));
    SB_CARRY div_11_unary_minus_4_add_3_13 (.CI(n36970), .I0(GND_net), .I1(n14_adj_4121), 
            .CO(n36971));
    SB_LUT4 add_2996_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n36749), 
            .O(n6873)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_93[23]), 
            .I2(n3_adj_4067), .I3(n36176), .O(displacement_23__N_1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_15 (.CI(n36749), .I0(n2171), .I1(n87), .CO(n36750));
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_93[22]), 
            .I2(n3_adj_4067), .I3(n36175), .O(displacement_23__N_1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2996_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n36748), 
            .O(n6874)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_14 (.CI(n36748), .I0(n2172), .I1(n88), .CO(n36749));
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n36175), .I0(displacement_23__N_93[22]), 
            .I1(n3_adj_4067), .CO(n36176));
    SB_LUT4 add_2996_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n36747), 
            .O(n6875)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2996_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2996_13 (.CI(n36747), .I0(n2173), .I1(n89), .CO(n36748));
    SB_LUT4 i10513_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n42405), 
            .I3(GND_net), .O(n23927));   // verilog/coms.v(126[12] 289[6])
    defparam i10513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4122), .I3(n36969), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_11_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10514_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n42405), 
            .I3(GND_net), .O(n23928));   // verilog/coms.v(126[12] 289[6])
    defparam i10514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10515_3_lut (.I0(\data_in_frame[1] [1]), .I1(rx_data[1]), .I2(n42405), 
            .I3(GND_net), .O(n23929));   // verilog/coms.v(126[12] 289[6])
    defparam i10515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10516_3_lut (.I0(\data_in_frame[1] [0]), .I1(rx_data[0]), .I2(n42405), 
            .I3(GND_net), .O(n23930));   // verilog/coms.v(126[12] 289[6])
    defparam i10516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_22_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[0]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_27[0]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[1]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_27[1]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1411 (.I0(\data_in_frame[8] [0]), .I1(n5_adj_4028), 
            .I2(GND_net), .I3(GND_net), .O(n43032));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1411.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[10] [2]), .I1(n43032), .I2(n42920), 
            .I3(\data_in_frame[8] [2]), .O(n42559));   // verilog/coms.v(94[12:25])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42633));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1413 (.I0(n22538), .I1(n42633), .I2(\data_in_frame[12] [4]), 
            .I3(n22908), .O(n10_adj_4027));   // verilog/coms.v(94[12:25])
    defparam i4_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1414 (.I0(n42559), .I1(n10_adj_4027), .I2(\data_in_frame[6] [1]), 
            .I3(GND_net), .O(n22589));   // verilog/coms.v(94[12:25])
    defparam i5_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 mux_22_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[2]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_27[2]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[3]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n22283), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_4032));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 mux_21_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_27[3]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[4]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_27[4]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1415 (.I0(control_mode[0]), .I1(n22283), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_4031));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i1_2_lut_3_lut_adj_1415.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_22_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[5]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_27[5]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[6]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_27[6]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[7]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_27[7]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[8]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_27[8]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1524_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6891), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_22_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[9]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_27[9]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[10]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_27[10]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1539_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6906), .I2(n385), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_22_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[11]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_27[11]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10657_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24071));   // verilog/coms.v(126[12] 289[6])
    defparam i10657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_26));   // verilog/TinyFPGA_B.v(73[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_22_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[12]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_27[12]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[13]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_27[13]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10658_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24072));   // verilog/coms.v(126[12] 289[6])
    defparam i10658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[14]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_27[14]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_539_i15_2_lut (.I0(pwm_count[7]), .I1(pwm[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4099));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_539_i9_2_lut (.I0(pwm_count[4]), .I1(pwm[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4095));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_539_i13_2_lut (.I0(pwm_count[6]), .I1(pwm[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4097));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_539_i11_2_lut (.I0(pwm_count[5]), .I1(pwm[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4096));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_539_i4_4_lut (.I0(pwm_count[0]), .I1(pwm[1]), .I2(pwm_count[1]), 
            .I3(pwm[0]), .O(n4_adj_4092));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i33108_3_lut (.I0(n4_adj_4092), .I1(pwm[5]), .I2(n11_adj_4096), 
            .I3(GND_net), .O(n48669));   // verilog/motorControl.v(65[19:32])
    defparam i33108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33109_3_lut (.I0(n48669), .I1(pwm[6]), .I2(n13_adj_4097), 
            .I3(GND_net), .O(n48670));   // verilog/motorControl.v(65[19:32])
    defparam i33109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31976_4_lut (.I0(n13_adj_4097), .I1(n11_adj_4096), .I2(n9_adj_4095), 
            .I3(n46779), .O(n47537));
    defparam i31976_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_539_i8_3_lut (.I0(n6_adj_4093), .I1(pwm[4]), .I2(n9_adj_4095), 
            .I3(GND_net), .O(n8_adj_4094));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32947_3_lut (.I0(n48670), .I1(pwm[7]), .I2(n15_adj_4099), 
            .I3(GND_net), .O(n14_adj_4098));   // verilog/motorControl.v(65[19:32])
    defparam i32947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32650_4_lut (.I0(n14_adj_4098), .I1(n8_adj_4094), .I2(n15_adj_4099), 
            .I3(n47537), .O(n48211));   // verilog/motorControl.v(65[19:32])
    defparam i32650_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 LessThan_542_i9_2_lut (.I0(pwm_count[4]), .I1(n872), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4107));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_542_i4_3_lut (.I0(n46619), .I1(n875), .I2(pwm_count[1]), 
            .I3(GND_net), .O(n4_adj_4104));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_11_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4132));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1406_3_lut (.I0(n2081), .I1(n6864), .I2(n2093), .I3(GND_net), 
            .O(n2180));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_542_i8_3_lut (.I0(n6_adj_4105), .I1(n872), .I2(n9_adj_4107), 
            .I3(GND_net), .O(n8_adj_4106));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33401_4_lut (.I0(n8_adj_4106), .I1(n4_adj_4104), .I2(n9_adj_4107), 
            .I3(n46762), .O(n48962));   // verilog/motorControl.v(86[28:44])
    defparam i33401_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33402_3_lut (.I0(n48962), .I1(n871), .I2(pwm_count[5]), .I3(GND_net), 
            .O(n48963));   // verilog/motorControl.v(86[28:44])
    defparam i33402_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_11_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4131));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1405_3_lut (.I0(n2080), .I1(n6863), .I2(n2093), .I3(GND_net), 
            .O(n2179));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33305_3_lut (.I0(n48963), .I1(n870), .I2(pwm_count[6]), .I3(GND_net), 
            .O(n48866));   // verilog/motorControl.v(86[28:44])
    defparam i33305_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33209_3_lut (.I0(n48866), .I1(n869), .I2(pwm_count[7]), .I3(GND_net), 
            .O(n16_adj_4108));   // verilog/motorControl.v(86[28:44])
    defparam i33209_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i12_4_lut (.I0(n857), .I1(n855), .I2(n865), .I3(n866), .O(n28_adj_4433));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_542_i18_3_lut (.I0(n16_adj_4108), .I1(n868), .I2(pwm_count[8]), 
            .I3(GND_net), .O(n2311));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i18_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i10_4_lut (.I0(n861), .I1(n856), .I2(n859), .I3(n860), .O(n26_adj_4434));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n21_adj_4436), .I1(n28_adj_4433), .I2(n862), 
            .I3(n853), .O(n30_adj_4432));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4052));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_4_lut (.I0(n2311), .I1(n864), .I2(n863), .I3(n867), .O(n25_adj_4435));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_2_lut (.I0(n400), .I1(\PID_CONTROLLER.result [20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4090));   // verilog/motorControl.v(32[23:29])
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_2_lut (.I0(n399), .I1(\PID_CONTROLLER.result [21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4091));   // verilog/motorControl.v(32[23:29])
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i17_2_lut (.I0(n406), .I1(\PID_CONTROLLER.result [14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4089));   // verilog/motorControl.v(32[23:29])
    defparam i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_22_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4056), .I3(n15_adj_4032), .O(motor_state_23__N_27[15]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_22_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_21_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_27[15]), 
            .I2(n15_adj_4031), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_2_lut_adj_1416 (.I0(n415), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4086));   // verilog/motorControl.v(32[23:29])
    defparam i6_2_lut_adj_1416.LUT_INIT = 16'h6666;
    SB_LUT4 i13_2_lut (.I0(n413), .I1(\PID_CONTROLLER.result [7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4087));   // verilog/motorControl.v(32[23:29])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10659_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24073));   // verilog/coms.v(126[12] 289[6])
    defparam i10659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10660_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24074));   // verilog/coms.v(126[12] 289[6])
    defparam i10660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10661_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24075));   // verilog/coms.v(126[12] 289[6])
    defparam i10661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10662_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24076));   // verilog/coms.v(126[12] 289[6])
    defparam i10662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31736_4_lut (.I0(n27_adj_4243), .I1(n25_adj_4241), .I2(n23_adj_4239), 
            .I3(n21_adj_4237), .O(n47297));
    defparam i31736_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_i1534_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6901), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1404_3_lut (.I0(n2079), .I1(n6862), .I2(n2093), .I3(GND_net), 
            .O(n2178));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4130));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4053));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4129));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1527_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6894), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4128));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1403_3_lut (.I0(n2078), .I1(n6861), .I2(n2093), .I3(GND_net), 
            .O(n2177));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1402_3_lut (.I0(n2077), .I1(n6860), .I2(n2093), .I3(GND_net), 
            .O(n2176));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4127));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1401_3_lut (.I0(n2076), .I1(n6859), .I2(n2093), .I3(GND_net), 
            .O(n2175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1327_3_lut (.I0(n1967), .I1(n6835), .I2(n1991), .I3(GND_net), 
            .O(n2069));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n381));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1271_3_lut (.I0(n381), .I1(n6832), .I2(n1886), .I3(GND_net), 
            .O(n1980));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i725_3_lut (.I0(n374), .I1(n6218), .I2(n1067), .I3(GND_net), 
            .O(n1175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i808_3_lut (.I0(n1175), .I1(n6579), .I2(n1193), .I3(GND_net), 
            .O(n1298));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i889_3_lut (.I0(n1298), .I1(n6650), .I2(n1316), .I3(GND_net), 
            .O(n1418));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i968_3_lut (.I0(n1418), .I1(n6690), .I2(n1436), .I3(GND_net), 
            .O(n1535));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1045_3_lut (.I0(n1535), .I1(n6730), .I2(n1553), .I3(GND_net), 
            .O(n1649));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1120_3_lut (.I0(n1649), .I1(n6743), .I2(n1667), .I3(GND_net), 
            .O(n1760));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1193_3_lut (.I0(n1760), .I1(n6784), .I2(n1778), .I3(GND_net), 
            .O(n1868));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1264_3_lut (.I0(n1868), .I1(n6825), .I2(n1886), .I3(GND_net), 
            .O(n1973));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1328_3_lut (.I0(n1968), .I1(n6836), .I2(n1991), .I3(GND_net), 
            .O(n2070));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1329_3_lut (.I0(n1969), .I1(n6837), .I2(n1991), .I3(GND_net), 
            .O(n2071));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31732_4_lut (.I0(n33_adj_4248), .I1(n31_adj_4246), .I2(n29_adj_4245), 
            .I3(n47297), .O(n47293));
    defparam i31732_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_i1330_3_lut (.I0(n1970), .I1(n6838), .I2(n1991), .I3(GND_net), 
            .O(n2072));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4252));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10649_4_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n5017), .I3(n22277), .O(n24063));   // verilog/coms.v(126[12] 289[6])
    defparam i10649_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 div_11_i1331_3_lut (.I0(n1971), .I1(n6839), .I2(n1991), .I3(GND_net), 
            .O(n2073));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4251));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1332_3_lut (.I0(n1972), .I1(n6840), .I2(n1991), .I3(GND_net), 
            .O(n2074));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4250));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4249));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n382));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1341_3_lut (.I0(n382), .I1(n6849), .I2(n1991), .I3(GND_net), 
            .O(n2083));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1341_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n383));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n376));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i891_3_lut (.I0(n376), .I1(n6652), .I2(n1316), .I3(GND_net), 
            .O(n1420));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i970_3_lut (.I0(n1420), .I1(n6692), .I2(n1436), .I3(GND_net), 
            .O(n1537));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1047_3_lut (.I0(n1537), .I1(n6732), .I2(n1553), .I3(GND_net), 
            .O(n1651));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1122_3_lut (.I0(n1651), .I1(n6745), .I2(n1667), .I3(GND_net), 
            .O(n1762));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1195_3_lut (.I0(n1762), .I1(n6786), .I2(n1778), .I3(GND_net), 
            .O(n1870));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1266_3_lut (.I0(n1870), .I1(n6827), .I2(n1886), .I3(GND_net), 
            .O(n1975));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1335_3_lut (.I0(n1975), .I1(n6843), .I2(n1991), .I3(GND_net), 
            .O(n2077));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1335_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n377));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i971_3_lut (.I0(n377), .I1(n6693), .I2(n1436), .I3(GND_net), 
            .O(n1538));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1048_3_lut (.I0(n1538), .I1(n6733), .I2(n1553), .I3(GND_net), 
            .O(n1652));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1123_3_lut (.I0(n1652), .I1(n6746), .I2(n1667), .I3(GND_net), 
            .O(n1763));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1196_3_lut (.I0(n1763), .I1(n6787), .I2(n1778), .I3(GND_net), 
            .O(n1871));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10756_3_lut (.I0(encoder1_position[1]), .I1(n2249), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24170));   // quad.v(35[10] 41[6])
    defparam i10756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1267_3_lut (.I0(n1871), .I1(n6828), .I2(n1886), .I3(GND_net), 
            .O(n1976));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21958_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4024));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i21958_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10757_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4030), 
            .I3(n22411), .O(n24171));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10757_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10758_4_lut (.I0(pwm_23__N_2957), .I1(n471), .I2(PWMLimit[0]), 
            .I3(n387), .O(n24172));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10758_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_i1336_3_lut (.I0(n1976), .I1(n6844), .I2(n1991), .I3(GND_net), 
            .O(n2078));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1336_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10269_3_lut (.I0(n23545), .I1(r_Bit_Index[0]), .I2(n23457), 
            .I3(GND_net), .O(n23683));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10269_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i10266_3_lut (.I0(n23547), .I1(r_Bit_Index_adj_4478[0]), .I2(n23463), 
            .I3(GND_net), .O(n23680));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10266_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 div_11_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4161));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1334_3_lut (.I0(n1974), .I1(n6842), .I2(n1991), .I3(GND_net), 
            .O(n2076));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1334_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4164));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4167));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4245));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4246));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4168));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10767_3_lut (.I0(encoder1_position[2]), .I1(n2248), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24181));   // quad.v(35[10] 41[6])
    defparam i10767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4248));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10768_3_lut (.I0(encoder1_position[3]), .I1(n2247), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24182));   // quad.v(35[10] 41[6])
    defparam i10768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n380));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10769_3_lut (.I0(encoder1_position[4]), .I1(n2246), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24183));   // quad.v(35[10] 41[6])
    defparam i10769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1199_3_lut (.I0(n380), .I1(n6790), .I2(n1778), .I3(GND_net), 
            .O(n1874));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10770_3_lut (.I0(encoder1_position[5]), .I1(n2245), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24184));   // quad.v(35[10] 41[6])
    defparam i10770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4177));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10771_3_lut (.I0(encoder1_position[6]), .I1(n2244), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24185));   // quad.v(35[10] 41[6])
    defparam i10771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4178));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4181));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4179));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4182));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10772_3_lut (.I0(encoder1_position[7]), .I1(n2243), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24186));   // quad.v(35[10] 41[6])
    defparam i10772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1270_3_lut (.I0(n1874), .I1(n6831), .I2(n1886), .I3(GND_net), 
            .O(n1979));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4187));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10773_3_lut (.I0(encoder1_position[8]), .I1(n2242), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24187));   // quad.v(35[10] 41[6])
    defparam i10773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1338_3_lut (.I0(n1978), .I1(n6846), .I2(n1991), .I3(GND_net), 
            .O(n2080));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1338_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4185));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4188));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10774_3_lut (.I0(encoder1_position[9]), .I1(n2241), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24188));   // quad.v(35[10] 41[6])
    defparam i10774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4189));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4192));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4190));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4193));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10775_3_lut (.I0(encoder1_position[10]), .I1(n2240), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24189));   // quad.v(35[10] 41[6])
    defparam i10775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n378));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4198));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10776_3_lut (.I0(encoder1_position[11]), .I1(n2239), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24190));   // quad.v(35[10] 41[6])
    defparam i10776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1049_3_lut (.I0(n378), .I1(n6734), .I2(n1553), .I3(GND_net), 
            .O(n1653));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4196));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4199));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10777_3_lut (.I0(encoder1_position[12]), .I1(n2238), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24191));   // quad.v(35[10] 41[6])
    defparam i10777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4200));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4203));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4201));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4204));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1124_3_lut (.I0(n1653), .I1(n6747), .I2(n1667), .I3(GND_net), 
            .O(n1764));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10778_3_lut (.I0(encoder1_position[13]), .I1(n2237), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24192));   // quad.v(35[10] 41[6])
    defparam i10778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4210));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10779_3_lut (.I0(encoder1_position[14]), .I1(n2236), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24193));   // quad.v(35[10] 41[6])
    defparam i10779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1197_3_lut (.I0(n1764), .I1(n6788), .I2(n1778), .I3(GND_net), 
            .O(n1872));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4208));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4212));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10780_3_lut (.I0(encoder1_position[15]), .I1(n2235), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24194));   // quad.v(35[10] 41[6])
    defparam i10780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4214));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4217));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4215));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4218));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10781_3_lut (.I0(encoder1_position[16]), .I1(n2234), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24195));   // quad.v(35[10] 41[6])
    defparam i10781_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10782_3_lut (.I0(encoder1_position[17]), .I1(n2233), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24196));   // quad.v(35[10] 41[6])
    defparam i10782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4226));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4228));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10783_3_lut (.I0(encoder1_position[18]), .I1(n2232), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24197));   // quad.v(35[10] 41[6])
    defparam i10783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4224));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4231));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i22014_3_lut (.I0(n648), .I1(n98), .I2(n4), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i22014_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i10784_3_lut (.I0(encoder1_position[19]), .I1(n2231), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24198));   // quad.v(35[10] 41[6])
    defparam i10784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i458_4_lut (.I0(n43088), .I1(n6), .I2(n671), .I3(n97), 
            .O(n43090));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i458_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i10785_3_lut (.I0(encoder1_position[20]), .I1(n2230), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24199));   // quad.v(35[10] 41[6])
    defparam i10785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10786_3_lut (.I0(encoder1_position[21]), .I1(n2229), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24200));   // quad.v(35[10] 41[6])
    defparam i10786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22054_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4101), .I3(GND_net), 
            .O(n8_adj_4100));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i22054_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_11_i547_4_lut (.I0(n43090), .I1(n8_adj_4100), .I2(n806), 
            .I3(n96), .O(n914));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i547_4_lut.LUT_INIT = 16'h5659;
    SB_LUT4 i10787_3_lut (.I0(encoder1_position[22]), .I1(n2228), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24201));   // quad.v(35[10] 41[6])
    defparam i10787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i634_3_lut (.I0(n914), .I1(n5820), .I2(n938), .I3(GND_net), 
            .O(n1043));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10788_3_lut (.I0(encoder1_position[23]), .I1(n2227), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n24202));   // quad.v(35[10] 41[6])
    defparam i10788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i719_3_lut (.I0(n1043), .I1(n6212), .I2(n1067), .I3(GND_net), 
            .O(n1169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10789_4_lut (.I0(pwm_23__N_2957), .I1(n470), .I2(PWMLimit[1]), 
            .I3(n387), .O(n24203));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10789_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10790_4_lut (.I0(pwm_23__N_2957), .I1(n469), .I2(PWMLimit[2]), 
            .I3(n387), .O(n24204));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10790_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_i802_3_lut (.I0(n1169), .I1(n6573), .I2(n1193), .I3(GND_net), 
            .O(n1292));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10791_4_lut (.I0(pwm_23__N_2957), .I1(n468), .I2(PWMLimit[3]), 
            .I3(n387), .O(n24205));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10791_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10792_4_lut (.I0(pwm_23__N_2957), .I1(n467), .I2(PWMLimit[4]), 
            .I3(n387), .O(n24206));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10792_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_i883_3_lut (.I0(n1292), .I1(n6644), .I2(n1316), .I3(GND_net), 
            .O(n1412));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i883_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10156_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n23570));   // verilog/coms.v(126[12] 289[6])
    defparam i10156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10794_4_lut (.I0(pwm_23__N_2957), .I1(n465), .I2(PWMLimit[6]), 
            .I3(n387), .O(n24208));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10794_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_i962_3_lut (.I0(n1412), .I1(n6684), .I2(n1436), .I3(GND_net), 
            .O(n1529));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1039_3_lut (.I0(n1529), .I1(n6724), .I2(n1553), .I3(GND_net), 
            .O(n1643));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10796_4_lut (.I0(pwm_23__N_2957), .I1(n463), .I2(PWMLimit[8]), 
            .I3(n387), .O(n24210));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10796_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10160_3_lut (.I0(\PID_CONTROLLER.err_prev [0]), .I1(\PID_CONTROLLER.err [0]), 
            .I2(n43357), .I3(GND_net), .O(n23574));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10160_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10797_4_lut (.I0(pwm_23__N_2957), .I1(n462), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24211));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10797_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10798_4_lut (.I0(pwm_23__N_2957), .I1(n461), .I2(PWMLimit[10]), 
            .I3(n387), .O(n24212));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10798_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i2_4_lut_adj_1417 (.I0(n22303), .I1(n43181), .I2(n2857), .I3(n42428), 
            .O(n44294));
    defparam i2_4_lut_adj_1417.LUT_INIT = 16'hff37;
    SB_LUT4 i10799_4_lut (.I0(pwm_23__N_2957), .I1(n460), .I2(PWMLimit[11]), 
            .I3(n387), .O(n24213));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10799_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10800_4_lut (.I0(pwm_23__N_2957), .I1(n459), .I2(PWMLimit[12]), 
            .I3(n387), .O(n24214));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10800_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_i1114_3_lut (.I0(n1643), .I1(n6737), .I2(n1667), .I3(GND_net), 
            .O(n1754));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1418 (.I0(n22309), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n44294), .I3(n20088), .O(n41786));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1418.LUT_INIT = 16'hd5f5;
    SB_LUT4 div_11_i1187_3_lut (.I0(n1754), .I1(n6778), .I2(n1778), .I3(GND_net), 
            .O(n1862));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10803_4_lut (.I0(pwm_23__N_2957), .I1(n456), .I2(PWMLimit[15]), 
            .I3(n387), .O(n24217));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10803_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10804_4_lut (.I0(pwm_23__N_2957), .I1(n455), .I2(PWMLimit[16]), 
            .I3(n387), .O(n24218));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10804_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10805_4_lut (.I0(pwm_23__N_2957), .I1(n454), .I2(PWMLimit[17]), 
            .I3(n387), .O(n24219));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10805_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10162_3_lut (.I0(encoder0_position[0]), .I1(n2300), .I2(count_enable), 
            .I3(GND_net), .O(n23576));   // quad.v(35[10] 41[6])
    defparam i10162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10163_3_lut (.I0(encoder1_position[0]), .I1(n2250), .I2(count_enable_adj_4059), 
            .I3(GND_net), .O(n23577));   // quad.v(35[10] 41[6])
    defparam i10163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10806_4_lut (.I0(pwm_23__N_2957), .I1(n453), .I2(PWMLimit[18]), 
            .I3(n387), .O(n24220));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10806_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_11_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10164_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n44196), 
            .I3(GND_net), .O(n23578));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10807_4_lut (.I0(pwm_23__N_2957), .I1(n452), .I2(PWMLimit[19]), 
            .I3(n387), .O(n24221));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10807_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1419 (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n22405));
    defparam i1_2_lut_adj_1419.LUT_INIT = 16'hdddd;
    SB_LUT4 i10165_4_lut (.I0(r_SM_Main[2]), .I1(n1), .I2(n28925), .I3(r_SM_Main[1]), 
            .O(n23579));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10165_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i10166_3_lut (.I0(quadB_debounced_adj_4058), .I1(reg_B_adj_4485[0]), 
            .I2(n43884), .I3(GND_net), .O(n23580));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12360_3_lut (.I0(r_SM_Main_adj_4476[0]), .I1(o_Tx_Serial_N_2784), 
            .I2(r_SM_Main_adj_4476[1]), .I3(GND_net), .O(n25767));   // verilog/uart_tx.v(31[16:25])
    defparam i12360_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i12361_3_lut (.I0(tx_o), .I1(n25767), .I2(r_SM_Main_adj_4476[2]), 
            .I3(GND_net), .O(n23581));
    defparam i12361_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10810_4_lut (.I0(pwm_23__N_2957), .I1(n449), .I2(PWMLimit[22]), 
            .I3(n387), .O(n24224));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10810_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10_2_lut (.I0(deadband[20]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(32[23:29])
    defparam i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10169_4_lut (.I0(r_SM_Main_adj_4476[2]), .I1(n49), .I2(r_SM_Main_2__N_2753[1]), 
            .I3(r_SM_Main_adj_4476[0]), .O(n23583));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10169_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 div_11_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(n81), .I1(n22399), .I2(GND_net), .I3(GND_net), 
            .O(n22396));
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'hdddd;
    SB_LUT4 i10170_3_lut (.I0(setpoint[0]), .I1(n3790), .I2(n43935), .I3(GND_net), 
            .O(n23584));   // verilog/coms.v(126[12] 289[6])
    defparam i10170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_2_lut (.I0(deadband[14]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(32[23:29])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i5_2_lut (.I0(deadband[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4077));   // verilog/motorControl.v(32[23:29])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1421 (.I0(n84), .I1(n22390), .I2(GND_net), .I3(GND_net), 
            .O(n22387));
    defparam i1_2_lut_adj_1421.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_2_lut (.I0(deadband[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4078));   // verilog/motorControl.v(32[23:29])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4121));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_i1258_3_lut (.I0(n1862), .I1(n6819), .I2(n1886), .I3(GND_net), 
            .O(n1967));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4120));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_2_lut_adj_1422 (.I0(deadband[21]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/motorControl.v(32[23:29])
    defparam i5_2_lut_adj_1422.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4119));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_1423 (.I0(r_SM_Main_adj_4476[1]), .I1(r_SM_Main_adj_4476[0]), 
            .I2(r_SM_Main_adj_4476[2]), .I3(r_SM_Main_2__N_2753[1]), .O(n49982));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_adj_1423.LUT_INIT = 16'h0800;
    SB_LUT4 i22046_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4102), .I3(GND_net), 
            .O(n6_adj_4101));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i22046_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_11_i459_4_lut (.I0(n648), .I1(n4), .I2(n671), .I3(n98), 
            .O(n783));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i459_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i548_4_lut (.I0(n783), .I1(n6_adj_4101), .I2(n806), 
            .I3(n97), .O(n915));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i548_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i8_2_lut (.I0(PWMLimit[20]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4083));   // verilog/motorControl.v(32[23:29])
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_i635_3_lut (.I0(n915), .I1(n5821), .I2(n938), .I3(GND_net), 
            .O(n1044));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i635_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4118));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i720_3_lut (.I0(n1044), .I1(n6213), .I2(n1067), .I3(GND_net), 
            .O(n1170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_2_lut_adj_1424 (.I0(PWMLimit[21]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4084));   // verilog/motorControl.v(32[23:29])
    defparam i8_2_lut_adj_1424.LUT_INIT = 16'h6666;
    SB_LUT4 i10230_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n28462), 
            .I3(n22416), .O(n23644));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10230_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i13_2_lut_adj_1425 (.I0(PWMLimit[14]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4082));   // verilog/motorControl.v(32[23:29])
    defparam i13_2_lut_adj_1425.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_i803_3_lut (.I0(n1170), .I1(n6574), .I2(n1193), .I3(GND_net), 
            .O(n1293));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i803_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i884_3_lut (.I0(n1293), .I1(n6645), .I2(n1316), .I3(GND_net), 
            .O(n1413));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i963_3_lut (.I0(n1413), .I1(n6685), .I2(n1436), .I3(GND_net), 
            .O(n1530));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i963_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_2_lut_adj_1426 (.I0(PWMLimit[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4079));   // verilog/motorControl.v(32[23:29])
    defparam i9_2_lut_adj_1426.LUT_INIT = 16'h6666;
    SB_LUT4 i17_2_lut_adj_1427 (.I0(PWMLimit[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4080));   // verilog/motorControl.v(32[23:29])
    defparam i17_2_lut_adj_1427.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_i1040_3_lut (.I0(n1530), .I1(n6725), .I2(n1553), .I3(GND_net), 
            .O(n1644));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1115_3_lut (.I0(n1644), .I1(n6738), .I2(n1667), .I3(GND_net), 
            .O(n1755));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1188_3_lut (.I0(n1755), .I1(n6779), .I2(n1778), .I3(GND_net), 
            .O(n1863));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1259_3_lut (.I0(n1863), .I1(n6820), .I2(n1886), .I3(GND_net), 
            .O(n1968));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n379));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1125_3_lut (.I0(n379), .I1(n6748), .I2(n1667), .I3(GND_net), 
            .O(n1765));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1198_3_lut (.I0(n1765), .I1(n6789), .I2(n1778), .I3(GND_net), 
            .O(n1873));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1269_3_lut (.I0(n1873), .I1(n6830), .I2(n1886), .I3(GND_net), 
            .O(n1978));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21998_2_lut (.I0(n371), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i21998_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i31779_3_lut (.I0(n370), .I1(n558), .I2(n533), .I3(GND_net), 
            .O(n649));
    defparam i31779_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_11_i460_4_lut (.I0(n649), .I1(n2), .I2(n671), .I3(n99), 
            .O(n784));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i460_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i549_4_lut (.I0(n784), .I1(n4_adj_4102), .I2(n806), 
            .I3(n98), .O(n916));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i549_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i636_3_lut (.I0(n916), .I1(n5822), .I2(n938), .I3(GND_net), 
            .O(n1045));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i721_3_lut (.I0(n1045), .I1(n6214), .I2(n1067), .I3(GND_net), 
            .O(n1171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10231_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n28462), 
            .I3(n22411), .O(n23645));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10231_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i10232_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4055), 
            .I3(n22416), .O(n23646));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10232_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_11_i804_3_lut (.I0(n1171), .I1(n6575), .I2(n1193), .I3(GND_net), 
            .O(n1294));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i804_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10233_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4055), 
            .I3(n22411), .O(n23647));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10233_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10234_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4054), 
            .I3(n22416), .O(n23648));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10234_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_11_i885_3_lut (.I0(n1294), .I1(n6646), .I2(n1316), .I3(GND_net), 
            .O(n1414));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10235_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4054), 
            .I3(n22411), .O(n23649));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10235_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10236_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4030), 
            .I3(n22416), .O(n23650));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10236_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_11_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4117));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i964_3_lut (.I0(n1414), .I1(n6686), .I2(n1436), .I3(GND_net), 
            .O(n1531));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1041_3_lut (.I0(n1531), .I1(n6726), .I2(n1553), .I3(GND_net), 
            .O(n1645));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1116_3_lut (.I0(n1645), .I1(n6739), .I2(n1667), .I3(GND_net), 
            .O(n1756));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1189_3_lut (.I0(n1756), .I1(n6780), .I2(n1778), .I3(GND_net), 
            .O(n1864));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4116));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1260_3_lut (.I0(n1864), .I1(n6821), .I2(n1886), .I3(GND_net), 
            .O(n1969));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4235));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n375));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i809_3_lut (.I0(n375), .I1(n6580), .I2(n1193), .I3(GND_net), 
            .O(n1299));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1538_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6905), .I2(n2280_adj_4072), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i890_3_lut (.I0(n1299), .I1(n6651), .I2(n1316), .I3(GND_net), 
            .O(n1419));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i890_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15_rep_276_2_lut (.I0(pwm_23__N_2960[14]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(GND_net), .I3(GND_net), .O(n50258));   // verilog/motorControl.v(32[23:29])
    defparam i15_rep_276_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_11_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4115));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4114));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4113));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i969_3_lut (.I0(n1419), .I1(n6691), .I2(n1436), .I3(GND_net), 
            .O(n1536));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10270_3_lut (.I0(encoder0_position[23]), .I1(n2277), .I2(count_enable), 
            .I3(GND_net), .O(n23684));   // quad.v(35[10] 41[6])
    defparam i10270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10271_3_lut (.I0(encoder0_position[22]), .I1(n2278), .I2(count_enable), 
            .I3(GND_net), .O(n23685));   // quad.v(35[10] 41[6])
    defparam i10271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10272_3_lut (.I0(encoder0_position[21]), .I1(n2279), .I2(count_enable), 
            .I3(GND_net), .O(n23686));   // quad.v(35[10] 41[6])
    defparam i10272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1046_3_lut (.I0(n1536), .I1(n6731), .I2(n1553), .I3(GND_net), 
            .O(n1650));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10273_3_lut (.I0(encoder0_position[20]), .I1(n2280), .I2(count_enable), 
            .I3(GND_net), .O(n23687));   // quad.v(35[10] 41[6])
    defparam i10273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10274_3_lut (.I0(encoder0_position[19]), .I1(n2281), .I2(count_enable), 
            .I3(GND_net), .O(n23688));   // quad.v(35[10] 41[6])
    defparam i10274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_rep_264_2_lut (.I0(pwm_23__N_2960[20]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(GND_net), .I3(GND_net), .O(n50246));   // verilog/motorControl.v(32[23:29])
    defparam i7_rep_264_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10275_3_lut (.I0(encoder0_position[18]), .I1(n2282), .I2(count_enable), 
            .I3(GND_net), .O(n23689));   // quad.v(35[10] 41[6])
    defparam i10275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1121_3_lut (.I0(n1650), .I1(n6744), .I2(n1667), .I3(GND_net), 
            .O(n1761));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10276_3_lut (.I0(encoder0_position[17]), .I1(n2283), .I2(count_enable), 
            .I3(GND_net), .O(n23690));   // quad.v(35[10] 41[6])
    defparam i10276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10277_3_lut (.I0(encoder0_position[16]), .I1(n2284), .I2(count_enable), 
            .I3(GND_net), .O(n23691));   // quad.v(35[10] 41[6])
    defparam i10277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10278_3_lut (.I0(encoder0_position[15]), .I1(n2285), .I2(count_enable), 
            .I3(GND_net), .O(n23692));   // quad.v(35[10] 41[6])
    defparam i10278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10279_3_lut (.I0(encoder0_position[14]), .I1(n2286), .I2(count_enable), 
            .I3(GND_net), .O(n23693));   // quad.v(35[10] 41[6])
    defparam i10279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10280_3_lut (.I0(encoder0_position[13]), .I1(n2287), .I2(count_enable), 
            .I3(GND_net), .O(n23694));   // quad.v(35[10] 41[6])
    defparam i10280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10281_3_lut (.I0(encoder0_position[12]), .I1(n2288), .I2(count_enable), 
            .I3(GND_net), .O(n23695));   // quad.v(35[10] 41[6])
    defparam i10281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1194_3_lut (.I0(n1761), .I1(n6785), .I2(n1778), .I3(GND_net), 
            .O(n1869));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10282_3_lut (.I0(encoder0_position[11]), .I1(n2289), .I2(count_enable), 
            .I3(GND_net), .O(n23696));   // quad.v(35[10] 41[6])
    defparam i10282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10283_3_lut (.I0(encoder0_position[10]), .I1(n2290), .I2(count_enable), 
            .I3(GND_net), .O(n23697));   // quad.v(35[10] 41[6])
    defparam i10283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10284_3_lut (.I0(encoder0_position[9]), .I1(n2291), .I2(count_enable), 
            .I3(GND_net), .O(n23698));   // quad.v(35[10] 41[6])
    defparam i10284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10285_3_lut (.I0(encoder0_position[8]), .I1(n2292), .I2(count_enable), 
            .I3(GND_net), .O(n23699));   // quad.v(35[10] 41[6])
    defparam i10285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10286_3_lut (.I0(encoder0_position[7]), .I1(n2293), .I2(count_enable), 
            .I3(GND_net), .O(n23700));   // quad.v(35[10] 41[6])
    defparam i10286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_i1265_3_lut (.I0(n1869), .I1(n6826), .I2(n1886), .I3(GND_net), 
            .O(n1974));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10287_3_lut (.I0(encoder0_position[6]), .I1(n2294), .I2(count_enable), 
            .I3(GND_net), .O(n23701));   // quad.v(35[10] 41[6])
    defparam i10287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10288_3_lut (.I0(encoder0_position[5]), .I1(n2295), .I2(count_enable), 
            .I3(GND_net), .O(n23702));   // quad.v(35[10] 41[6])
    defparam i10288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10289_3_lut (.I0(encoder0_position[4]), .I1(n2296), .I2(count_enable), 
            .I3(GND_net), .O(n23703));   // quad.v(35[10] 41[6])
    defparam i10289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4229));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10290_3_lut (.I0(encoder0_position[3]), .I1(n2297), .I2(count_enable), 
            .I3(GND_net), .O(n23704));   // quad.v(35[10] 41[6])
    defparam i10290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10291_3_lut (.I0(encoder0_position[2]), .I1(n2298), .I2(count_enable), 
            .I3(GND_net), .O(n23705));   // quad.v(35[10] 41[6])
    defparam i10291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10292_3_lut (.I0(encoder0_position[1]), .I1(n2299), .I2(count_enable), 
            .I3(GND_net), .O(n23706));   // quad.v(35[10] 41[6])
    defparam i10292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1428 (.I0(\FRAME_MATCHER.state_31__N_1861 [2]), .I1(n7_adj_4076), 
            .I2(n22303), .I3(n2857), .O(n6_adj_4438));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1428.LUT_INIT = 16'hcfce;
    SB_LUT4 div_11_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i3_4_lut_adj_1429 (.I0(n22296), .I1(n6_adj_4438), .I2(n16810), 
            .I3(n123), .O(n8_adj_4085));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_1429.LUT_INIT = 16'hdccc;
    SB_LUT4 i4_4_lut_adj_1430 (.I0(\FRAME_MATCHER.state_31__N_1861 [2]), .I1(n8_adj_4085), 
            .I2(n22309), .I3(n42425), .O(n49981));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1430.LUT_INIT = 16'hefcf;
    SB_LUT4 i1_3_lut (.I0(n2103), .I1(n89_adj_4033), .I2(n22424), .I3(GND_net), 
            .O(n42425));   // verilog/coms.v(126[12] 289[6])
    defparam i1_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i1_3_lut_adj_1431 (.I0(n3761), .I1(n42425), .I2(n22422), .I3(GND_net), 
            .O(n42428));   // verilog/coms.v(126[12] 289[6])
    defparam i1_3_lut_adj_1431.LUT_INIT = 16'hcdcd;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(n88), .I1(n22378), .I2(GND_net), .I3(GND_net), 
            .O(n22375));
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_3_lut_adj_1433 (.I0(n124), .I1(n42428), .I2(n63_adj_4075), 
            .I3(GND_net), .O(n7_adj_4439));   // verilog/coms.v(126[12] 289[6])
    defparam i1_3_lut_adj_1433.LUT_INIT = 16'h8c8c;
    SB_LUT4 i2_4_lut_adj_1434 (.I0(n7_adj_4439), .I1(n124), .I2(n22296), 
            .I3(n16810), .O(n6_adj_4430));   // verilog/coms.v(126[12] 289[6])
    defparam i2_4_lut_adj_1434.LUT_INIT = 16'haeaf;
    SB_LUT4 i3_4_lut_adj_1435 (.I0(n22309), .I1(n6_adj_4430), .I2(n22303), 
            .I3(\FRAME_MATCHER.state_31__N_1989 [1]), .O(n49980));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_1435.LUT_INIT = 16'hdfdd;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(n91), .I1(n22369), .I2(GND_net), .I3(GND_net), 
            .O(n22366));
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'hdddd;
    SB_LUT4 div_11_i1537_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6904), .I2(n2279_adj_4071), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10295_3_lut (.I0(\PID_CONTROLLER.err_prev [31]), .I1(\PID_CONTROLLER.err [31]), 
            .I2(n43357), .I3(GND_net), .O(n23709));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10295_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4112));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10296_3_lut (.I0(\PID_CONTROLLER.err_prev [23]), .I1(\PID_CONTROLLER.err [23]), 
            .I2(n43357), .I3(GND_net), .O(n23710));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10296_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10297_3_lut (.I0(\PID_CONTROLLER.err_prev [22]), .I1(\PID_CONTROLLER.err [22]), 
            .I2(n43357), .I3(GND_net), .O(n23711));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10297_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10298_3_lut (.I0(\PID_CONTROLLER.err_prev [21]), .I1(\PID_CONTROLLER.err [21]), 
            .I2(n43357), .I3(GND_net), .O(n23712));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10298_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10299_3_lut (.I0(\PID_CONTROLLER.err_prev [20]), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n43357), .I3(GND_net), .O(n23713));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10299_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10300_3_lut (.I0(\PID_CONTROLLER.err_prev [19]), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n43357), .I3(GND_net), .O(n23714));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10300_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10301_3_lut (.I0(\PID_CONTROLLER.err_prev [18]), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n43357), .I3(GND_net), .O(n23715));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10301_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1437 (.I0(n94), .I1(n22360), .I2(GND_net), .I3(GND_net), 
            .O(n22357));
    defparam i1_2_lut_adj_1437.LUT_INIT = 16'hdddd;
    SB_LUT4 i10302_3_lut (.I0(\PID_CONTROLLER.err_prev [17]), .I1(\PID_CONTROLLER.err [17]), 
            .I2(n43357), .I3(GND_net), .O(n23716));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10302_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10303_3_lut (.I0(\PID_CONTROLLER.err_prev [16]), .I1(\PID_CONTROLLER.err [16]), 
            .I2(n43357), .I3(GND_net), .O(n23717));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10303_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10304_3_lut (.I0(\PID_CONTROLLER.err_prev [15]), .I1(\PID_CONTROLLER.err [15]), 
            .I2(n43357), .I3(GND_net), .O(n23718));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10304_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10305_3_lut (.I0(\PID_CONTROLLER.err_prev [14]), .I1(\PID_CONTROLLER.err [14]), 
            .I2(n43357), .I3(GND_net), .O(n23719));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1438 (.I0(n224), .I1(n99), .I2(n22345), .I3(n558), 
            .O(n5_adj_4437));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i1_4_lut_adj_1438.LUT_INIT = 16'h555d;
    SB_LUT4 i10306_3_lut (.I0(\PID_CONTROLLER.err_prev [13]), .I1(\PID_CONTROLLER.err [13]), 
            .I2(n43357), .I3(GND_net), .O(n23720));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10307_3_lut (.I0(\PID_CONTROLLER.err_prev [12]), .I1(\PID_CONTROLLER.err [12]), 
            .I2(n43357), .I3(GND_net), .O(n23721));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10308_3_lut (.I0(\PID_CONTROLLER.err_prev [11]), .I1(\PID_CONTROLLER.err [11]), 
            .I2(n43357), .I3(GND_net), .O(n23722));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10309_3_lut (.I0(\PID_CONTROLLER.err_prev [10]), .I1(\PID_CONTROLLER.err [10]), 
            .I2(n43357), .I3(GND_net), .O(n23723));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31154_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n46620));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i31154_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i10310_3_lut (.I0(\PID_CONTROLLER.err_prev [9]), .I1(\PID_CONTROLLER.err [9]), 
            .I2(n43357), .I3(GND_net), .O(n23724));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10311_3_lut (.I0(\PID_CONTROLLER.err_prev [8]), .I1(\PID_CONTROLLER.err [8]), 
            .I2(n43357), .I3(GND_net), .O(n23725));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10312_3_lut (.I0(\PID_CONTROLLER.err_prev [7]), .I1(\PID_CONTROLLER.err [7]), 
            .I2(n43357), .I3(GND_net), .O(n23726));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1439 (.I0(n46620), .I1(n22345), .I2(n99), .I3(n5_adj_4437), 
            .O(n392));
    defparam i1_4_lut_adj_1439.LUT_INIT = 16'hefce;
    SB_LUT4 i10313_3_lut (.I0(\PID_CONTROLLER.err_prev [6]), .I1(\PID_CONTROLLER.err [6]), 
            .I2(n43357), .I3(GND_net), .O(n23727));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10314_3_lut (.I0(\PID_CONTROLLER.err_prev [5]), .I1(\PID_CONTROLLER.err [5]), 
            .I2(n43357), .I3(GND_net), .O(n23728));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4026), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10315_3_lut (.I0(\PID_CONTROLLER.err_prev [4]), .I1(\PID_CONTROLLER.err [4]), 
            .I2(n43357), .I3(GND_net), .O(n23729));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_297_i46_4_lut (.I0(n370), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i10316_3_lut (.I0(\PID_CONTROLLER.err_prev [3]), .I1(\PID_CONTROLLER.err [3]), 
            .I2(n43357), .I3(GND_net), .O(n23730));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10317_3_lut (.I0(\PID_CONTROLLER.err_prev [2]), .I1(\PID_CONTROLLER.err [2]), 
            .I2(n43357), .I3(GND_net), .O(n23731));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10318_3_lut (.I0(\PID_CONTROLLER.err_prev [1]), .I1(\PID_CONTROLLER.err [1]), 
            .I2(n43357), .I3(GND_net), .O(n23732));   // verilog/motorControl.v(38[14] 59[8])
    defparam i10318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1440 (.I0(n46), .I1(n22348), .I2(n98), .I3(n43086), 
            .O(n533));
    defparam i1_4_lut_adj_1440.LUT_INIT = 16'hefce;
    SB_LUT4 i21974_2_lut (.I0(n370), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4023));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i21974_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i31852_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n47413));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i31852_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i31786_3_lut (.I0(n369), .I1(n558), .I2(n392), .I3(GND_net), 
            .O(n510));
    defparam i31786_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_11_LessThan_1350_i20_4_lut (.I0(n383), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4236));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_i368_4_lut (.I0(n510), .I1(n2_adj_4023), .I2(n533), 
            .I3(n99), .O(n648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i368_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_LessThan_1350_i28_3_lut (.I0(n26_adj_4242), .I1(n93), 
            .I2(n31_adj_4246), .I3(GND_net), .O(n28_adj_4244));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31163_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n46722));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i31163_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4165));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4111));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4162));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31171_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n46730));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i31171_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4159));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31185_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n46744));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i31185_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4157));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1350_i32_3_lut (.I0(n24_adj_4240), .I1(n91), 
            .I2(n35_adj_4249), .I3(GND_net), .O(n32_adj_4247));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33328_4_lut (.I0(n32_adj_4247), .I1(n22_adj_4238), .I2(n35_adj_4249), 
            .I3(n47289), .O(n48889));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33328_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33329_3_lut (.I0(n48889), .I1(n90), .I2(n37_adj_4250), .I3(GND_net), 
            .O(n48890));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33329_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33153_3_lut (.I0(n48890), .I1(n89), .I2(n39_adj_4251), .I3(GND_net), 
            .O(n48714));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33153_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33063_4_lut (.I0(n39_adj_4251), .I1(n37_adj_4250), .I2(n35_adj_4249), 
            .I3(n47293), .O(n48624));
    defparam i33063_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_11_i367_4_lut (.I0(n43086), .I1(n4_adj_4022), .I2(n533), 
            .I3(n98), .O(n43088));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i367_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i33405_4_lut (.I0(n28_adj_4244), .I1(n20_adj_4236), .I2(n31_adj_4246), 
            .I3(n47295), .O(n48966));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33405_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i31189_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n46748));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i31189_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4110));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32164_3_lut (.I0(n48714), .I1(n88), .I2(n41_adj_4252), .I3(GND_net), 
            .O(n47725));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32164_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33482_4_lut (.I0(n47725), .I1(n48966), .I2(n41_adj_4252), 
            .I3(n48624), .O(n49043));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33482_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_adj_1441 (.I0(n96), .I1(n22354), .I2(GND_net), .I3(GND_net), 
            .O(n22351));
    defparam i1_2_lut_adj_1441.LUT_INIT = 16'hdddd;
    SB_LUT4 LessThan_542_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(GND_net), .O(n6_adj_4105));   // verilog/motorControl.v(86[28:44])
    defparam LessThan_542_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_11_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4109));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_390_i44_4_lut (.I0(n371), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i31203_3_lut_4_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(pwm_count[2]), .O(n46762));   // verilog/motorControl.v(86[28:44])
    defparam i31203_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32660_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n48221));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32660_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1442 (.I0(n48221), .I1(n22351), .I2(n97), .I3(n43088), 
            .O(n671));
    defparam i1_4_lut_adj_1442.LUT_INIT = 16'hefce;
    SB_LUT4 i10349_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n42422), .I3(GND_net), .O(n23763));   // verilog/coms.v(126[12] 289[6])
    defparam i10349_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10350_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n42422), .I3(GND_net), .O(n23764));   // verilog/coms.v(126[12] 289[6])
    defparam i10350_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10351_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n42422), .I3(GND_net), .O(n23765));   // verilog/coms.v(126[12] 289[6])
    defparam i10351_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10352_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n42422), .I3(GND_net), .O(n23766));   // verilog/coms.v(126[12] 289[6])
    defparam i10352_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10353_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n42422), .I3(GND_net), .O(n23767));   // verilog/coms.v(126[12] 289[6])
    defparam i10353_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22030_2_lut (.I0(n372), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4103));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i22030_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10354_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n42422), .I3(GND_net), .O(n23768));   // verilog/coms.v(126[12] 289[6])
    defparam i10354_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4156));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10355_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n42422), .I3(GND_net), .O(n23769));   // verilog/coms.v(126[12] 289[6])
    defparam i10355_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31778_3_lut (.I0(n371), .I1(n558), .I2(n671), .I3(GND_net), 
            .O(n785));
    defparam i31778_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i10356_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n42422), .I3(GND_net), .O(n23770));   // verilog/coms.v(126[12] 289[6])
    defparam i10356_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i550_4_lut (.I0(n785), .I1(n2_adj_4103), .I2(n806), 
            .I3(n99), .O(n917));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i550_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_11_i637_3_lut (.I0(n917), .I1(n5823), .I2(n938), .I3(GND_net), 
            .O(n1046));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i722_3_lut (.I0(n1046), .I1(n6215), .I2(n1067), .I3(GND_net), 
            .O(n1172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i805_3_lut (.I0(n1172), .I1(n6576), .I2(n1193), .I3(GND_net), 
            .O(n1295));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i805_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10365_3_lut (.I0(\data_in_frame[19] [7]), .I1(rx_data[7]), 
            .I2(n42421), .I3(GND_net), .O(n23779));   // verilog/coms.v(126[12] 289[6])
    defparam i10365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10366_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n42421), .I3(GND_net), .O(n23780));   // verilog/coms.v(126[12] 289[6])
    defparam i10366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4155));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4154));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10367_3_lut (.I0(\data_in_frame[19] [5]), .I1(rx_data[5]), 
            .I2(n42421), .I3(GND_net), .O(n23781));   // verilog/coms.v(126[12] 289[6])
    defparam i10367_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10368_3_lut (.I0(\data_in_frame[19] [4]), .I1(rx_data[4]), 
            .I2(n42421), .I3(GND_net), .O(n23782));   // verilog/coms.v(126[12] 289[6])
    defparam i10368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i886_3_lut (.I0(n1295), .I1(n6647), .I2(n1316), .I3(GND_net), 
            .O(n1415));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10369_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n42421), .I3(GND_net), .O(n23783));   // verilog/coms.v(126[12] 289[6])
    defparam i10369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10370_3_lut (.I0(\data_in_frame[19] [2]), .I1(rx_data[2]), 
            .I2(n42421), .I3(GND_net), .O(n23784));   // verilog/coms.v(126[12] 289[6])
    defparam i10370_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10371_3_lut (.I0(\data_in_frame[19] [1]), .I1(rx_data[1]), 
            .I2(n42421), .I3(GND_net), .O(n23785));   // verilog/coms.v(126[12] 289[6])
    defparam i10371_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4153));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4152));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10372_3_lut (.I0(\data_in_frame[19] [0]), .I1(rx_data[0]), 
            .I2(n42421), .I3(GND_net), .O(n23786));   // verilog/coms.v(126[12] 289[6])
    defparam i10372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i965_3_lut (.I0(n1415), .I1(n6687), .I2(n1436), .I3(GND_net), 
            .O(n1532));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i965_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4293));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31624_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n47185));
    defparam i31624_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4295));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4297));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31604_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n47165));
    defparam i31604_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4299));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4315));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31588_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n47149));
    defparam i31588_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4317));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4319));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31566_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n47127));
    defparam i31566_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4321));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4337));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31548_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n47109));
    defparam i31548_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4339));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4341));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31528_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n47089));
    defparam i31528_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4343));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4359));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4363));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31427_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n46987));
    defparam i31427_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4365));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4361));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31475_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n47035));
    defparam i31475_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4151));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4150));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4149));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4148));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4147));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4381));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4385));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31275_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n46834));
    defparam i31275_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4146));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4387));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4383));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31322_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n46881));
    defparam i31322_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4225));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_i1042_3_lut (.I0(n1532), .I1(n6727), .I2(n1553), .I3(GND_net), 
            .O(n1646));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4145));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n86), .I1(n85), .I2(n84), .I3(n22390), 
            .O(n22381));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i27624_2_lut_3_lut_4_lut (.I0(n22289), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n740), .O(n43181));
    defparam i27624_2_lut_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 div_11_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4144));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4143));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4142));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4141));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1117_3_lut (.I0(n1646), .I1(n6740), .I2(n1667), .I3(GND_net), 
            .O(n1757));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1190_3_lut (.I0(n1757), .I1(n6781), .I2(n1778), .I3(GND_net), 
            .O(n1865));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1261_3_lut (.I0(n1865), .I1(n6822), .I2(n1886), .I3(GND_net), 
            .O(n1970));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4140));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4234));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_481_i42_4_lut (.I0(n372), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n24202(n24202), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n24201(n24201), .n24200(n24200), .n24199(n24199), 
            .n24198(n24198), .n24197(n24197), .n24196(n24196), .n24195(n24195), 
            .n24194(n24194), .n24193(n24193), .n24192(n24192), .n24191(n24191), 
            .n24190(n24190), .n24189(n24189), .n24188(n24188), .n24187(n24187), 
            .n24186(n24186), .n24185(n24185), .n24184(n24184), .n24183(n24183), 
            .n24182(n24182), .n24181(n24181), .n24170(n24170), .data_o({quadA_debounced_adj_4057, 
            quadB_debounced_adj_4058}), .n2226({n2227, n2228, n2229, 
            n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
            n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
            n2246, n2247, n2248, n2249, n2250}), .GND_net(GND_net), 
            .n23577(n23577), .count_enable(count_enable_adj_4059), .n24231(n24231), 
            .reg_B({reg_B_adj_4485}), .n43884(n43884), .PIN_18_c_1(PIN_18_c_1), 
            .PIN_19_c_0(PIN_19_c_0), .n23580(n23580)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(174[15] 179[4])
    SB_LUT4 i33483_3_lut (.I0(n49043), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n49044));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33483_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_11_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4139));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4067));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1399_3_lut_3_lut (.I0(n2093), .I1(n6857), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1397_3_lut_3_lut (.I0(n2093), .I1(n6855), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4238));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33210_3_lut (.I0(n42), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n48771));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33210_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33211_3_lut (.I0(n48771), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n48772));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33211_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1443 (.I0(n48772), .I1(n22354), .I2(n96), .I3(n43090), 
            .O(n806));
    defparam i1_4_lut_adj_1443.LUT_INIT = 16'hefce;
    SB_LUT4 div_11_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i21982_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n370), .I3(n558), 
            .O(n4_adj_4022));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i21982_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_11_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4025), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n372));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31728_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n47289));
    defparam i31728_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i31766_3_lut (.I0(n372), .I1(n558), .I2(n806), .I3(GND_net), 
            .O(n918));
    defparam i31766_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_11_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4240));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31734_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n47295));
    defparam i31734_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4242));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_4_lut (.I0(n98), .I1(n97), .I2(n96), .I3(n22354), 
            .O(n22345));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1444 (.I0(n97), .I1(n96), .I2(n22354), 
            .I3(GND_net), .O(n22348));
    defparam i1_2_lut_3_lut_adj_1444.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1445 (.I0(n95), .I1(n94), .I2(n22360), 
            .I3(GND_net), .O(n22354));
    defparam i1_2_lut_3_lut_adj_1445.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_11_i638_3_lut (.I0(n918), .I1(n5824), .I2(n938), .I3(GND_net), 
            .O(n1047));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i638_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4138));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i723_3_lut (.I0(n1047), .I1(n6216), .I2(n1067), .I3(GND_net), 
            .O(n1173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1536_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6903), .I2(n2278_adj_4070), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1446 (.I0(n93), .I1(n92), .I2(n91), .I3(n22369), 
            .O(n22360));
    defparam i1_2_lut_4_lut_adj_1446.LUT_INIT = 16'hff7f;
    SB_LUT4 div_11_i806_3_lut (.I0(n1173), .I1(n6577), .I2(n1193), .I3(GND_net), 
            .O(n1296));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1447 (.I0(n92), .I1(n91), .I2(n22369), 
            .I3(GND_net), .O(n22363));
    defparam i1_2_lut_3_lut_adj_1447.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1448 (.I0(n90), .I1(n89), .I2(n88), .I3(n22378), 
            .O(n22369));
    defparam i1_2_lut_4_lut_adj_1448.LUT_INIT = 16'hff7f;
    SB_LUT4 div_11_i887_3_lut (.I0(n1296), .I1(n6648), .I2(n1316), .I3(GND_net), 
            .O(n1416));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10381_3_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(n42424), .I3(GND_net), .O(n23795));   // verilog/coms.v(126[12] 289[6])
    defparam i10381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10382_3_lut (.I0(\data_in_frame[17] [6]), .I1(rx_data[6]), 
            .I2(n42424), .I3(GND_net), .O(n23796));   // verilog/coms.v(126[12] 289[6])
    defparam i10382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i966_3_lut (.I0(n1416), .I1(n6688), .I2(n1436), .I3(GND_net), 
            .O(n1533));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i966_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1043_3_lut (.I0(n1533), .I1(n6728), .I2(n1553), .I3(GND_net), 
            .O(n1647));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10383_3_lut (.I0(\data_in_frame[17] [5]), .I1(rx_data[5]), 
            .I2(n42424), .I3(GND_net), .O(n23797));   // verilog/coms.v(126[12] 289[6])
    defparam i10383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10384_3_lut (.I0(\data_in_frame[17] [4]), .I1(rx_data[4]), 
            .I2(n42424), .I3(GND_net), .O(n23798));   // verilog/coms.v(126[12] 289[6])
    defparam i10384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10655_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24069));   // verilog/coms.v(126[12] 289[6])
    defparam i10655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10385_3_lut (.I0(\data_in_frame[17] [3]), .I1(rx_data[3]), 
            .I2(n42424), .I3(GND_net), .O(n23799));   // verilog/coms.v(126[12] 289[6])
    defparam i10385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10386_3_lut (.I0(\data_in_frame[17] [2]), .I1(rx_data[2]), 
            .I2(n42424), .I3(GND_net), .O(n23800));   // verilog/coms.v(126[12] 289[6])
    defparam i10386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10387_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n42424), .I3(GND_net), .O(n23801));   // verilog/coms.v(126[12] 289[6])
    defparam i10387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1396_3_lut_3_lut (.I0(n2093), .I1(n6854), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1449 (.I0(n89), .I1(n88), .I2(n22378), 
            .I3(GND_net), .O(n22372));
    defparam i1_2_lut_3_lut_adj_1449.LUT_INIT = 16'hf7f7;
    SB_LUT4 i10388_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(n42424), .I3(GND_net), .O(n23802));   // verilog/coms.v(126[12] 289[6])
    defparam i10388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1118_3_lut (.I0(n1647), .I1(n6741), .I2(n1667), .I3(GND_net), 
            .O(n1758));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1118_3_lut.LUT_INIT = 16'hacac;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    coms setpoint_23__I_0 (.clk32MHz(clk32MHz), .gearBoxRatio({gearBoxRatio}), 
         .GND_net(GND_net), .n24099(n24099), .\data_in[0] ({\data_in[0] }), 
         .n24098(n24098), .n24097(n24097), .n24096(n24096), .n24095(n24095), 
         .n24094(n24094), .n24093(n24093), .n24092(n24092), .\data_in[1] ({\data_in[1] }), 
         .n24091(n24091), .n24090(n24090), .n24089(n24089), .n24088(n24088), 
         .n24087(n24087), .n24086(n24086), .n24085(n24085), .n24084(n24084), 
         .\data_in[2] ({\data_in[2] }), .n24083(n24083), .n24082(n24082), 
         .n24081(n24081), .n24080(n24080), .n24079(n24079), .n24078(n24078), 
         .n24077(n24077), .deadband({deadband}), .n24258(n24258), .setpoint({setpoint}), 
         .n24257(n24257), .n24256(n24256), .n24255(n24255), .n24254(n24254), 
         .n24253(n24253), .n24252(n24252), .n24251(n24251), .n24250(n24250), 
         .n24249(n24249), .n24248(n24248), .n24247(n24247), .n24246(n24246), 
         .n24245(n24245), .n24244(n24244), .n24243(n24243), .n24242(n24242), 
         .n24241(n24241), .n24240(n24240), .n24239(n24239), .n24238(n24238), 
         .n24237(n24237), .n24236(n24236), .VCC_net(VCC_net), .IntegralLimit({IntegralLimit}), 
         .n24063(n24063), .\data_out_frame[5][2] (\data_out_frame[5] [2]), 
         .rx_data({rx_data}), .n24076(n24076), .\data_in[3] ({\data_in[3] }), 
         .n24075(n24075), .n24074(n24074), .n24073(n24073), .rx_data_ready(rx_data_ready), 
         .n24072(n24072), .\Kd[7] (Kd[7]), .n24071(n24071), .n23930(n23930), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .n23929(n23929), .n23928(n23928), 
         .n23927(n23927), .n23926(n23926), .n23925(n23925), .n23924(n23924), 
         .n23923(n23923), .n23914(n23914), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .n23913(n23913), .n23912(n23912), .n23911(n23911), .n23910(n23910), 
         .n23909(n23909), .n23908(n23908), .n23907(n23907), .\FRAME_MATCHER.state ({Open_0, 
         Open_1, Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, 
         Open_8, Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
         Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, Open_21, 
         Open_22, Open_23, Open_24, Open_25, Open_26, Open_27, Open_28, 
         Open_29, Open_30, \FRAME_MATCHER.state [0]}), .\FRAME_MATCHER.state[2] (\FRAME_MATCHER.state [2]), 
         .n23898(n23898), .\data_in_frame[5] ({\data_in_frame[5] }), .n23897(n23897), 
         .n23896(n23896), .n23895(n23895), .n23894(n23894), .n23893(n23893), 
         .n23892(n23892), .n23891(n23891), .\Kp[1] (Kp[1]), .\data_in_frame[6][1] (\data_in_frame[6] [1]), 
         .n23882(n23882), .\data_in_frame[7] ({\data_in_frame[7] }), .n23881(n23881), 
         .n23880(n23880), .n23879(n23879), .n23878(n23878), .n23877(n23877), 
         .n23876(n23876), .n23875(n23875), .\data_in_frame[8] ({Open_31, 
         Open_32, Open_33, Open_34, Open_35, Open_36, Open_37, \data_in_frame[8] [0]}), 
         .\data_in_frame[8][2] (\data_in_frame[8] [2]), .\Kp[2] (Kp[2]), 
         .n22501(n22501), .n2(n2_adj_4029), .n42614(n42614), .\Kp[3] (Kp[3]), 
         .\Kp[4] (Kp[4]), .n5(n5_adj_4028), .n23866(n23866), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .n43935(n43935), .\Kp[5] (Kp[5]), .n23865(n23865), .n42406(n42406), 
         .n23864(n23864), .n23863(n23863), .n23862(n23862), .n23861(n23861), 
         .n23860(n23860), .n23859(n23859), .\data_in_frame[12][4] (\data_in_frame[12] [4]), 
         .n23858(n23858), .\data_in_frame[10] ({\data_in_frame[10] }), .n23857(n23857), 
         .n23856(n23856), .n23855(n23855), .n23854(n23854), .n23853(n23853), 
         .n23852(n23852), .n23851(n23851), .n23850(n23850), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n23849(n23849), .\Kp[6] (Kp[6]), .n20435(n20435), .\data_in_frame[12][1] (\data_in_frame[12] [1]), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n42421(n42421), 
         .n23848(n23848), .n24070(n24070), .\Kp[7] (Kp[7]), .n22289(n22289), 
         .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .n23847(n23847), 
         .n22303(n22303), .n23846(n23846), .n28374(n28374), .n23844(n23844), 
         .n23843(n23843), .n63(n63_adj_4075), .n20088(n20088), .n23834(n23834), 
         .\data_in_frame[13] ({\data_in_frame[13] }), .n23833(n23833), .n23832(n23832), 
         .n23831(n23831), .n23830(n23830), .n26846(n26846), .n23828(n23828), 
         .n23827(n23827), .n23818(n23818), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .n124(n124), .n23817(n23817), .n23816(n23816), .n23815(n23815), 
         .n23814(n23814), .n23813(n23813), .n23812(n23812), .n23811(n23811), 
         .n2857(n2857), .n89(n89_adj_4033), .n22424(n22424), .n23802(n23802), 
         .\data_in_frame[17] ({\data_in_frame[17] }), .n23801(n23801), .n23800(n23800), 
         .n23799(n23799), .n24069(n24069), .n23798(n23798), .n23797(n23797), 
         .n23796(n23796), .n23795(n23795), .n23786(n23786), .\data_in_frame[19] ({\data_in_frame[19] }), 
         .n23785(n23785), .n23784(n23784), .n23783(n23783), .n23782(n23782), 
         .n23781(n23781), .n23780(n23780), .n23779(n23779), .n23770(n23770), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .n23769(n23769), .n23768(n23768), 
         .n23767(n23767), .n23766(n23766), .n23765(n23765), .n23764(n23764), 
         .n23763(n23763), .control_mode({control_mode}), .n20195(n20195), 
         .\Ki[4] (Ki[4]), .n42422(n42422), .n20420(n20420), .n43035(n43035), 
         .PWMLimit({PWMLimit}), .n49980(n49980), .n49981(n49981), .n43032(n43032), 
         .\Ki[5] (Ki[5]), .n43011(n43011), .n24068(n24068), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n24067(n24067), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n24066(n24066), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Kd[1] (Kd[1]), 
         .\Kd[2] (Kd[2]), .\Kd[3] (Kd[3]), .\Kd[4] (Kd[4]), .\Kd[5] (Kd[5]), 
         .\Kd[6] (Kd[6]), .LED_c(LED_c), .n22277(n22277), .encoder1_position({encoder1_position}), 
         .n38879(n38879), .n23013(n23013), .n22538(n22538), .n3346(n3346), 
         .encoder0_position({encoder0_position}), .n22589(n22589), .n23584(n23584), 
         .n41786(n41786), .n23570(n23570), .\Kd[0] (Kd[0]), .\Ki[0] (Ki[0]), 
         .\Kp[0] (Kp[0]), .n42896(n42896), .n42559(n42559), .n42920(n42920), 
         .displacement({displacement}), .n42621(n42621), .pwm({pwm}), 
         .n20471(n20471), .n42418(n42418), .n3790(n3790), .n407(n407), 
         .\PID_CONTROLLER.result[13] (\PID_CONTROLLER.result [13]), .n27(n27_adj_4088), 
         .n3791(n3791), .n3792(n3792), .n3793(n3793), .n3794(n3794), 
         .n5017(n5017), .n3795(n3795), .n3796(n3796), .n3797(n3797), 
         .n3798(n3798), .n3799(n3799), .r_SM_Main({r_SM_Main_adj_4476}), 
         .n3800(n3800), .n27_adj_3(n27), .n3801(n3801), .n27_adj_4(n27_adj_4081), 
         .n3802(n3802), .n3803(n3803), .\pwm_23__N_2960[13] (pwm_23__N_2960[13]), 
         .n50261(n50261), .n23444(n23444), .n3804(n3804), .n3805(n3805), 
         .n3806(n3806), .n123(n123), .n740(n740), .n16810(n16810), .\FRAME_MATCHER.state_31__N_1989[1] (\FRAME_MATCHER.state_31__N_1989 [1]), 
         .n3807(n3807), .n3808(n3808), .n3809(n3809), .n3810(n3810), 
         .n3811(n3811), .n3812(n3812), .n3813(n3813), .n22296(n22296), 
         .n22422(n22422), .n3761(n3761), .n2103(n2103), .n22309(n22309), 
         .\FRAME_MATCHER.state_31__N_1861[2] (\FRAME_MATCHER.state_31__N_1861 [2]), 
         .n7(n7_adj_4076), .n22908(n22908), .n42400(n42400), .n42424(n42424), 
         .n42405(n42405), .n42413(n42413), .n23609(n23609), .\r_Clock_Count[8] (r_Clock_Count_adj_4477[8]), 
         .n23612(n23612), .\r_Clock_Count[7] (r_Clock_Count_adj_4477[7]), 
         .n23615(n23615), .\r_Clock_Count[6] (r_Clock_Count_adj_4477[6]), 
         .n23618(n23618), .\r_Clock_Count[5] (r_Clock_Count_adj_4477[5]), 
         .n23621(n23621), .\r_Clock_Count[4] (r_Clock_Count_adj_4477[4]), 
         .n23624(n23624), .\r_Clock_Count[3] (r_Clock_Count_adj_4477[3]), 
         .n23627(n23627), .\r_Clock_Count[2] (r_Clock_Count_adj_4477[2]), 
         .n23630(n23630), .\r_Clock_Count[1] (r_Clock_Count_adj_4477[1]), 
         .n23634(n23634), .r_Bit_Index({r_Bit_Index_adj_4478}), .n23637(n23637), 
         .n24235(n24235), .n23680(n23680), .n313(n313), .n314(n314), 
         .n315(n315), .n316(n316), .n317(n317), .n318(n318), .\r_SM_Main_2__N_2753[1] (r_SM_Main_2__N_2753[1]), 
         .n319(n319), .n320(n320), .n23629(n23629), .n23463(n23463), 
         .n23547(n23547), .n4032(n4032), .o_Tx_Serial_N_2784(o_Tx_Serial_N_2784), 
         .n49982(n49982), .n23583(n23583), .n23581(n23581), .tx_o(tx_o), 
         .n49(n49), .tx_enable(tx_enable), .n23640(n23640), .r_Bit_Index_adj_12({r_Bit_Index}), 
         .n23643(n23643), .n28961(n28961), .\r_SM_Main[1]_adj_8 (r_SM_Main[1]), 
         .n23683(n23683), .n24171(n24171), .r_Rx_Data(r_Rx_Data), .PIN_13_N_26(PIN_13_N_26), 
         .n46671(n46671), .n46670(n46670), .\r_SM_Main[2]_adj_9 (r_SM_Main[2]), 
         .n23457(n23457), .n23545(n23545), .n4010(n4010), .n23650(n23650), 
         .n23649(n23649), .n23648(n23648), .n23647(n23647), .n23646(n23646), 
         .n23645(n23645), .n23644(n23644), .n23579(n23579), .n22411(n22411), 
         .n4(n4_adj_4030), .n28925(n28925), .n1(n1), .n28462(n28462), 
         .n4_adj_10(n4_adj_4055), .n4_adj_11(n4_adj_4054), .n22416(n22416)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(68[8] 88[4])
    SB_LUT4 div_11_i1191_3_lut (.I0(n1758), .I1(n6782), .I2(n1778), .I3(GND_net), 
            .O(n1866));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(n87), .I1(n86), .I2(n85), .I3(n22387), 
            .O(n22378));
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'hff7f;
    SB_LUT4 div_11_i1262_3_lut (.I0(n1866), .I1(n6823), .I2(n1886), .I3(GND_net), 
            .O(n1971));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4233));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4137));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10654_3_lut_4_lut (.I0(\data_out_frame[0] [2]), .I1(n3346), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23444), .O(n24068));   // verilog/coms.v(126[12] 289[6])
    defparam i10654_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 div_11_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4136));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4135));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4134));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4133));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10653_3_lut_4_lut (.I0(\data_out_frame[0] [3]), .I1(n3346), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23444), .O(n24067));   // verilog/coms.v(126[12] 289[6])
    defparam i10653_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i10397_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n42418), .I3(GND_net), .O(n23811));   // verilog/coms.v(126[12] 289[6])
    defparam i10397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10398_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n42418), .I3(GND_net), .O(n23812));   // verilog/coms.v(126[12] 289[6])
    defparam i10398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10399_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n42418), .I3(GND_net), .O(n23813));   // verilog/coms.v(126[12] 289[6])
    defparam i10399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10400_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n42418), .I3(GND_net), .O(n23814));   // verilog/coms.v(126[12] 289[6])
    defparam i10400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10401_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n42418), .I3(GND_net), .O(n23815));   // verilog/coms.v(126[12] 289[6])
    defparam i10401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10402_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n42418), .I3(GND_net), .O(n23816));   // verilog/coms.v(126[12] 289[6])
    defparam i10402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10403_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n42418), .I3(GND_net), .O(n23817));   // verilog/coms.v(126[12] 289[6])
    defparam i10403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10404_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n42418), .I3(GND_net), .O(n23818));   // verilog/coms.v(126[12] 289[6])
    defparam i10404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10652_3_lut_4_lut (.I0(\data_out_frame[0] [4]), .I1(n3346), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n23444), .O(n24066));   // verilog/coms.v(126[12] 289[6])
    defparam i10652_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i22038_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n372), .I3(n558), 
            .O(n4_adj_4102));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i22038_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i10413_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n20420), .I3(GND_net), .O(n23827));   // verilog/coms.v(126[12] 289[6])
    defparam i10413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10414_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n20420), .I3(GND_net), .O(n23828));   // verilog/coms.v(126[12] 289[6])
    defparam i10414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13447_3_lut (.I0(n20420), .I1(rx_data[5]), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n26846));   // verilog/coms.v(89[13:20])
    defparam i13447_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10416_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n20420), .I3(GND_net), .O(n23830));   // verilog/coms.v(126[12] 289[6])
    defparam i10416_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10417_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n20420), .I3(GND_net), .O(n23831));   // verilog/coms.v(126[12] 289[6])
    defparam i10417_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10418_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n20420), .I3(GND_net), .O(n23832));   // verilog/coms.v(126[12] 289[6])
    defparam i10418_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10419_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n20420), .I3(GND_net), .O(n23833));   // verilog/coms.v(126[12] 289[6])
    defparam i10419_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10420_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n20420), .I3(GND_net), .O(n23834));   // verilog/coms.v(126[12] 289[6])
    defparam i10420_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22006_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n371), .I3(n558), 
            .O(n4));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i22006_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(n85), .I1(n84), .I2(n22390), 
            .I3(GND_net), .O(n22384));
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1452 (.I0(n83), .I1(n82), .I2(n81), .I3(n22399), 
            .O(n22390));
    defparam i1_2_lut_4_lut_adj_1452.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1453 (.I0(n82), .I1(n81), .I2(n22399), 
            .I3(GND_net), .O(n22393));
    defparam i1_2_lut_3_lut_adj_1453.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1454 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n22399));
    defparam i1_2_lut_4_lut_adj_1454.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1455 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n22402));
    defparam i1_2_lut_3_lut_adj_1455.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_11_LessThan_570_i40_4_lut (.I0(n373), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_570_i44_3_lut (.I0(n42_adj_4157), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4158));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32662_4_lut (.I0(n44_adj_4158), .I1(n40), .I2(n45), .I3(n46748), 
            .O(n48223));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32662_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1456 (.I0(n48223), .I1(n22357), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1456.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n373));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_657_i38_4_lut (.I0(n374), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_657_i42_3_lut (.I0(n40_adj_4159), .I1(n96), 
            .I2(n43_adj_4161), .I3(GND_net), .O(n42_adj_4160));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33106_4_lut (.I0(n42_adj_4160), .I1(n38), .I2(n43_adj_4161), 
            .I3(n46744), .O(n48667));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33106_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33107_3_lut (.I0(n48667), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n48668));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33107_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1457 (.I0(n48668), .I1(n22360), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1457.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1395_3_lut_3_lut (.I0(n2093), .I1(n6853), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i639_3_lut (.I0(n373), .I1(n5825), .I2(n938), .I3(GND_net), 
            .O(n1048));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1398_3_lut_3_lut (.I0(n2093), .I1(n6856), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10429_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n20435), .I3(GND_net), .O(n23843));   // verilog/coms.v(126[12] 289[6])
    defparam i10429_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10430_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n20435), .I3(GND_net), .O(n23844));   // verilog/coms.v(126[12] 289[6])
    defparam i10430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14982_3_lut (.I0(n20435), .I1(rx_data[5]), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n28374));   // verilog/coms.v(89[13:20])
    defparam i14982_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10432_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n20435), .I3(GND_net), .O(n23846));   // verilog/coms.v(126[12] 289[6])
    defparam i10432_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10433_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n20435), .I3(GND_net), .O(n23847));   // verilog/coms.v(126[12] 289[6])
    defparam i10433_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_742_i36_4_lut (.I0(n375), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_11_LessThan_742_i40_3_lut (.I0(n38_adj_4162), .I1(n96), 
            .I2(n41_adj_4164), .I3(GND_net), .O(n40_adj_4163));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33403_4_lut (.I0(n40_adj_4163), .I1(n36), .I2(n41_adj_4164), 
            .I3(n46730), .O(n48964));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33403_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33438_3_lut (.I0(n49044), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n48999));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33438_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_11_i1394_3_lut_3_lut (.I0(n2093), .I1(n6852), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33404_3_lut (.I0(n48964), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n48965));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33404_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33303_3_lut (.I0(n48965), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n48864));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33303_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i10656_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24070));   // verilog/coms.v(126[12] 289[6])
    defparam i10656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1458 (.I0(n48864), .I1(n22363), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1458.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i724_3_lut (.I0(n1048), .I1(n6217), .I2(n1067), .I3(GND_net), 
            .O(n1174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10434_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n20435), .I3(GND_net), .O(n23848));   // verilog/coms.v(126[12] 289[6])
    defparam i10434_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10435_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n20435), .I3(GND_net), .O(n23849));   // verilog/coms.v(126[12] 289[6])
    defparam i10435_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10436_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n20435), .I3(GND_net), .O(n23850));   // verilog/coms.v(126[12] 289[6])
    defparam i10436_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10437_3_lut (.I0(\data_in_frame[10] [7]), .I1(rx_data[7]), 
            .I2(n42400), .I3(GND_net), .O(n23851));   // verilog/coms.v(126[12] 289[6])
    defparam i10437_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10438_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n42400), .I3(GND_net), .O(n23852));   // verilog/coms.v(126[12] 289[6])
    defparam i10438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10439_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n42400), .I3(GND_net), .O(n23853));   // verilog/coms.v(126[12] 289[6])
    defparam i10439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10440_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n42400), .I3(GND_net), .O(n23854));   // verilog/coms.v(126[12] 289[6])
    defparam i10440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10441_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n42400), .I3(GND_net), .O(n23855));   // verilog/coms.v(126[12] 289[6])
    defparam i10441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10442_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n42400), .I3(GND_net), .O(n23856));   // verilog/coms.v(126[12] 289[6])
    defparam i10442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10443_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n42400), .I3(GND_net), .O(n23857));   // verilog/coms.v(126[12] 289[6])
    defparam i10443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1471_3_lut_3_lut (.I0(n2192), .I1(n6882), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1459_3_lut_3_lut (.I0(n2192), .I1(n6870), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[7] [3]), 
            .I2(n2_adj_4029), .I3(n42614), .O(n42621));   // verilog/coms.v(94[12:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 div_11_i1470_3_lut_3_lut (.I0(n2192), .I1(n6881), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10444_3_lut (.I0(\data_in_frame[10] [0]), .I1(rx_data[0]), 
            .I2(n42400), .I3(GND_net), .O(n23858));   // verilog/coms.v(126[12] 289[6])
    defparam i10444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10445_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n42413), 
            .I3(GND_net), .O(n23859));   // verilog/coms.v(126[12] 289[6])
    defparam i10445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10446_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n42413), 
            .I3(GND_net), .O(n23860));   // verilog/coms.v(126[12] 289[6])
    defparam i10446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10447_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n42413), 
            .I3(GND_net), .O(n23861));   // verilog/coms.v(126[12] 289[6])
    defparam i10447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1467_3_lut_3_lut (.I0(n2192), .I1(n6878), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10448_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n42413), 
            .I3(GND_net), .O(n23862));   // verilog/coms.v(126[12] 289[6])
    defparam i10448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10449_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n42413), 
            .I3(GND_net), .O(n23863));   // verilog/coms.v(126[12] 289[6])
    defparam i10449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10450_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n42413), 
            .I3(GND_net), .O(n23864));   // verilog/coms.v(126[12] 289[6])
    defparam i10450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_i1465_3_lut_3_lut (.I0(n2192), .I1(n6876), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n7002), 
            .I3(n2724), .O(n41_adj_4427));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n7003), 
            .I3(n2724), .O(n39_adj_4425));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_i1475_3_lut_3_lut (.I0(n2192), .I1(n6886), .I2(n384), 
            .I3(GND_net), .O(n2280_adj_4072));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n391));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n7000), 
            .I3(n2724), .O(n45_adj_4429));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n7004), 
            .I3(n2724), .O(n37_adj_4424));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_i1463_3_lut_3_lut (.I0(n2192), .I1(n6874), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n7008), 
            .I3(n2724), .O(n29_adj_4419));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n7007), 
            .I3(n2724), .O(n31_adj_4421));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n7001), 
            .I3(n2724), .O(n43_adj_4428));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n7012), 
            .I3(n2724), .O(n21_adj_4414));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n7011), 
            .I3(n2724), .O(n23_adj_4415));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n7010), 
            .I3(n2724), .O(n25_adj_4417));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n7014), 
            .I3(n2724), .O(n17_adj_4412));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n7013), 
            .I3(n2724), .O(n19_adj_4413));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n7018), 
            .I3(n2724), .O(n9_adj_4405));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n7019), 
            .I3(n2724), .O(n7_adj_4403));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n7005), 
            .I3(n2724), .O(n35_adj_4423));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n7006), 
            .I3(n2724), .O(n33_adj_4422));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n7017), 
            .I3(n2724), .O(n11_adj_4407));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n7016), 
            .I3(n2724), .O(n13_adj_4409));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n7015), 
            .I3(n2724), .O(n15_adj_4410));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n7009), 
            .I3(n2724), .O(n27_adj_4418));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_11_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1462_3_lut_3_lut (.I0(n2192), .I1(n6873), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31183_4_lut (.I0(n27_adj_4418), .I1(n15_adj_4410), .I2(n13_adj_4409), 
            .I3(n11_adj_4407), .O(n46742));
    defparam i31183_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4422), 
            .I3(GND_net), .O(n12_adj_4408));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i31165_2_lut (.I0(n33_adj_4422), .I1(n15_adj_4410), .I2(GND_net), 
            .I3(GND_net), .O(n46724));
    defparam i31165_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_11_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4409), 
            .I3(GND_net), .O(n10_adj_4406));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1830_i30_3_lut (.I0(n12_adj_4408), .I1(n83), 
            .I2(n35_adj_4423), .I3(GND_net), .O(n30_adj_4420));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1828_3_lut (.I0(n2720), .I1(n7020), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31239_3_lut (.I0(n7_adj_4403), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n46798));
    defparam i31239_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i31988_4_lut (.I0(n13_adj_4409), .I1(n11_adj_4407), .I2(n9_adj_4405), 
            .I3(n46798), .O(n47549));
    defparam i31988_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i31978_4_lut (.I0(n19_adj_4413), .I1(n17_adj_4412), .I2(n15_adj_4410), 
            .I3(n47549), .O(n47539));
    defparam i31978_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33132_4_lut (.I0(n25_adj_4417), .I1(n23_adj_4415), .I2(n21_adj_4414), 
            .I3(n47539), .O(n48693));
    defparam i33132_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32590_4_lut (.I0(n31_adj_4421), .I1(n29_adj_4419), .I2(n27_adj_4418), 
            .I3(n48693), .O(n48151));
    defparam i32590_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33344_4_lut (.I0(n37_adj_4424), .I1(n35_adj_4423), .I2(n33_adj_4422), 
            .I3(n48151), .O(n48905));
    defparam i33344_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_11_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4428), 
            .I3(GND_net), .O(n16_adj_4411));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4403), 
            .I3(GND_net), .O(n6_adj_4402));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i33085_3_lut (.I0(n6_adj_4402), .I1(n90), .I2(n21_adj_4414), 
            .I3(GND_net), .O(n48646));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33085_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33086_3_lut (.I0(n48646), .I1(n89), .I2(n23_adj_4415), .I3(GND_net), 
            .O(n48647));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33086_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31205_4_lut (.I0(n21_adj_4414), .I1(n19_adj_4413), .I2(n17_adj_4412), 
            .I3(n9_adj_4405), .O(n46764));
    defparam i31205_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31918_2_lut (.I0(n43_adj_4428), .I1(n19_adj_4413), .I2(GND_net), 
            .I3(GND_net), .O(n47479));
    defparam i31918_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_11_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4412), 
            .I3(GND_net), .O(n8_adj_4404));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_11_LessThan_1830_i24_3_lut (.I0(n16_adj_4411), .I1(n78), 
            .I2(n45_adj_4429), .I3(GND_net), .O(n24_adj_4416));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31923_4_lut (.I0(n43_adj_4428), .I1(n25_adj_4417), .I2(n23_adj_4415), 
            .I3(n46764), .O(n47484));
    defparam i31923_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33015_4_lut (.I0(n24_adj_4416), .I1(n8_adj_4404), .I2(n45_adj_4429), 
            .I3(n47479), .O(n48576));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33015_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33010_3_lut (.I0(n48647), .I1(n88), .I2(n25_adj_4417), .I3(GND_net), 
            .O(n48571));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33010_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1829_3_lut (.I0(n390), .I1(n7021), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1830_i4_4_lut (.I0(n391), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4401));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33083_3_lut (.I0(n4_adj_4401), .I1(n87), .I2(n27_adj_4418), 
            .I3(GND_net), .O(n48644));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33083_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33084_3_lut (.I0(n48644), .I1(n86), .I2(n29_adj_4419), .I3(GND_net), 
            .O(n48645));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33084_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31173_4_lut (.I0(n33_adj_4422), .I1(n31_adj_4421), .I2(n29_adj_4419), 
            .I3(n46742), .O(n46732));
    defparam i31173_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33391_4_lut (.I0(n30_adj_4420), .I1(n10_adj_4406), .I2(n35_adj_4423), 
            .I3(n46724), .O(n48952));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33391_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33012_3_lut (.I0(n48645), .I1(n85), .I2(n31_adj_4421), .I3(GND_net), 
            .O(n48573));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33012_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33538_4_lut (.I0(n48573), .I1(n48952), .I2(n35_adj_4423), 
            .I3(n46732), .O(n49099));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33538_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33539_3_lut (.I0(n49099), .I1(n82), .I2(n37_adj_4424), .I3(GND_net), 
            .O(n49100));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33539_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1461_3_lut_3_lut (.I0(n2192), .I1(n6872), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33473_3_lut (.I0(n49100), .I1(n81), .I2(n39_adj_4425), .I3(GND_net), 
            .O(n49034));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33473_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31148_4_lut (.I0(n43_adj_4428), .I1(n41_adj_4427), .I2(n39_adj_4425), 
            .I3(n48905), .O(n46707));
    defparam i31148_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33369_4_lut (.I0(n48571), .I1(n48576), .I2(n45_adj_4429), 
            .I3(n47484), .O(n48930));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33369_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33453_3_lut (.I0(n49034), .I1(n80), .I2(n41_adj_4427), .I3(GND_net), 
            .O(n40_adj_4426));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33453_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1807_3_lut (.I0(n2699), .I1(n6999), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33371_4_lut (.I0(n40_adj_4426), .I1(n48930), .I2(n45_adj_4429), 
            .I3(n46707), .O(n48932));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33371_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33372_3_lut (.I0(n48932), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33372_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_11_i1464_3_lut_3_lut (.I0(n2192), .I1(n6875), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10451_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n42413), 
            .I3(GND_net), .O(n23865));   // verilog/coms.v(126[12] 289[6])
    defparam i10451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(\data_in_frame[10] [1]), .I3(\data_in_frame[7] [5]), .O(n43035));   // verilog/coms.v(94[12:25])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 div_11_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4398));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4400));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4396));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4399));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n390));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4393));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4394));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4391));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1460_3_lut_3_lut (.I0(n2192), .I1(n6871), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4392));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1474_3_lut_3_lut (.I0(n2192), .I1(n6885), .I2(n2183), 
            .I3(GND_net), .O(n2279_adj_4071));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4382));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4384));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4390));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4386));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4388));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4389));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4395));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31303_4_lut (.I0(n29_adj_4395), .I1(n17_adj_4389), .I2(n15_adj_4388), 
            .I3(n13_adj_4386), .O(n46862));
    defparam i31303_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32120_4_lut (.I0(n11_adj_4384), .I1(n9_adj_4382), .I2(n2719), 
            .I3(n98), .O(n47681));
    defparam i32120_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32644_4_lut (.I0(n17_adj_4389), .I1(n15_adj_4388), .I2(n13_adj_4386), 
            .I3(n47681), .O(n48205));
    defparam i32644_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_11_i1472_3_lut_3_lut (.I0(n2192), .I1(n6883), .I2(n2181), 
            .I3(GND_net), .O(n2277_adj_4069));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32636_4_lut (.I0(n23_adj_4392), .I1(n21_adj_4391), .I2(n19_adj_4390), 
            .I3(n48205), .O(n48197));
    defparam i32636_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31306_4_lut (.I0(n29_adj_4395), .I1(n27_adj_4394), .I2(n25_adj_4393), 
            .I3(n48197), .O(n46865));
    defparam i31306_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1777_i6_4_lut (.I0(n390), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4380));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33091_3_lut (.I0(n6_adj_4380), .I1(n87), .I2(n29_adj_4395), 
            .I3(GND_net), .O(n48652));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33091_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_i1473_3_lut_3_lut (.I0(n2192), .I1(n6884), .I2(n2182), 
            .I3(GND_net), .O(n2278_adj_4070));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1469_3_lut_3_lut (.I0(n2192), .I1(n6880), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1777_i32_3_lut (.I0(n14_adj_4387), .I1(n83), 
            .I2(n37_adj_4400), .I3(GND_net), .O(n32_adj_4397));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33092_3_lut (.I0(n48652), .I1(n86), .I2(n31_adj_4396), .I3(GND_net), 
            .O(n48653));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33092_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31285_4_lut (.I0(n35_adj_4399), .I1(n33_adj_4398), .I2(n31_adj_4396), 
            .I3(n46862), .O(n46844));
    defparam i31285_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33409_4_lut (.I0(n32_adj_4397), .I1(n12_adj_4385), .I2(n37_adj_4400), 
            .I3(n46834), .O(n48970));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33409_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33002_3_lut (.I0(n48653), .I1(n85), .I2(n33_adj_4398), .I3(GND_net), 
            .O(n48563));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33002_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33093_3_lut (.I0(n8_adj_4381), .I1(n90), .I2(n23_adj_4392), 
            .I3(GND_net), .O(n48654));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33093_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33094_3_lut (.I0(n48654), .I1(n89), .I2(n25_adj_4393), .I3(GND_net), 
            .O(n48655));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33094_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32050_4_lut (.I0(n25_adj_4393), .I1(n23_adj_4392), .I2(n21_adj_4391), 
            .I3(n46881), .O(n47611));
    defparam i32050_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32999_3_lut (.I0(n10_adj_4383), .I1(n91), .I2(n21_adj_4391), 
            .I3(GND_net), .O(n48560));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32999_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32998_3_lut (.I0(n48655), .I1(n88), .I2(n27_adj_4394), .I3(GND_net), 
            .O(n48559));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32998_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32892_4_lut (.I0(n35_adj_4399), .I1(n33_adj_4398), .I2(n31_adj_4396), 
            .I3(n46865), .O(n48453));
    defparam i32892_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33536_4_lut (.I0(n48563), .I1(n48970), .I2(n37_adj_4400), 
            .I3(n46844), .O(n49097));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33536_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33087_4_lut (.I0(n48559), .I1(n48560), .I2(n27_adj_4394), 
            .I3(n47611), .O(n48648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33087_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_11_i1468_3_lut_3_lut (.I0(n2192), .I1(n6879), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33558_4_lut (.I0(n48648), .I1(n49097), .I2(n37_adj_4400), 
            .I3(n48453), .O(n49119));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33558_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33559_3_lut (.I0(n49119), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n49120));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33559_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33555_3_lut (.I0(n49120), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n49116));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33555_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33342_3_lut (.I0(n49116), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n48903));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33342_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33343_3_lut (.I0(n48903), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n48904));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33343_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1804_4_lut (.I0(n48904), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1804_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4377));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1466_3_lut_3_lut (.I0(n2192), .I1(n6877), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4379));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4375));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n389));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4372));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4373));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4378));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1533_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6900), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4360));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22345), 
            .O(n249));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 div_11_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4362));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4364));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4366));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4367));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31448_4_lut (.I0(n31_adj_4374), .I1(n19_adj_4367), .I2(n17_adj_4366), 
            .I3(n15_adj_4364), .O(n47008));
    defparam i31448_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32255_4_lut (.I0(n13_adj_4362), .I1(n11_adj_4360), .I2(n2637), 
            .I3(n98), .O(n47816));
    defparam i32255_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32690_4_lut (.I0(n19_adj_4367), .I1(n17_adj_4366), .I2(n15_adj_4364), 
            .I3(n47816), .O(n48251));
    defparam i32690_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_11_i1522_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6889), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32686_4_lut (.I0(n25_adj_4371), .I1(n23_adj_4370), .I2(n21_adj_4369), 
            .I3(n48251), .O(n48247));
    defparam i32686_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31452_4_lut (.I0(n31_adj_4374), .I1(n29_adj_4373), .I2(n27_adj_4372), 
            .I3(n48247), .O(n47012));
    defparam i31452_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1722_i8_4_lut (.I0(n389), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4358));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32836_3_lut (.I0(n8_adj_4358), .I1(n87), .I2(n31_adj_4374), 
            .I3(GND_net), .O(n48397));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32836_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32837_3_lut (.I0(n48397), .I1(n86), .I2(n33_adj_4375), .I3(GND_net), 
            .O(n48398));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32837_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1722_i34_3_lut (.I0(n16_adj_4365), .I1(n83), 
            .I2(n39_adj_4379), .I3(GND_net), .O(n34_adj_4376));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31437_4_lut (.I0(n37_adj_4378), .I1(n35_adj_4377), .I2(n33_adj_4375), 
            .I3(n47008), .O(n46997));
    defparam i31437_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33407_4_lut (.I0(n34_adj_4376), .I1(n14_adj_4363), .I2(n39_adj_4379), 
            .I3(n46987), .O(n48968));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33407_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32212_3_lut (.I0(n48398), .I1(n85), .I2(n35_adj_4377), .I3(GND_net), 
            .O(n47773));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32212_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32838_3_lut (.I0(n10_adj_4359), .I1(n90), .I2(n25_adj_4371), 
            .I3(GND_net), .O(n48399));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32838_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32839_3_lut (.I0(n48399), .I1(n89), .I2(n27_adj_4372), .I3(GND_net), 
            .O(n48400));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32839_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32237_4_lut (.I0(n27_adj_4372), .I1(n25_adj_4371), .I2(n23_adj_4370), 
            .I3(n47035), .O(n47798));
    defparam i32237_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_11_LessThan_1722_i20_3_lut (.I0(n12_adj_4361), .I1(n91), 
            .I2(n23_adj_4370), .I3(GND_net), .O(n20_adj_4368));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32210_3_lut (.I0(n48400), .I1(n88), .I2(n29_adj_4373), .I3(GND_net), 
            .O(n47771));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32210_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33017_4_lut (.I0(n37_adj_4378), .I1(n35_adj_4377), .I2(n33_adj_4375), 
            .I3(n47012), .O(n48578));
    defparam i33017_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33534_4_lut (.I0(n47773), .I1(n48968), .I2(n39_adj_4379), 
            .I3(n46997), .O(n49095));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33534_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32993_4_lut (.I0(n47771), .I1(n20_adj_4368), .I2(n29_adj_4373), 
            .I3(n47798), .O(n48554));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32993_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33560_4_lut (.I0(n48554), .I1(n49095), .I2(n39_adj_4379), 
            .I3(n48578), .O(n49121));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33560_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i31220_3_lut_4_lut (.I0(pwm_count[3]), .I1(pwm[3]), .I2(pwm[2]), 
            .I3(pwm_count[2]), .O(n46779));   // verilog/motorControl.v(65[19:32])
    defparam i31220_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_539_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(pwm[3]), 
            .I2(pwm[2]), .I3(GND_net), .O(n6_adj_4093));   // verilog/motorControl.v(65[19:32])
    defparam LessThan_539_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i33561_3_lut (.I0(n49121), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n49122));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33561_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33553_3_lut (.I0(n49122), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n49114));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33553_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i32995_3_lut (.I0(n49114), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n48556));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32995_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1459 (.I0(n48556), .I1(n22405), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1459.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4355));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4357));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1525_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6892), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4353));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n388));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4356));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4350));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4351));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4347));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4348));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4349));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4342));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4344));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4345));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4352));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4338));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4340));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31536_4_lut (.I0(n33_adj_4352), .I1(n21_adj_4345), .I2(n19_adj_4344), 
            .I3(n17_adj_4342), .O(n47097));
    defparam i31536_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32297_4_lut (.I0(n15_adj_4340), .I1(n13_adj_4338), .I2(n2552), 
            .I3(n98), .O(n47858));
    defparam i32297_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32710_4_lut (.I0(n21_adj_4345), .I1(n19_adj_4344), .I2(n17_adj_4342), 
            .I3(n47858), .O(n48271));
    defparam i32710_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32708_4_lut (.I0(n27_adj_4349), .I1(n25_adj_4348), .I2(n23_adj_4347), 
            .I3(n48271), .O(n48269));
    defparam i32708_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31538_4_lut (.I0(n33_adj_4352), .I1(n31_adj_4351), .I2(n29_adj_4350), 
            .I3(n48269), .O(n47099));
    defparam i31538_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1665_i10_4_lut (.I0(n388), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4336));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32844_3_lut (.I0(n10_adj_4336), .I1(n87), .I2(n33_adj_4352), 
            .I3(GND_net), .O(n48405));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32844_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_4_lut_adj_1460 (.I0(n48999), .I1(n22387), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1460.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_i1523_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6890), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32845_3_lut (.I0(n48405), .I1(n86), .I2(n35_adj_4353), .I3(GND_net), 
            .O(n48406));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32845_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_825_i34_4_lut (.I0(n376), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33102_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4167), .I3(GND_net), 
            .O(n48663));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33102_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1665_i36_3_lut (.I0(n18_adj_4343), .I1(n83), 
            .I2(n41_adj_4357), .I3(GND_net), .O(n36_adj_4354));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31532_4_lut (.I0(n39_adj_4356), .I1(n37_adj_4355), .I2(n35_adj_4353), 
            .I3(n47097), .O(n47093));
    defparam i31532_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33340_4_lut (.I0(n36_adj_4354), .I1(n16_adj_4341), .I2(n41_adj_4357), 
            .I3(n47089), .O(n48901));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33340_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33103_3_lut (.I0(n48663), .I1(n94), .I2(n43_adj_4168), .I3(GND_net), 
            .O(n48664));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33103_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31934_4_lut (.I0(n43_adj_4168), .I1(n41_adj_4167), .I2(n39), 
            .I3(n46722), .O(n47495));
    defparam i31934_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32200_3_lut (.I0(n48406), .I1(n85), .I2(n37_adj_4355), .I3(GND_net), 
            .O(n47761));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32200_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_825_i38_3_lut (.I0(n36_adj_4165), .I1(n96), 
            .I2(n39), .I3(GND_net), .O(n38_adj_4166));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32963_3_lut (.I0(n48664), .I1(n93), .I2(n45_adj_4170), .I3(GND_net), 
            .O(n44_adj_4169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32963_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32666_4_lut (.I0(n44_adj_4169), .I1(n38_adj_4166), .I2(n45_adj_4170), 
            .I3(n47495), .O(n48227));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32666_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_11_LessThan_1665_i22_3_lut (.I0(n14_adj_4339), .I1(n91), 
            .I2(n25_adj_4348), .I3(GND_net), .O(n22_adj_4346));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33338_4_lut (.I0(n22_adj_4346), .I1(n12_adj_4337), .I2(n25_adj_4348), 
            .I3(n47109), .O(n48899));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33338_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33339_3_lut (.I0(n48899), .I1(n90), .I2(n27_adj_4349), .I3(GND_net), 
            .O(n48900));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33339_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33137_3_lut (.I0(n48900), .I1(n89), .I2(n29_adj_4350), .I3(GND_net), 
            .O(n48698));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33137_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33029_4_lut (.I0(n39_adj_4356), .I1(n37_adj_4355), .I2(n35_adj_4353), 
            .I3(n47099), .O(n48590));
    defparam i33029_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33496_4_lut (.I0(n47761), .I1(n48901), .I2(n41_adj_4357), 
            .I3(n47093), .O(n49057));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33496_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32198_3_lut (.I0(n48698), .I1(n88), .I2(n31_adj_4351), .I3(GND_net), 
            .O(n47759));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32198_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33564_4_lut (.I0(n47759), .I1(n49057), .I2(n41_adj_4357), 
            .I3(n48590), .O(n49125));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33564_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33565_3_lut (.I0(n49125), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n49126));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33565_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33557_3_lut (.I0(n49126), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n49118));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33557_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1461 (.I0(n49118), .I1(n22402), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1461.LUT_INIT = 16'hceef;
    SB_LUT4 i10452_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n42413), 
            .I3(GND_net), .O(n23866));   // verilog/coms.v(126[12] 289[6])
    defparam i10452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4221));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31754_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n47315));
    defparam i31754_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4333));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4223));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4331));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31760_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n47321));
    defparam i31760_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4335));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4334));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n387_adj_4068));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31791_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n47352));
    defparam i31791_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4211));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4328));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4329));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4207));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31782_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n47343));
    defparam i31782_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4209));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4325));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4326));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4327));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4195));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31805_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n47366));
    defparam i31805_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4197));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4316));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4318));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4184));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31820_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n47381));
    defparam i31820_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4186));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4320));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4322));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4323));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4330));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31576_4_lut (.I0(n35_adj_4330), .I1(n23_adj_4323), .I2(n21_adj_4322), 
            .I3(n19_adj_4320), .O(n47137));
    defparam i31576_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32333_4_lut (.I0(n17_adj_4318), .I1(n15_adj_4316), .I2(n2464), 
            .I3(n98), .O(n47894));
    defparam i32333_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32730_4_lut (.I0(n23_adj_4323), .I1(n21_adj_4322), .I2(n19_adj_4320), 
            .I3(n47894), .O(n48291));
    defparam i32730_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32726_4_lut (.I0(n29_adj_4327), .I1(n27_adj_4326), .I2(n25_adj_4325), 
            .I3(n48291), .O(n48287));
    defparam i32726_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31580_4_lut (.I0(n35_adj_4330), .I1(n33_adj_4329), .I2(n31_adj_4328), 
            .I3(n48287), .O(n47141));
    defparam i31580_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_LessThan_1606_i12_4_lut (.I0(n387_adj_4068), .I1(n99), 
            .I2(n2465), .I3(n558), .O(n12_adj_4314));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32848_3_lut (.I0(n12_adj_4314), .I1(n87), .I2(n35_adj_4330), 
            .I3(GND_net), .O(n48409));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32848_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4123));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1526_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6893), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1535_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6902), .I2(n2277_adj_4069), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1606_i38_3_lut (.I0(n20_adj_4321), .I1(n83), 
            .I2(n43_adj_4335), .I3(GND_net), .O(n38_adj_4332));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32849_3_lut (.I0(n48409), .I1(n86), .I2(n37_adj_4331), .I3(GND_net), 
            .O(n48410));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32849_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31570_4_lut (.I0(n41_adj_4334), .I1(n39_adj_4333), .I2(n37_adj_4331), 
            .I3(n47137), .O(n47131));
    defparam i31570_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33294_4_lut (.I0(n38_adj_4332), .I1(n18_adj_4319), .I2(n43_adj_4335), 
            .I3(n47127), .O(n48855));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33294_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32194_3_lut (.I0(n48410), .I1(n85), .I2(n39_adj_4333), .I3(GND_net), 
            .O(n47755));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32194_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1606_i24_3_lut (.I0(n16_adj_4317), .I1(n91), 
            .I2(n27_adj_4326), .I3(GND_net), .O(n24_adj_4324));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33336_4_lut (.I0(n24_adj_4324), .I1(n14_adj_4315), .I2(n27_adj_4326), 
            .I3(n47149), .O(n48897));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33336_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33337_3_lut (.I0(n48897), .I1(n90), .I2(n29_adj_4327), .I3(GND_net), 
            .O(n48898));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33337_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33139_3_lut (.I0(n48898), .I1(n89), .I2(n31_adj_4328), .I3(GND_net), 
            .O(n48700));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33139_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33041_4_lut (.I0(n41_adj_4334), .I1(n39_adj_4333), .I2(n37_adj_4331), 
            .I3(n47141), .O(n48602));
    defparam i33041_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33478_4_lut (.I0(n47755), .I1(n48855), .I2(n43_adj_4335), 
            .I3(n47131), .O(n49039));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33478_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32192_3_lut (.I0(n48700), .I1(n88), .I2(n33_adj_4329), .I3(GND_net), 
            .O(n47753));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32192_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33544_4_lut (.I0(n47753), .I1(n49039), .I2(n43_adj_4335), 
            .I3(n48602), .O(n49105));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33544_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33545_3_lut (.I0(n49105), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n49106));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33545_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1462 (.I0(n49106), .I1(n22399), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1462.LUT_INIT = 16'hceef;
    SB_LUT4 div_11_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31834_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n47395));
    defparam i31834_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4176));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4311));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n2276({n2277, n2278, n2279, 
            n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
            n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
            n2296, n2297, n2298, n2299, n2300}), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .data_o({quadA_debounced, quadB_debounced}), 
            .clk32MHz(clk32MHz), .n23706(n23706), .n23705(n23705), .n23704(n23704), 
            .n23703(n23703), .n23702(n23702), .n23701(n23701), .n23700(n23700), 
            .n23699(n23699), .n23698(n23698), .n23697(n23697), .n23696(n23696), 
            .n23695(n23695), .n23694(n23694), .n23693(n23693), .n23692(n23692), 
            .n23691(n23691), .n23690(n23690), .n23689(n23689), .n23688(n23688), 
            .n23687(n23687), .n23686(n23686), .n23685(n23685), .n23684(n23684), 
            .n23576(n23576), .count_enable(count_enable), .n24227(n24227), 
            .reg_B({reg_B}), .n44196(n44196), .PIN_23_c_1(PIN_23_c_1), 
            .PIN_24_c_0(PIN_24_c_0), .n23578(n23578)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(166[15] 171[4])
    SB_LUT4 div_11_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4313));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4309));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10821_3_lut_4_lut (.I0(r_SM_Main_adj_4476[2]), .I1(r_SM_Main_2__N_2753[1]), 
            .I2(r_SM_Main_adj_4476[0]), .I3(r_SM_Main_adj_4476[1]), .O(n24235));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10821_3_lut_4_lut.LUT_INIT = 16'h1540;
    SB_LUT4 div_11_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n386));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_11_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4255));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4312));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31698_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n47259));
    defparam i31698_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4306));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4307));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4257));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4259));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31704_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n47265));
    defparam i31704_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4303));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4304));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4305));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278_adj_4070), 
            .I3(GND_net), .O(n18_adj_4275));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31660_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277_adj_4069), 
            .I3(n96), .O(n47221));
    defparam i31660_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4277));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_11_i1595_3_lut_3_lut (.I0(n2381), .I1(n6921), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4294));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1333_3_lut (.I0(n1973), .I1(n6841), .I2(n1991), .I3(GND_net), 
            .O(n2075));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1333_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_11_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4122));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4296));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4279));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31670_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n47231));
    defparam i31670_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_11_i1583_3_lut_3_lut (.I0(n2381), .I1(n6909), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1584_3_lut_3_lut (.I0(n2381), .I1(n6910), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4298));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1587_3_lut_3_lut (.I0(n2381), .I1(n6913), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4300));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4301));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4308));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_11_i1588_3_lut_3_lut (.I0(n2381), .I1(n6914), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1585_3_lut_3_lut (.I0(n2381), .I1(n6911), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_11_i1532_3_lut_3_lut (.I0(n2288_adj_4073), .I1(n6899), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31614_4_lut (.I0(n37_adj_4308), .I1(n25_adj_4301), .I2(n23_adj_4300), 
            .I3(n21_adj_4298), .O(n47175));
    defparam i31614_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32371_4_lut (.I0(n19_adj_4296), .I1(n17_adj_4294), .I2(n2373), 
            .I3(n98), .O(n47932));
    defparam i32371_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i32748_4_lut (.I0(n25_adj_4301), .I1(n23_adj_4300), .I2(n21_adj_4298), 
            .I3(n47932), .O(n48309));
    defparam i32748_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_11_i1586_3_lut_3_lut (.I0(n2381), .I1(n6912), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32746_4_lut (.I0(n31_adj_4305), .I1(n29_adj_4304), .I2(n27_adj_4303), 
            .I3(n48309), .O(n48307));
    defparam i32746_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31616_4_lut (.I0(n37_adj_4308), .I1(n35_adj_4307), .I2(n33_adj_4306), 
            .I3(n48307), .O(n47177));
    defparam i31616_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_11_i1601_3_lut_3_lut (.I0(n2381), .I1(n6927), .I2(n386), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_11_LessThan_1545_i14_4_lut (.I0(n386), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4292));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i32854_3_lut (.I0(n14_adj_4292), .I1(n87), .I2(n37_adj_4308), 
            .I3(GND_net), .O(n48415));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32854_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32855_3_lut (.I0(n48415), .I1(n86), .I2(n39_adj_4309), .I3(GND_net), 
            .O(n48416));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32855_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1545_i40_3_lut (.I0(n22_adj_4299), .I1(n83), 
            .I2(n45_adj_4313), .I3(GND_net), .O(n40_adj_4310));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31608_4_lut (.I0(n43_adj_4312), .I1(n41_adj_4311), .I2(n39_adj_4309), 
            .I3(n47175), .O(n47169));
    defparam i31608_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32987_4_lut (.I0(n40_adj_4310), .I1(n20_adj_4297), .I2(n45_adj_4313), 
            .I3(n47165), .O(n48548));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32987_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32186_3_lut (.I0(n48416), .I1(n85), .I2(n41_adj_4311), .I3(GND_net), 
            .O(n47747));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32186_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_11_LessThan_1545_i26_3_lut (.I0(n18_adj_4295), .I1(n91), 
            .I2(n29_adj_4304), .I3(GND_net), .O(n26_adj_4302));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_11_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33334_4_lut (.I0(n26_adj_4302), .I1(n16_adj_4293), .I2(n29_adj_4304), 
            .I3(n47185), .O(n48895));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33334_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33335_3_lut (.I0(n48895), .I1(n90), .I2(n31_adj_4305), .I3(GND_net), 
            .O(n48896));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33335_3_lut.LUT_INIT = 16'h3a3a;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, deadband, \PID_CONTROLLER.result[13] , n459, 
            n460, \PID_CONTROLLER.err[9] , n461, \PID_CONTROLLER.err[8] , 
            \PID_CONTROLLER.err[7] , n462, \PID_CONTROLLER.err[6] , n463, 
            \PID_CONTROLLER.err[5] , \PID_CONTROLLER.result[7] , n465, 
            \PID_CONTROLLER.err[4] , \PID_CONTROLLER.err[3] , \PID_CONTROLLER.err[2] , 
            \PID_CONTROLLER.err[1] , \PID_CONTROLLER.err[0] , pwm_count, 
            \pwm_23__N_2960[13] , VCC_net, \PID_CONTROLLER.result[5] , 
            \pwm_23__N_2960[14] , \PID_CONTROLLER.result[14] , n467, n468, 
            n469, n470, n50246, \PID_CONTROLLER.result[21] , \pwm_23__N_2960[20] , 
            \PID_CONTROLLER.result[20] , n27, n29, n471, \motor_state[23] , 
            \motor_state[22] , \motor_state[21] , \motor_state[20] , \motor_state[19] , 
            \motor_state[18] , \motor_state[17] , n41, pwm_23__N_2957, 
            \motor_state[16] , n399, n24225, pwm, clk32MHz, n24224, 
            n24221, n24220, n24219, n24218, n24217, n24214, n24213, 
            n24212, n24211, n24210, n24208, n24206, n24205, n24204, 
            n24203, n24172, n400, \motor_state[15] , PIN_7_c_1, \motor_state[14] , 
            PIN_6_c_0, \motor_state[13] , \motor_state[12] , \motor_state[11] , 
            \motor_state[10] , \motor_state[9] , \motor_state[8] , \motor_state[7] , 
            \motor_state[6] , \motor_state[5] , \motor_state[4] , \motor_state[3] , 
            \motor_state[2] , n406, \motor_state[1] , n407, \motor_state[0] , 
            \PID_CONTROLLER.err_prev[31] , \PID_CONTROLLER.err_prev[23] , 
            \PID_CONTROLLER.err_prev[22] , \PID_CONTROLLER.err_prev[21] , 
            \PID_CONTROLLER.err_prev[20] , \PID_CONTROLLER.err_prev[19] , 
            \PID_CONTROLLER.err_prev[18] , \PID_CONTROLLER.err_prev[17] , 
            \PID_CONTROLLER.err_prev[16] , n413, \PID_CONTROLLER.err_prev[15] , 
            \PID_CONTROLLER.err_prev[14] , \PID_CONTROLLER.err_prev[13] , 
            \PID_CONTROLLER.err_prev[12] , \PID_CONTROLLER.err_prev[11] , 
            \Kd[4] , \Kp[7] , \PID_CONTROLLER.err[17] , n415, \PID_CONTROLLER.err_prev[10] , 
            \PID_CONTROLLER.err_prev[9] , \PID_CONTROLLER.err_prev[8] , 
            \PID_CONTROLLER.err_prev[7] , \PID_CONTROLLER.err[31] , \PID_CONTROLLER.err_prev[6] , 
            \Kp[1] , \PID_CONTROLLER.err[20] , \Kp[0] , \PID_CONTROLLER.err[21] , 
            \PID_CONTROLLER.err_prev[5] , \Kd[0] , \Kd[1] , \Kd[2] , 
            \PID_CONTROLLER.err_prev[4] , \PID_CONTROLLER.err_prev[3] , 
            \Kp[2] , \Kd[5] , \Kp[3] , hall1, hall2, \Kp[4] , \PID_CONTROLLER.err[10] , 
            \Kp[5] , \PID_CONTROLLER.err_prev[2] , \PID_CONTROLLER.err_prev[1] , 
            \PID_CONTROLLER.err_prev[0] , \Kp[6] , \PID_CONTROLLER.err[11] , 
            n853, n21, n855, n856, n857, n859, n860, n861, n862, 
            n863, n864, n865, n866, \PID_CONTROLLER.err[12] , PWMLimit, 
            setpoint, \Kd[6] , \PID_CONTROLLER.err[16] , n867, \PID_CONTROLLER.err[13] , 
            n868, n869, \Ki[3] , \Kd[7] , \Ki[7] , \Kd[3] , n870, 
            n871, n872, n873, n874, n875, \PID_CONTROLLER.err[15] , 
            n46619, \Ki[4] , \Ki[5] , \Ki[6] , \PID_CONTROLLER.err[14] , 
            \Ki[1] , \Ki[0] , \PID_CONTROLLER.err[18] , \PID_CONTROLLER.err[19] , 
            \Ki[2] , \PID_CONTROLLER.err[22] , n448, n449, \PID_CONTROLLER.err[23] , 
            n23732, n23731, n23730, n23729, n23728, n23727, n23726, 
            n23725, n23724, n23723, n23722, n23721, n23720, n23719, 
            n23718, n23717, n23716, n23715, n23714, n23713, n23712, 
            n23711, n23710, n23709, n452, PIN_8_c_2, PIN_9_c_3, 
            PIN_10_c_4, PIN_11_c_5, n453, n454, n455, n456, n23574, 
            hall3, n48211, n25, n30, n26, n27_adj_13, n15, n11, 
            n29_adj_14, n43, n41_adj_15, n387, n27_adj_16, n15_adj_17, 
            n11_adj_18, n29_adj_19, n43_adj_20, n41_adj_21, n43_adj_22, 
            n50261, n16, n50258, n15_adj_23, n11_adj_24, n43357, 
            IntegralLimit) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input [23:0]deadband;
    output \PID_CONTROLLER.result[13] ;
    output n459;
    output n460;
    output \PID_CONTROLLER.err[9] ;
    output n461;
    output \PID_CONTROLLER.err[8] ;
    output \PID_CONTROLLER.err[7] ;
    output n462;
    output \PID_CONTROLLER.err[6] ;
    output n463;
    output \PID_CONTROLLER.err[5] ;
    output \PID_CONTROLLER.result[7] ;
    output n465;
    output \PID_CONTROLLER.err[4] ;
    output \PID_CONTROLLER.err[3] ;
    output \PID_CONTROLLER.err[2] ;
    output \PID_CONTROLLER.err[1] ;
    output \PID_CONTROLLER.err[0] ;
    output [8:0]pwm_count;
    output \pwm_23__N_2960[13] ;
    input VCC_net;
    output \PID_CONTROLLER.result[5] ;
    output \pwm_23__N_2960[14] ;
    output \PID_CONTROLLER.result[14] ;
    output n467;
    output n468;
    output n469;
    output n470;
    input n50246;
    output \PID_CONTROLLER.result[21] ;
    output \pwm_23__N_2960[20] ;
    output \PID_CONTROLLER.result[20] ;
    input n27;
    input n29;
    output n471;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input n41;
    output pwm_23__N_2957;
    input \motor_state[16] ;
    output n399;
    input n24225;
    output [23:0]pwm;
    input clk32MHz;
    input n24224;
    input n24221;
    input n24220;
    input n24219;
    input n24218;
    input n24217;
    input n24214;
    input n24213;
    input n24212;
    input n24211;
    input n24210;
    input n24208;
    input n24206;
    input n24205;
    input n24204;
    input n24203;
    input n24172;
    output n400;
    input \motor_state[15] ;
    output PIN_7_c_1;
    input \motor_state[14] ;
    output PIN_6_c_0;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    output n406;
    input \motor_state[1] ;
    output n407;
    input \motor_state[0] ;
    output \PID_CONTROLLER.err_prev[31] ;
    output \PID_CONTROLLER.err_prev[23] ;
    output \PID_CONTROLLER.err_prev[22] ;
    output \PID_CONTROLLER.err_prev[21] ;
    output \PID_CONTROLLER.err_prev[20] ;
    output \PID_CONTROLLER.err_prev[19] ;
    output \PID_CONTROLLER.err_prev[18] ;
    output \PID_CONTROLLER.err_prev[17] ;
    output \PID_CONTROLLER.err_prev[16] ;
    output n413;
    output \PID_CONTROLLER.err_prev[15] ;
    output \PID_CONTROLLER.err_prev[14] ;
    output \PID_CONTROLLER.err_prev[13] ;
    output \PID_CONTROLLER.err_prev[12] ;
    output \PID_CONTROLLER.err_prev[11] ;
    input \Kd[4] ;
    input \Kp[7] ;
    output \PID_CONTROLLER.err[17] ;
    output n415;
    output \PID_CONTROLLER.err_prev[10] ;
    output \PID_CONTROLLER.err_prev[9] ;
    output \PID_CONTROLLER.err_prev[8] ;
    output \PID_CONTROLLER.err_prev[7] ;
    output \PID_CONTROLLER.err[31] ;
    output \PID_CONTROLLER.err_prev[6] ;
    input \Kp[1] ;
    output \PID_CONTROLLER.err[20] ;
    input \Kp[0] ;
    output \PID_CONTROLLER.err[21] ;
    output \PID_CONTROLLER.err_prev[5] ;
    input \Kd[0] ;
    input \Kd[1] ;
    input \Kd[2] ;
    output \PID_CONTROLLER.err_prev[4] ;
    output \PID_CONTROLLER.err_prev[3] ;
    input \Kp[2] ;
    input \Kd[5] ;
    input \Kp[3] ;
    input hall1;
    input hall2;
    input \Kp[4] ;
    output \PID_CONTROLLER.err[10] ;
    input \Kp[5] ;
    output \PID_CONTROLLER.err_prev[2] ;
    output \PID_CONTROLLER.err_prev[1] ;
    output \PID_CONTROLLER.err_prev[0] ;
    input \Kp[6] ;
    output \PID_CONTROLLER.err[11] ;
    output n853;
    output n21;
    output n855;
    output n856;
    output n857;
    output n859;
    output n860;
    output n861;
    output n862;
    output n863;
    output n864;
    output n865;
    output n866;
    output \PID_CONTROLLER.err[12] ;
    input [23:0]PWMLimit;
    input [23:0]setpoint;
    input \Kd[6] ;
    output \PID_CONTROLLER.err[16] ;
    output n867;
    output \PID_CONTROLLER.err[13] ;
    output n868;
    output n869;
    input \Ki[3] ;
    input \Kd[7] ;
    input \Ki[7] ;
    input \Kd[3] ;
    output n870;
    output n871;
    output n872;
    output n873;
    output n874;
    output n875;
    output \PID_CONTROLLER.err[15] ;
    output n46619;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    output \PID_CONTROLLER.err[14] ;
    input \Ki[1] ;
    input \Ki[0] ;
    output \PID_CONTROLLER.err[18] ;
    output \PID_CONTROLLER.err[19] ;
    input \Ki[2] ;
    output \PID_CONTROLLER.err[22] ;
    output n448;
    output n449;
    output \PID_CONTROLLER.err[23] ;
    input n23732;
    input n23731;
    input n23730;
    input n23729;
    input n23728;
    input n23727;
    input n23726;
    input n23725;
    input n23724;
    input n23723;
    input n23722;
    input n23721;
    input n23720;
    input n23719;
    input n23718;
    input n23717;
    input n23716;
    input n23715;
    input n23714;
    input n23713;
    input n23712;
    input n23711;
    input n23710;
    input n23709;
    output n452;
    output PIN_8_c_2;
    output PIN_9_c_3;
    output PIN_10_c_4;
    output PIN_11_c_5;
    output n453;
    output n454;
    output n455;
    output n456;
    input n23574;
    input hall3;
    input n48211;
    input n25;
    input n30;
    input n26;
    input n27_adj_13;
    input n15;
    input n11;
    input n29_adj_14;
    input n43;
    input n41_adj_15;
    output n387;
    input n27_adj_16;
    input n15_adj_17;
    input n11_adj_18;
    input n29_adj_19;
    input n43_adj_20;
    input n41_adj_21;
    input n43_adj_22;
    input n50261;
    input n16;
    input n50258;
    input n15_adj_23;
    input n11_adj_24;
    output n43357;
    input [23:0]IntegralLimit;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n37226;
    wire [24:0]n8104;
    
    wire n37227;
    wire [15:0]n8311;
    
    wire n50, n143;
    wire [21:0]n8446;
    wire [20:0]n8470;
    
    wire n37524, n37772;
    wire [22:0]n1802;
    
    wire n37773, n37412;
    wire [25:0]n8076;
    
    wire n37225, n37224;
    wire [16:0]n8292;
    
    wire n37411, n16_c;
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(32[23:29])
    
    wire n45, n24;
    wire [22:0]n1801;
    
    wire n37771, n37674;
    wire [22:0]n1798;
    
    wire n37675, n37223;
    wire [22:0]n1797;
    
    wire n37673;
    wire [15:0]n15397;
    wire [14:0]n15638;
    
    wire n434, n37601, n37602, n37525, n37410, n37770, n37523, 
        n37409;
    wire [31:0]n57;
    wire [8:0]n7063;
    wire [55:0]n58;
    
    wire n35914, n37222, n37672, n8, n47135, n48879, n6, n48461, 
        n35915, n36434;
    wire [9:0]n14910;
    
    wire n36435;
    wire [10:0]n14558;
    
    wire n36433, n37769, n337, n37600, n25_c, n47822, n37221, 
        n54, n37408, n37768, n37671, n36048, n49815;
    wire [31:0]n60;
    
    wire n36049, n545, n36432, n2, n36047, n37220, n36046, n36045, 
        n37219, n37522, n37407, n37218, n37217, n240, n37599, 
        n472, n37521, n37767, n37406, n37216, n37215, n399_c, 
        n37520, n37405, n37670, n50_adj_3379, n143_adj_3380, n37214, 
        n326, n37519, n37404, n37213, n36431;
    wire [9:0]n61;
    wire [9:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(33[22:30])
    
    wire n36959, n695, n37212, n598, n37211, n47842, n47091, n253, 
        n37518, n37403, n36044, n35913, n36430, n36958, n501, 
        n37210, n50234, n28894, n37402, n36957, n36043, n36956, 
        n18, n48487, n37766, n37765, n404, n37209, n36429, n36042, 
        n36955, n36428, n180, n36427, n1, n36041, n36040, n47662, 
        n37764;
    wire [5:0]n16627;
    
    wire n43968, n658, n37598, n722, n37401, n307, n37208, n37517, 
        n210, n37207;
    wire [4:0]n16635;
    
    wire n558, n37597, n625, n37400, n20_adj_3384, n113, n35, 
        n107;
    wire [26:0]n8047;
    
    wire n37206, n37205, n37669, n528, n37399, n37204;
    wire [6:0]n8437;
    wire [5:0]n9317;
    
    wire n752, n37516;
    wire [31:0]n63;
    
    wire n37203, n464, n37596, n655, n37515, n431, n37398, n37668, 
        n37202, n558_adj_3386, n37514, n35912, n48880, n37763, n370, 
        n37595, n334, n37397, n47848, n48592, n461_adj_3387, n37513, 
        n237, n37396, n364, n37512, n37762, n37667, n276, n37594, 
        n47_adj_3388, n140, n267, n37511;
    wire [17:0]n8272;
    
    wire n37395, n86, n170, n37394, n86_adj_3389, n182, n37761, 
        n37201, n37393, n48917;
    wire [13:0]n15848;
    
    wire n37593;
    wire [7:0]n8427;
    
    wire n37510, n37592, n37200, n36954, n749, n37509, n47660;
    wire [31:0]pwm_23__N_2960;
    
    wire n43891, n37199, n37392, n36953, n37198, n36952, n652, 
        n37508, n37197, n37391, n36951, n37196, n37390, n37195;
    wire [8:0]n64;
    
    wire n36950, n36949, n37194, n36948, n37666, n37591, n555, 
        n37507, n37389, n37193, n36947, n37192, n36946, n37388, 
        n37191, n36945, n37190, n36944, n458, n37506, n46591, 
        n4, n37387, n37189, n48457, n36943, n37188, n37386, n37187;
    wire [29:0]n7954;
    wire [28:0]n7986;
    
    wire n36942, n692, n37186, n36941, n37590, n361, n37505, n37385, 
        n595, n37185;
    wire [24:0]n11356;
    wire [23:0]n11990;
    
    wire n36426, n36425, n719, n37384, n26834, n36039, n498, n37184, 
        n36424, n48458, n36423, n36422, n50255, n47784, n46999, 
        n264, n37504, n622, n37383, n50243, n37760, n401, n37183, 
        n36421, n36420, n30_c, n10, n46995, n48881, n36419, n525, 
        n37382, n304, n37182, n36418, n36417, n36038, n36416, 
        n36037, n515, n37665, n37589, n74, n167, n428, n37381, 
        n207, n37181, n36415, n36414, n36413, n331, n37380, n47666, 
        n17, n110, n36412, n36411, n36036, n36410;
    wire [8:0]n8416;
    
    wire n37503, n234, n37379;
    wire [27:0]n8017;
    
    wire n37180, n36409, n37179, n698, n36408, n601, n36407, n37502, 
        n44_adj_3398, n137, n504, n36406, n37178, n407_c, n36405, 
        n36035, n49053, n37759, n37588;
    wire [18:0]n8251;
    
    wire n37378, n49054, n37177, n37377, n48987, n37176, n746, 
        n37501, n49004, n46958, n37175, n37376, n37174, n442, 
        n37664, n37587, n37173, n37375, n37172, n649, n37500, 
        n37171, n37374, n37170, n37758, n37586, n37373, n552, 
        n37499, n37372, n369, n37663, n728, n37585, n47664, n48954, 
        n50239, n46953, n49103, n37371, n455_c, n37498, n37370, 
        n47672, n631, n37584, n37369, n37169, n358, n37497, n37168, 
        n36940, n36939, n37368, n37167, n36938, n49109, n36937, 
        n37166, n37367, n37165, n261, n37496, n37164, n36936, 
        n36935, n716, n37366, n37163, n36934, n36933, n296, n37662, 
        n534, n37583, n8_adj_3401, n37162, n619, n37365, n37161, 
        n71, n164, n44147, n37160, n36932, n36931, n36930, n522, 
        n37364, n49110, n689, n37159, n36929, n4_adj_3402, n36928, 
        n48471;
    wire [9:0]n8404;
    
    wire n37495, n425, n37363, n592_adj_3404, n37158, n48472, n495, 
        n37157, n37494, n328, n37362, n398, n37156, n36927, n33, 
        n31_adj_3406, n47187, n47171, n36926, n301, n37155, n36925, 
        n527, n37757, n437, n37582, n231, n37361, n204, n37154, 
        n37493, n41_c, n134, n36924, n310, n36404, n14, n107_adj_3409, 
        n213, n36403, n23_adj_3410, n116;
    wire [8:0]n15224;
    
    wire n36402, n37153, n36401, n36400;
    wire [24:0]\PID_CONTROLLER.err_31__N_2825 ;
    wire [24:0]n66;
    
    wire n36153;
    wire [19:0]n8229;
    
    wire n37360, n37359, n743, n37492, n37152, n36399, n36398, 
        n36152, n36397, n37358, n37151, n36396, n36395, n36151;
    wire [31:0]n67;
    
    wire n36034, n36394, n36150, n36033, n223, n37661, n340, n37581, 
        n37357, n30_adj_3414, n10_adj_3415, n35_adj_3416, n47167, 
        n48877, n646, n37491, n37356, n37150, n37149, n36149, 
        n47650, n37355, n37148, n49051, n37, n49052, n36148, n36032, 
        n36147, n243, n37580, n549, n37490, n37354, n37147, n36146;
    wire [22:0]n12573;
    
    wire n36387, n36386, n37353, n37146, n36385, n36384, n39, 
        n48991, n49081, n49123, n48919, n47656, pwm_23__N_2959, 
        n48921, n36145, n36031, n452_c, n37489, n24223, n24222, 
        n24216, n24215, n24209, n24207, n37145, n454_c, n37756, 
        n150, n37660, n36030, n37352, n381, n37755, n36923, n37144, 
        n308, n37754, n37143, n36383, n35911, n37142, n36922, 
        n36921, n53_adj_3424, n146, n37351, n37141, n37140, n36920, 
        n683, n36919, n355, n37488, n37350, n37139, n37138, n586, 
        n36918, n489, n36917, n235, n37753, n37349, n37137, n37348, 
        n392, n36916, n36144, n258, n37487;
    wire [31:0]\PID_CONTROLLER.result_31__N_3003 ;
    wire [5:0]GATES_5__N_2788;
    
    wire n37136, n36029, n36143, n36382, n36381, n713, n37347, 
        n36380, n37135, n36379, n616, n37346, n36142, n36141;
    wire [6:0]n16618;
    
    wire n752_adj_3431, n37579, n36378, n295, n36915, n37134, n198, 
        n36914, n36140, n36028, n8_adj_3433, n101, n36377, n37578, 
        n68, n161, n519_adj_3434, n37345, n36139, n36376, n37133, 
        n162, n37752, n36375, n36138, n36374, n422, n37344, n36373, 
        n37132, n36027, n36137, n36372, n20_adj_3439, n89, n36026, 
        n36136, n36371, n8_adj_3443, n77;
    wire [10:0]n8391;
    
    wire n37486, n325, n37343, n37577, n701, n36370, n686, n37131, 
        n604_adj_3444, n36369, n36135, n507, n36368, n37485, n228, 
        n37342, n410, n36367, n589_adj_3446, n37130, n36134, n313, 
        n36366, n36133, n36025, n216, n36365, n37484, n38, n131_adj_3450, 
        n492, n37129, n26_adj_3451, n119, n36364, n36132, n583, 
        n36363, n510, n36362;
    wire [20:0]n8206;
    
    wire n37341, n37340, n35910, n395, n37128, n437_adj_3453, n36361, 
        n36131, n36024, n364_adj_3455, n36360;
    wire [14:0]n12730;
    wire [13:0]n13254;
    
    wire n36913, n35909, n36912, n291, n36359;
    wire [22:0]n1800;
    
    wire n37750, n1699, n37749;
    wire [22:0]n1796;
    
    wire n37658, n37576, n37483, n298, n37127, n37339, n201, n37126, 
        n11_adj_3457, n104, n37338;
    wire [0:0]n7059;
    
    wire n37125;
    wire [31:0]n69;
    wire [55:0]n191;
    
    wire n37124, n1683, n37575, n740, n37482, n37123, n37337, 
        n37122, n37121, n37336;
    wire [33:0]n282;
    
    wire n37657, n37574, n643, n37481, n37335, n37334, n546, n37480, 
        n37333, n37332, n37748, n37656;
    wire [12:0]n16029;
    
    wire n37573, n449_c, n37479, n37120, n37331, n37119, n36911, 
        n37118, n36910, n37330, n36909, n37117, n36908, n37572, 
        n352, n37478, n37329, n37116, n37115, n36130, n37328, 
        n37114, n36907, n36906, n218_adj_3463, n36358, n37113, n36905, 
        n36904, n37112, n255, n37477, n710, n37327, n37111, n37747, 
        n36023, n36903, n145, n36357, n36902, n36901, n37110, 
        n36022, n37109, n72, n613, n37326, n36900;
    wire [21:0]n13107;
    
    wire n36356, n37108;
    wire [6:0]n70;
    wire [6:0]Kd_delay_counter;   // verilog/motorControl.v(27[13:29])
    
    wire n36899, n36898, n37107, n36897, n37106, n516_adj_3471, 
        n37325, n36129, n36896, n36021, n37571, n36895, n65, n158, 
        n37105, n36128, n36355, n419, n37324, n37104, n36020, 
        n36127, n37103, n36894, n322, n37323, n37102, n37746, 
        n37655, n37570;
    wire [11:0]n8377;
    
    wire n37476, n680, n37101, n225_adj_3485, n37322, n37475, n36354, 
        n583_adj_3486, n37100, n36353, n36352, n35_adj_3487, n128, 
        n36351, n486, n37099, n36126, n36350, n36125, n36349;
    wire [21:0]n8182;
    
    wire n37321, n37474, n37320, n36348, n389, n37098, n36124, 
        n36347, n36346, n36345, n292, n37097, n36123, n36019, 
        n36344, n36122, n36018, n36343, n37569, n37319, n37473, 
        n37318, n36342, n195, n37096, n36121, n36341, n704, n36340, 
        n607, n36339, n5_adj_3496, n98, n36120, n36017, n510_adj_3498, 
        n36338, n36119, n413_adj_3500, n36337, n37317, n37472, n37316, 
        n316, n36336;
    wire [19:0]n9325;
    wire [18:0]n10116;
    
    wire n37095, n36118, n219_adj_3502, n36335, n37654, n35908, 
        n37653, n37568, n29_adj_3505, n122, n737, n37471, n36117;
    wire [10:0]n16312;
    wire [9:0]n16418;
    
    wire n36334, n36333, n640, n37470, n37652, n37651, n37094, 
        n37745, n36332, n36116, n37744, n37093, n36016, n37650, 
        n37315, n36331, n37743, n37649, n35907, n36115, n740_adj_3511, 
        n36330, n446_adj_3512, n37742, n731, n37741, n643_adj_3513, 
        n36329, n37092, n546_adj_3514, n36328, n37091, n36015, n37648, 
        n37740, n35906, n36114, n449_adj_3518, n36327, n37739, n36113, 
        n352_adj_3520, n36326, n543, n37469, n36014, n36112, n37314, 
        n37090, n36013, n255_adj_3523, n36325, n35905, n37567, n65_adj_3524, 
        n158_adj_3525, n37089, n36111, n36012;
    wire [0:0]n5784;
    wire [29:0]n6540;
    
    wire n36644, n36643, n37313, n36642;
    wire [20:0]n13592;
    
    wire n36324, n36323, n37088, n36641, n36322, n36640, n36321, 
        n36320, n37566, n36639, n37468, n37312, n36638, n36319, 
        n36637, n36011, n37738, n37087, n36636, n36318, n36635, 
        n36317, n36110, n36634, n46593, n37086, n37311, n36633, 
        n37647, n36632, n37737, n37736, n36316, n36109, n36315, 
        n36631, n37085;
    wire [4:0]n10109;
    
    wire n35704;
    wire [22:0]n1804;
    
    wire n1711, n37870;
    wire [23:0]n73;
    wire [23:0]n75;
    
    wire n36010, n36314, n36313;
    wire [22:0]n1803;
    
    wire n1707, n37869, n36630, n37735, n524, n37734, n1703, n37868, 
        n36108, n451, n37733, n378, n37732, n37867, n37646, n305_adj_3538, 
        n37731, n1695, n37866, n36629, n45_adj_3539, n36009;
    wire [22:0]n1799;
    
    wire n1691, n37865, n36107, n36312, n36628, n1687, n37864, 
        n35904, n37863, n37084, n232_adj_3543, n37730, n370_adj_3544, 
        n4_adj_3545, n7_adj_3546, n36311, n35903, n36627, n36310, 
        n36626, n37862, n37861, n159, n37729, n37860, n634, n37565, 
        n37645, n349, n37467, n37310, n37083, n37859, n37309, 
        n37082, n537, n37564;
    wire [5:0]GATES_5__N_3048;
    
    wire n5_adj_3549, n252, n37466, n37308, n37081, n37858, n62, 
        n155, n37080;
    wire [12:0]n8362;
    
    wire n37465, n37079, n37307, n37078, n37464, n36625, n707, 
        n37306, n37077, n440, n37563, n37463, n610, n37305, n36624, 
        n707_adj_3552, n36309, n43988, n658_adj_3553, n37076, n564, 
        n37075, n17_adj_3554, n86_adj_3555, n37644, n343, n37562, 
        n37462, n513, n37304, n37461, n416_adj_3557, n37303, n246_adj_3558, 
        n37561, n37460, n319, n37302, n37727, n36623, n610_adj_3559, 
        n36308, n734, n37459, n222_adj_3560, n37301, n37857, n37643, 
        n56, n149, n637, n37458, n32_adj_3562, n125;
    wire [3:0]n10844;
    
    wire n464_adj_3563, n37074, n37073;
    wire [22:0]n8157;
    
    wire n37300, n276_adj_3564, n37072, n37726, n37856, n37299, 
        n36622, n182_adj_3565, n540, n37457;
    wire [17:0]n10850;
    
    wire n37071, n37070, n37298, n37069, n37068, n37297, n43_adj_3566, 
        n36008, n36106, n36621, n35902, n513_adj_3570, n36307, n37067, 
        n36105;
    wire [11:0]n16183;
    
    wire n37560, n443_adj_3572, n37456, n37066, n37296, n37065, 
        n680_adj_3574, n36620, n37064, n416_adj_3575, n36306, n37295, 
        n41_adj_3576, n36007, n583_adj_3579, n36619, n319_adj_3580, 
        n36305, n37063, n37559, n346, n37455, n37062, n37294, 
        n37061, n486_adj_3581, n36618, n37060, n37293, n37059, n389_adj_3583, 
        n36617, n512, n37642, n249, n37454, n37292, n37058, n222_adj_3585, 
        n36304, n292_adj_3587, n36616, n37057, n32_adj_3588, n125_adj_3589;
    wire [19:0]n14033;
    
    wire n36303, n36302, n37558, n39_adj_3590, n36006, n195_adj_3593, 
        n36615, GATES_5__N_3055, n36104, n37_adj_3594, n36005, n37291, 
        n37056, n5_adj_3596, n98_adj_3597, n36301;
    wire [23:0]n76;
    
    wire n36103;
    wire [23:0]n852;
    
    wire n36300, n36299, n36102, n36298, n59, n152_adj_3601, n36101, 
        n37290, n37055, n36297, n36296, n35_adj_3603, n36004, n37054, 
        n36295, n36100, n36294, n37289, n36293;
    wire [28:0]n7758;
    
    wire n36607, n36099, n36292, n37725, n33_adj_3607, n36003, n36606, 
        n36291, n31_adj_3609, n36002, n36098, n36605, n36290, n29_adj_3612, 
        n36001, n36097, n439, n37641, n37557;
    wire [16:0]n11529;
    
    wire n37053;
    wire [13:0]n8346;
    
    wire n37453, n37288, n37052, n366, n37640, n37287, n36604, 
        n710_adj_3616, n36289, n36603, n613_adj_3617, n36288, n516_adj_3618, 
        n36287, n36096, n37452, n37051, n37286, n36602, n419_adj_3620, 
        n36286, n36601, n322_adj_3621, n36285, n37050, n36095, n225_adj_3623, 
        n36284, n36600, n35_adj_3624, n128_adj_3625, n27_adj_3626, 
        n36000, n36094, n37285, n37049, n36599;
    wire [8:0]n16503;
    
    wire n36283, n36282, n36598, n36093, n36281, n36597, n36092, 
        n743_adj_3631, n36280, n37724, n37451, n704_adj_3632, n37284, 
        n37048, n37855, n36596, n646_adj_3633, n36279, n36595, n25_adj_3634, 
        n35999, n36091, n549_adj_3637, n36278, n37854, n37853, n37723, 
        n37852, n37450, n37556, n37851, n37722, n607_adj_3638, n37283, 
        n293, n37639, n36594, n23_adj_3640, n35998, n37047, n510_adj_3642, 
        n37282, n37046, n37045, n37555, n37449, n413_adj_3643, n37281, 
        n452_adj_3644, n36277, n37044, n36593, n316_adj_3645, n37280, 
        n37043, n355_adj_3646, n36276, n36592, n258_adj_3647, n36275, 
        n36591, n68_adj_3648, n161_adj_3649, n36590;
    wire [18:0]n14432;
    
    wire n36274, n36589, n37042, n36273, n37041, n220_adj_3651, 
        n37638, n734_adj_3652, n37554, n37721, n37720, n37850, n147_adj_3653, 
        n37637, n37719, n36588, n36272, n36587, n37849, n37718, 
        n36271, n36586, n36270, n36585, n37448, n36269, n219_adj_3654, 
        n37279, n37040, n37039, n36268, n683_adj_3655, n36584, n37717, 
        n36267, n586_adj_3656, n36583, n36266, n489_adj_3657, n36582, 
        n36265, n392_adj_3658, n36581, n29_adj_3659, n122_adj_3660, 
        n37038, n36264, n295_adj_3661, n36580, n36263, n198_adj_3662, 
        n36579, n37037, n36262, n8_adj_3663, n101_adj_3664;
    wire [27:0]n9123;
    
    wire n36578, n713_adj_3665, n36261, n36577, n37447;
    wire [23:0]n8131;
    
    wire n37278, n36090, n616_adj_3667, n36260, n519_adj_3668, n36259, 
        n36576, n21_adj_3669, n35997, n36575, n637_adj_3671, n37553;
    wire [15:0]n12155;
    
    wire n37036, n35901, n37277, n37848, n35916, n35917, n37716, 
        n37847, n422_adj_3672, n36258, n36574, n5_adj_3673, n74_adj_3674, 
        n36089, n37715, n731_adj_3676, n37446, n37035, n37846, n35900, 
        n540_adj_3677, n37552, n36573, n325_adj_3678, n36257, n36572, 
        n228_adj_3679, n36256, n37276, n36571, n38_adj_3680, n131_adj_3681, 
        n36570;
    wire [17:0]n14791;
    
    wire n36255, n37034, n37275, n35899, n37845, n37033, n36569, 
        n36254, n36568, n36253, n36567, n634_adj_3682, n37445, n37032, 
        n36252, n36566, n36565, n36251, n36564, n37031, n19_adj_3683, 
        n35996, n36088, n37274, n37714;
    wire [16:0]n15112;
    
    wire n37636, n37273, n443_adj_3686, n37551, n537_adj_3687, n37444, 
        n37272, n37635, n36250, n36563, n36249, n37030, n36562, 
        n37844, n37271, n346_adj_3688, n37550, n440_adj_3689, n37443, 
        n36248, n36561, n36247, n36560, n36246, n37270, n343_adj_3690, 
        n37442, n37269, n37029, n36559, n37268, n37028, n37713, 
        n37267, n246_adj_3691, n37441, n37027, n36245, n249_adj_3692, 
        n37549, n37026, n37634, n59_adj_3693, n152_adj_3694, n37548, 
        n35898, n37266, n37025, n37547, n37024, n36087, n37023, 
        n56_adj_3696, n149_adj_3697, n37265, n17_adj_3698, n35995, 
        n36558, n37843, n37633, n37022, n37021, n36557, n35897, 
        n37546, n37264, n37842, n37712, n36244, n36086, n15_adj_3702, 
        n35994;
    wire [14:0]n8329;
    
    wire n37440, n686_adj_3704, n36556, n37841, n37632, n36085, 
        n35896, n35895, n35894, n589_adj_3706, n36555, n492_adj_3707, 
        n36554, n36084, n37263, n37439, n35893, n37020, n37262, 
        n37631, n701_adj_3709, n37261, n37438, n37545, n37019, n521, 
        n37711, n37630, n37840, n35892, n37544, n37629, n37839, 
        n448_c, n37710, n37838, n37018, n37017, n37016, n37437, 
        n604_adj_3712, n37260, n37015, n37014, n737_adj_3713, n37543, 
        n507_adj_3714, n37259, n37013, n37012, n37436, n410_adj_3715, 
        n37258, n37011, n37010, n375, n37709, n313_adj_3716, n37257, 
        n37435, n216_adj_3717, n37256, n37009, n395_adj_3718, n36553, 
        n716_adj_3719, n36243, n619_adj_3720, n36242, n298_adj_3721, 
        n36552, n201_adj_3722, n36551, n35891, n37837, n640_adj_3723, 
        n37542, n36083, n37628, n543_adj_3725, n37541, n55_adj_3726, 
        n36082, n522_adj_3728, n36241, n37008, n11_adj_3729, n104_adj_3730, 
        n28817, n35890, n37007, n425_adj_3732, n36240, n13_adj_3733, 
        n35993, n37836, n37835, n328_adj_3735, n36239, n302_adj_3737, 
        n37708;
    wire [12:0]n13732;
    
    wire n36550, n11_adj_3738, n35992, n26_adj_3740, n119_adj_3741, 
        n37834, n36549, n37833, n36548, n231_adj_3742, n36238, n9_adj_3743, 
        n35991, n35889, n7_adj_3745, n35990, n36547, n37006, n41_adj_3747, 
        n134_adj_3748, n37434, n36546, n37255, n37254, n229_adj_3750, 
        n37707;
    wire [7:0]n16569;
    
    wire n36237, n36545, n37832, n37627, n37831, n36544, n446_adj_3751, 
        n37540, n36236, n37253, n37252, n37433, n349_adj_3752, n37539, 
        n5_adj_3753, n35989, n746_adj_3755, n36235, n36543, n722_adj_3756, 
        n37626, n36542, n649_adj_3757, n36234, n3_adj_3758, n35988, 
        n728_adj_3760, n37432, n37251, n252_adj_3763, n37538, n631_adj_3764, 
        n37431, n37250, n625_adj_3765, n37625, n62_adj_3766, n155_adj_3767, 
        n36541, n552_adj_3768, n36233, n156_adj_3769, n37706, n36540, 
        n455_adj_3770, n36232, n36539, n534_adj_3771, n37430, n35888, 
        n437_adj_3772, n37429, n358_adj_3773, n36231, n36538, n37537, 
        n261_adj_3774, n36230, n37249, n37830;
    wire [26:0]n9927;
    
    wire n36537, n35887, n71_adj_3775, n164_adj_3776, n36536, n36535, 
        n37829;
    wire [31:0]n79;
    
    wire n35987, n35986, n36534, n14_adj_3778, n83, n37704, n37536, 
        n36533, n340_adj_3779, n37428, n35985, n528_adj_3783, n37624, 
        n243_adj_3784, n37427, n37248, n53_adj_3785, n146_adj_3786, 
        n37828, n37827, n431_adj_3789, n37623, n536, n37826, n37535, 
        n463_adj_3792, n37825, n36532, n37703, n37426, n334_adj_3793, 
        n37622, n36531, n37534, n37247, n36530, n36529, n36528, 
        n36527, n37425, n37246, n36526, n36224, n36223, n36525, 
        n35984, n36524, n36222, n36523, n36221, n35983, n36220, 
        n36522, n35982, n36521, n36520, n36519, n390, n37824, 
        n36219, n36518, n36517, n36218, n37245, n689_adj_3797, n36516, 
        n592_adj_3798, n36515, n36217, n37702, n237_adj_3799, n37621, 
        n35981, n495_adj_3801, n36514, n398_adj_3802, n36513, n36216, 
        n301_adj_3803, n36512, n35980, n204_adj_3805, n36511, n36215, 
        n14_adj_3806, n107_adj_3807, n35979, n36214;
    wire [11:0]n14166;
    
    wire n36510, n35978, n36509, n36213, n36508, n37244, n36507, 
        n317, n37823, n37701, n36506, n37424, n36212, n36505, 
        n37243, n244_adj_3811, n37822, n36211, n37242, n37700, n37533, 
        n36504, n36210, n36503, n36502, n36209, n36501, n37241, 
        n36208, n36500, n37423, n36207, n36499, n35977, n37699;
    wire [25:0]n10669;
    
    wire n36498, n47_adj_3813, n140_adj_3814, n35976, n36497, n36496, 
        n37532, n36206, n35975, n36495, n36205, n35974, n35561, 
        n37873, n37620, n37422, n37240, n171_adj_3819, n37821, n36204, 
        n37531, n37239, n37421, n98_adj_3820, n36494, n36203, n36202, 
        n36493, n35973, n7_adj_3822, n8_adj_3823, n8_adj_3824, n37819, 
        n749_adj_3825, n37619, n37818, n37530, n36201, n36492, n37238, 
        n37698, n37817, n37816, n37815, n37814, n652_adj_3826, n37618, 
        n37697, n37813, n37812, n37696, n37420, n698_adj_3827, n37237, 
        n555_adj_3828, n37617, n37419, n36200, n601_adj_3829, n37236, 
        n35972, n36491, n36490, n458_adj_3831, n37616, n35971, n361_adj_3833, 
        n37615, n37695, n36489, n36199, n36488, n37694, n37529, 
        n36487, n36198, n37811, n35970, n36486, n36485, n504_adj_3835, 
        n37235, n407_adj_3836, n37234, n36484, n36197, n264_adj_3837, 
        n37614, n37418, n36483, n37693, n37692, n35969, n37691, 
        n37810, n36196, n37809, n167_adj_3839, n36482, n37808, n37807, 
        n35968, n37806, n37805, n37613, n37612, n37611, n36481, 
        n37804, n533, n37803, n460_adj_3845, n37802, n36195, n37690, 
        n310_adj_3846, n37233, n36057, n36480, n37610, n36056, n35967, 
        n36479, n28362, n36055, n37528, n37689, n692_adj_3850, n36478, 
        n387_c, n37801, n518, n37688, n314_adj_3852, n37800, n241_adj_3854, 
        n37799, n168_adj_3856, n37798, n445, n37687, n26_adj_3857, 
        n95, n37609, n35966, n37527, n37796, n595_adj_3859, n36477, 
        n36194, n498_adj_3860, n36476, n725, n37417, n401_adj_3861, 
        n36475, n372, n37686, n37795, n37794, n213_adj_3862, n37232, 
        n304_adj_3863, n36474, n37526, n207_adj_3864, n36473, n17_adj_3865, 
        n110_adj_3866, n36193, n36472, n36471, n36192, n36470, n36469, 
        n36191, n37793, n36468, n36467, n36190, n628, n37416, 
        n23_adj_3867, n116_adj_3868, n37792, n36466, n36189, n1_adj_3869, 
        n36054, n35965, n37608, n36465, n299_adj_3871, n37685, n36188, 
        n36464, n531_adj_3872, n37415, n35964, n36463, n36462, n36187, 
        n37231, n36186, n36461, n36460, n36053, n36459, n36185, 
        n36458, n36457, n36184, n434_adj_3876, n37414, n37230, n36456, 
        n36455, n36183, n226_adj_3877, n37684, n36454, n36453, n719_adj_3878, 
        n36182, n36452, n36451, n37229, n36450, n337_adj_3879, n37413, 
        n622_adj_3880, n36181, n36449, n36448, n525_adj_3881, n36180, 
        n153_adj_3882, n37683, n36052, n11_adj_3883, n80, n37681, 
        n37680, n36447, n36446, n428_adj_3884, n36179, n36445, n331_adj_3885, 
        n36178, n37228, n36051, n36444, n37791, n36443, n695_adj_3887, 
        n36442, n37679, n37607, n36050, n598_adj_3889, n36441, n234_adj_3890, 
        n36177, n501_adj_3891, n36440, n404_adj_3892, n36439, n44_adj_3893, 
        n137_adj_3894, n37790, n307_adj_3895, n36438, n210_adj_3896, 
        n36437, n20_adj_3897, n113_adj_3898, n37789, n240_adj_3899, 
        n37788, n36436, n37787, n27734, n37786, n37606, n37678, 
        n37785, n37784, n37783, n37605, n37782, n37781, n37677, 
        n725_adj_3900, n37604, n37676, n530, n37780, n457, n37779, 
        n384, n37778, n311_adj_3901, n37777, n628_adj_3902, n37603, 
        n238_adj_3903, n37776, n165_adj_3904, n37775, n23_adj_3905, 
        n92, n531_adj_3906, n878, n17_adj_3907, n42366, n20_adj_3908, 
        n26_adj_3909, n24_adj_3910, n28_adj_3911, n23_adj_3912, n42312, 
        n39_adj_3916, n45_adj_3917, n43127, n46681, n37_adj_3918, 
        n18_adj_3919, n31_adj_3920, n21_adj_3921, n23_adj_3922, n25_adj_3923, 
        n17_adj_3924, n19_adj_3925, n9_adj_3926, n35_adj_3927, n33_adj_3928, 
        n13_adj_3929, n46817, n12_adj_3933, n10_adj_3934, n30_adj_3935, 
        n46851, n47591, n47585, n48723, n48175, n48907, n6_adj_3937, 
        n48757, n48758, n16_adj_3939, n8_adj_3940, n24_adj_3941, n46826, 
        n46793, n46791, n48960, n48500, n10_adj_3942, n8_adj_3943, 
        n12_adj_3944, n4_adj_3945, n48675, n48676, n46811, n46807, 
        n48958, n48502, n49093, n49094, n49046, n46795, n49101, 
        n48997, n49111, n43881, n49112, n7_adj_3948, n13_adj_3949, 
        n23_adj_3950, n9_adj_3951, n17_adj_3952, n19_adj_3953, n21_adj_3954, 
        n39_adj_3955, n45_adj_3956, n37_adj_3957, n31_adj_3958, n23_adj_3959, 
        n25_adj_3960, n35_adj_3961, n33_adj_3962, n9_adj_3963, n17_adj_3964, 
        n19_adj_3965, n21_adj_3966, n13_adj_3967, n46893, n46887, 
        n12_adj_3971, n30_adj_3972, n46916, n47677, n47673, n48745, 
        n48201, n48911, n6_adj_3974, n48681, n48682, n16_adj_3975, 
        n24_adj_3976, n46858, n8_adj_3978, n46854, n48497, n48492, 
        n4_adj_3979, n48679, n48680, n46878, n10_adj_3980, n46875, 
        n48956, n48494, n49091, n49092, n49048, n46860, n48753, 
        n40_adj_3982, n48755, n48_adj_3983, n44079, n44083, n56_adj_3984, 
        n44134, n44139, n47930, n47205, n47139, n48279, n48811, 
        n47041, n47806, n12_adj_3986, n47053, n50290, n47047, n50319, 
        n48249, n50293, n19_adj_3988, n44357, n44353, n44355, n47804, 
        n29_adj_3989, n50307, n6_adj_3990, n48584, n50302, n47010, 
        n46652, n48237, n50313, n48793, n50249, n16_adj_3991, n46950, 
        n8_adj_3992, n24_adj_3993, n47031, n47800, n6_adj_3994, n48459, 
        n48460, n47796, n12_adj_3997, n47960, n48323, n48317, n47191, 
        n48610, n49025, n47878, n48600, n48942, n12_adj_3998, n6_adj_3999, 
        n8_adj_4000, n8_adj_4001, n35689, n8_adj_4002, n18_adj_4003, 
        n24_adj_4004, n22_adj_4005, n26_adj_4006, n43653, n11_adj_4007, 
        n9_adj_4008, n17_adj_4009, n48056, n48054, n47257, n50541, 
        n48070, n48038, n47303, n50529, n10_adj_4010, n30_adj_4011, 
        n5_adj_4012, n48060, n47358, n47350, n48369, n48843, n48044, 
        n48628, n48950, n49085, n6_adj_4013, n47460, n24_adj_4014, 
        n48481, n47275, n50494, n48485, n47638, n4_adj_4015, n48475, 
        n48476, n8_adj_4016, n47241, n6_adj_4017, n16_adj_4018, n47247, 
        n48582, n47648, n48915, n4_adj_4019, n48479, n47307, n48875, 
        n47640, n49049, n49050, n48002, n48747, n47646, n48916, 
        n48913, n4_adj_4020, n6_adj_4021;
    
    SB_CARRY add_3058_22 (.CI(n37226), .I0(n8104[19]), .I1(GND_net), .CO(n37227));
    SB_LUT4 add_3068_2_lut (.I0(GND_net), .I1(n50), .I2(n143), .I3(GND_net), 
            .O(n8311[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_10_lut (.I0(GND_net), .I1(n8470[7]), .I2(GND_net), 
            .I3(n37524), .O(n8446[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_23 (.CI(n37772), .I0(n1802[20]), .I1(GND_net), 
            .CO(n37773));
    SB_CARRY add_3068_2 (.CI(GND_net), .I0(n50), .I1(n143), .CO(n37412));
    SB_LUT4 add_3058_21_lut (.I0(GND_net), .I1(n8104[18]), .I2(GND_net), 
            .I3(n37225), .O(n8076[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_21 (.CI(n37225), .I0(n8104[18]), .I1(GND_net), .CO(n37226));
    SB_LUT4 add_3058_20_lut (.I0(GND_net), .I1(n8104[17]), .I2(GND_net), 
            .I3(n37224), .O(n8076[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_18_lut (.I0(GND_net), .I1(n8311[15]), .I2(GND_net), 
            .I3(n37411), .O(n8292[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i24_3_lut  (.I0(n16_c), .I1(\PID_CONTROLLER.result [22]), 
            .I2(n45), .I3(GND_net), .O(n24));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_3058_20 (.CI(n37224), .I0(n8104[17]), .I1(GND_net), .CO(n37225));
    SB_LUT4 mult_14_add_1216_22_lut (.I0(GND_net), .I1(n1802[19]), .I2(GND_net), 
            .I3(n37771), .O(n1801[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_17 (.CI(n37674), .I0(n1798[14]), .I1(GND_net), 
            .CO(n37675));
    SB_LUT4 add_3058_19_lut (.I0(GND_net), .I1(n8104[16]), .I2(GND_net), 
            .I3(n37223), .O(n8076[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_16_lut (.I0(GND_net), .I1(n1798[13]), .I2(GND_net), 
            .I3(n37673), .O(n1797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3387_5_lut (.I0(GND_net), .I1(n15638[2]), .I2(n434), .I3(n37601), 
            .O(n15397[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_5 (.CI(n37601), .I0(n15638[2]), .I1(n434), .CO(n37602));
    SB_CARRY add_3058_19 (.CI(n37223), .I0(n8104[16]), .I1(GND_net), .CO(n37224));
    SB_CARRY mult_14_add_1212_16 (.CI(n37673), .I0(n1798[13]), .I1(GND_net), 
            .CO(n37674));
    SB_CARRY mult_14_add_1216_22 (.CI(n37771), .I0(n1802[19]), .I1(GND_net), 
            .CO(n37772));
    SB_CARRY add_3078_10 (.CI(n37524), .I0(n8470[7]), .I1(GND_net), .CO(n37525));
    SB_LUT4 add_3067_17_lut (.I0(GND_net), .I1(n8311[14]), .I2(GND_net), 
            .I3(n37410), .O(n8292[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_21_lut (.I0(GND_net), .I1(n1802[18]), .I2(GND_net), 
            .I3(n37770), .O(n1801[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_17 (.CI(n37410), .I0(n8311[14]), .I1(GND_net), .CO(n37411));
    SB_LUT4 add_3078_9_lut (.I0(GND_net), .I1(n8470[6]), .I2(GND_net), 
            .I3(n37523), .O(n8446[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_16_lut (.I0(GND_net), .I1(n8311[13]), .I2(GND_net), 
            .I3(n37409), .O(n8292[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_30_lut (.I0(GND_net), .I1(n7063[5]), 
            .I2(n58[28]), .I3(n35914), .O(n57[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_18_lut (.I0(GND_net), .I1(n8104[15]), .I2(GND_net), 
            .I3(n37222), .O(n8076[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_15_lut (.I0(GND_net), .I1(n1798[12]), .I2(GND_net), 
            .I3(n37672), .O(n1797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_21 (.CI(n37770), .I0(n1802[18]), .I1(GND_net), 
            .CO(n37771));
    SB_LUT4 i33318_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n47135), 
            .O(n48879));   // verilog/motorControl.v(44[10:27])
    defparam i33318_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32900_3_lut (.I0(n6), .I1(\PID_CONTROLLER.result [26]), .I2(deadband[23]), 
            .I3(GND_net), .O(n48461));   // verilog/motorControl.v(44[10:27])
    defparam i32900_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_13_add_1_21902_add_1_30 (.CI(n35914), .I0(n7063[5]), .I1(n58[28]), 
            .CO(n35915));
    SB_CARRY add_3340_10 (.CI(n36434), .I0(n14910[7]), .I1(GND_net), .CO(n36435));
    SB_CARRY add_3058_18 (.CI(n37222), .I0(n8104[15]), .I1(GND_net), .CO(n37223));
    SB_LUT4 add_3340_9_lut (.I0(GND_net), .I1(n14910[6]), .I2(GND_net), 
            .I3(n36433), .O(n14558[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_20_lut (.I0(GND_net), .I1(n1802[17]), .I2(GND_net), 
            .I3(n37769), .O(n1801[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_20 (.CI(n37769), .I0(n1802[17]), .I1(GND_net), 
            .CO(n37770));
    SB_LUT4 add_3387_4_lut (.I0(GND_net), .I1(n15638[1]), .I2(n337), .I3(n37600), 
            .O(n15397[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32261_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [29]), 
            .I2(\PID_CONTROLLER.result [30]), .I3(n25_c), .O(n47822));
    defparam i32261_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 add_3058_17_lut (.I0(GND_net), .I1(n8104[14]), .I2(GND_net), 
            .I3(n37221), .O(n8076[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_17 (.CI(n37221), .I0(n8104[14]), .I1(GND_net), .CO(n37222));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i54_4_lut  (.I0(\PID_CONTROLLER.result [12]), 
            .I1(\PID_CONTROLLER.result [30]), .I2(deadband[23]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n54));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i54_4_lut .LUT_INIT = 16'h8f0e;
    SB_CARRY add_3067_16 (.CI(n37409), .I0(n8311[13]), .I1(GND_net), .CO(n37410));
    SB_LUT4 add_3067_15_lut (.I0(GND_net), .I1(n8311[12]), .I2(GND_net), 
            .I3(n37408), .O(n8292[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_9 (.CI(n37523), .I0(n8470[6]), .I1(GND_net), .CO(n37524));
    SB_CARRY mult_14_add_1212_15 (.CI(n37672), .I0(n1798[12]), .I1(GND_net), 
            .CO(n37673));
    SB_LUT4 mult_14_add_1216_19_lut (.I0(GND_net), .I1(n1802[16]), .I2(GND_net), 
            .I3(n37768), .O(n1801[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_14_lut (.I0(GND_net), .I1(n1798[11]), .I2(GND_net), 
            .I3(n37671), .O(n1797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3340_9 (.CI(n36433), .I0(n14910[6]), .I1(GND_net), .CO(n36434));
    SB_CARRY unary_minus_23_add_3_16 (.CI(n36048), .I0(n49815), .I1(n60[14]), 
            .CO(n36049));
    SB_LUT4 add_3340_8_lut (.I0(GND_net), .I1(n14910[5]), .I2(n545), .I3(n36432), 
            .O(n14558[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_15_lut (.I0(\PID_CONTROLLER.result[13] ), 
            .I1(n49815), .I2(n60[13]), .I3(n36047), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3067_15 (.CI(n37408), .I0(n8311[12]), .I1(GND_net), .CO(n37409));
    SB_CARRY unary_minus_23_add_3_15 (.CI(n36047), .I0(n49815), .I1(n60[13]), 
            .CO(n36048));
    SB_LUT4 add_3058_16_lut (.I0(GND_net), .I1(n8104[13]), .I2(GND_net), 
            .I3(n37220), .O(n8076[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_16 (.CI(n37220), .I0(n8104[13]), .I1(GND_net), .CO(n37221));
    SB_LUT4 unary_minus_23_add_3_14_lut (.I0(\PID_CONTROLLER.result [12]), 
            .I1(n49815), .I2(n60[12]), .I3(n36046), .O(n459)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3340_8 (.CI(n36432), .I0(n14910[5]), .I1(n545), .CO(n36433));
    SB_CARRY unary_minus_23_add_3_14 (.CI(n36046), .I0(n49815), .I1(n60[12]), 
            .CO(n36047));
    SB_LUT4 unary_minus_23_add_3_13_lut (.I0(\PID_CONTROLLER.result [11]), 
            .I1(n49815), .I2(n60[11]), .I3(n36045), .O(n460)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mult_14_add_1216_19 (.CI(n37768), .I0(n1802[16]), .I1(GND_net), 
            .CO(n37769));
    SB_CARRY mult_14_add_1212_14 (.CI(n37671), .I0(n1798[11]), .I1(GND_net), 
            .CO(n37672));
    SB_LUT4 add_3058_15_lut (.I0(GND_net), .I1(n8104[12]), .I2(GND_net), 
            .I3(n37219), .O(n8076[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_4 (.CI(n37600), .I0(n15638[1]), .I1(n337), .CO(n37601));
    SB_LUT4 add_3078_8_lut (.I0(GND_net), .I1(n8470[5]), .I2(n545), .I3(n37522), 
            .O(n8446[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_14_lut (.I0(GND_net), .I1(n8311[11]), .I2(GND_net), 
            .I3(n37407), .O(n8292[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_15 (.CI(n37219), .I0(n8104[12]), .I1(GND_net), .CO(n37220));
    SB_LUT4 add_3058_14_lut (.I0(GND_net), .I1(n8104[11]), .I2(GND_net), 
            .I3(n37218), .O(n8076[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_8 (.CI(n37522), .I0(n8470[5]), .I1(n545), .CO(n37523));
    SB_CARRY add_3067_14 (.CI(n37407), .I0(n8311[11]), .I1(GND_net), .CO(n37408));
    SB_CARRY add_3058_14 (.CI(n37218), .I0(n8104[11]), .I1(GND_net), .CO(n37219));
    SB_LUT4 add_3058_13_lut (.I0(GND_net), .I1(n8104[10]), .I2(GND_net), 
            .I3(n37217), .O(n8076[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3387_3_lut (.I0(GND_net), .I1(n15638[0]), .I2(n240), .I3(n37599), 
            .O(n15397[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_7_lut (.I0(GND_net), .I1(n8470[4]), .I2(n472), .I3(n37521), 
            .O(n8446[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_18_lut (.I0(GND_net), .I1(n1802[15]), .I2(GND_net), 
            .I3(n37767), .O(n1801[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_18 (.CI(n37767), .I0(n1802[15]), .I1(GND_net), 
            .CO(n37768));
    SB_LUT4 add_3067_13_lut (.I0(GND_net), .I1(n8311[10]), .I2(GND_net), 
            .I3(n37406), .O(n8292[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_13 (.CI(n37217), .I0(n8104[10]), .I1(GND_net), .CO(n37218));
    SB_LUT4 add_3058_12_lut (.I0(GND_net), .I1(n8104[9]), .I2(GND_net), 
            .I3(n37216), .O(n8076[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_7 (.CI(n37521), .I0(n8470[4]), .I1(n472), .CO(n37522));
    SB_CARRY add_3067_13 (.CI(n37406), .I0(n8311[10]), .I1(GND_net), .CO(n37407));
    SB_CARRY add_3058_12 (.CI(n37216), .I0(n8104[9]), .I1(GND_net), .CO(n37217));
    SB_LUT4 add_3058_11_lut (.I0(GND_net), .I1(n8104[8]), .I2(GND_net), 
            .I3(n37215), .O(n8076[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_3 (.CI(n37599), .I0(n15638[0]), .I1(n240), .CO(n37600));
    SB_LUT4 add_3078_6_lut (.I0(GND_net), .I1(n8470[3]), .I2(n399_c), 
            .I3(n37520), .O(n8446[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_12_lut (.I0(GND_net), .I1(n8311[9]), .I2(GND_net), 
            .I3(n37405), .O(n8292[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_6 (.CI(n37520), .I0(n8470[3]), .I1(n399_c), .CO(n37521));
    SB_CARRY add_3067_12 (.CI(n37405), .I0(n8311[9]), .I1(GND_net), .CO(n37406));
    SB_CARRY add_3058_11 (.CI(n37215), .I0(n8104[8]), .I1(GND_net), .CO(n37216));
    SB_LUT4 mult_14_add_1212_13_lut (.I0(GND_net), .I1(n1798[10]), .I2(GND_net), 
            .I3(n37670), .O(n1797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3387_2_lut (.I0(GND_net), .I1(n50_adj_3379), .I2(n143_adj_3380), 
            .I3(GND_net), .O(n15397[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_10_lut (.I0(GND_net), .I1(n8104[7]), .I2(GND_net), 
            .I3(n37214), .O(n8076[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_5_lut (.I0(GND_net), .I1(n8470[2]), .I2(n326), .I3(n37519), 
            .O(n8446[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_11_lut (.I0(GND_net), .I1(n8311[8]), .I2(GND_net), 
            .I3(n37404), .O(n8292[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_10 (.CI(n37214), .I0(n8104[7]), .I1(GND_net), .CO(n37215));
    SB_LUT4 add_3058_9_lut (.I0(GND_net), .I1(n8104[6]), .I2(GND_net), 
            .I3(n37213), .O(n8076[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3340_7_lut (.I0(GND_net), .I1(n14910[4]), .I2(n472), .I3(n36431), 
            .O(n14558[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n36959), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_9 (.CI(n37213), .I0(n8104[6]), .I1(GND_net), .CO(n37214));
    SB_CARRY add_3078_5 (.CI(n37519), .I0(n8470[2]), .I1(n326), .CO(n37520));
    SB_LUT4 add_3058_8_lut (.I0(GND_net), .I1(n8104[5]), .I2(n695), .I3(n37212), 
            .O(n8076[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_11 (.CI(n37404), .I0(n8311[8]), .I1(GND_net), .CO(n37405));
    SB_CARRY add_3058_8 (.CI(n37212), .I0(n8104[5]), .I1(n695), .CO(n37213));
    SB_LUT4 add_3058_7_lut (.I0(GND_net), .I1(n8104[4]), .I2(n598), .I3(n37211), 
            .O(n8076[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31530_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [28]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(n47842), .O(n47091));
    defparam i31530_4_lut.LUT_INIT = 16'h5adb;
    SB_CARRY add_3387_2 (.CI(GND_net), .I0(n50_adj_3379), .I1(n143_adj_3380), 
            .CO(n37599));
    SB_LUT4 add_3078_4_lut (.I0(GND_net), .I1(n8470[1]), .I2(n253), .I3(n37518), 
            .O(n8446[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_10_lut (.I0(GND_net), .I1(n8311[7]), .I2(GND_net), 
            .I3(n37403), .O(n8292[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_13 (.CI(n36045), .I0(n49815), .I1(n60[11]), 
            .CO(n36046));
    SB_CARRY add_3340_7 (.CI(n36431), .I0(n14910[4]), .I1(n472), .CO(n36432));
    SB_CARRY add_3058_7 (.CI(n37211), .I0(n8104[4]), .I1(n598), .CO(n37212));
    SB_LUT4 unary_minus_23_add_3_12_lut (.I0(\PID_CONTROLLER.result [10]), 
            .I1(n49815), .I2(n60[10]), .I3(n36044), .O(n461)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_13_add_1_21902_add_1_29_lut (.I0(GND_net), .I1(n7063[4]), 
            .I2(n58[27]), .I3(n35913), .O(n57[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3340_6_lut (.I0(GND_net), .I1(n14910[3]), .I2(n399_c), 
            .I3(n36430), .O(n14558[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_10 (.CI(n37403), .I0(n8311[7]), .I1(GND_net), .CO(n37404));
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n36958), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_10  (.CI(n36958), .I0(\PID_CONTROLLER.err[8] ), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n36959));
    SB_LUT4 add_3058_6_lut (.I0(GND_net), .I1(n8104[3]), .I2(n501), .I3(n37210), 
            .O(n8076[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_12 (.CI(n36044), .I0(n49815), .I1(n60[10]), 
            .CO(n36045));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i61_rep_252_2_lut  (.I0(deadband[23]), 
            .I1(\PID_CONTROLLER.result [30]), .I2(GND_net), .I3(GND_net), 
            .O(n50234));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i61_rep_252_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 i15489_1_lut (.I0(\PID_CONTROLLER.result [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28894));   // verilog/motorControl.v(38[14] 59[8])
    defparam i15489_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_13_add_1_21902_add_1_29 (.CI(n35913), .I0(n7063[4]), .I1(n58[27]), 
            .CO(n35914));
    SB_LUT4 add_3067_9_lut (.I0(GND_net), .I1(n8311[6]), .I2(GND_net), 
            .I3(n37402), .O(n8292[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n36957), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_11_lut (.I0(\PID_CONTROLLER.result [9]), 
            .I1(n49815), .I2(n60[9]), .I3(n36043), .O(n462)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_9  (.CI(n36957), .I0(\PID_CONTROLLER.err[7] ), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n36958));
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n36956), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_11 (.CI(n36043), .I0(n49815), .I1(n60[9]), 
            .CO(n36044));
    SB_CARRY add_3058_6 (.CI(n37210), .I0(n8104[3]), .I1(n501), .CO(n37211));
    SB_LUT4 i32926_3_lut (.I0(n54), .I1(n18), .I2(n47822), .I3(GND_net), 
            .O(n48487));   // verilog/motorControl.v(44[10:27])
    defparam i32926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mult_14_add_1216_17_lut (.I0(GND_net), .I1(n1802[14]), .I2(GND_net), 
            .I3(n37766), .O(n1801[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_17 (.CI(n37766), .I0(n1802[14]), .I1(GND_net), 
            .CO(n37767));
    SB_LUT4 mult_14_add_1216_16_lut (.I0(GND_net), .I1(n1802[13]), .I2(GND_net), 
            .I3(n37765), .O(n1801[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3340_6 (.CI(n36430), .I0(n14910[3]), .I1(n399_c), .CO(n36431));
    SB_CARRY add_3067_9 (.CI(n37402), .I0(n8311[6]), .I1(GND_net), .CO(n37403));
    SB_LUT4 add_3058_5_lut (.I0(GND_net), .I1(n8104[2]), .I2(n404), .I3(n37209), 
            .O(n8076[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3340_5_lut (.I0(GND_net), .I1(n14910[2]), .I2(n326), .I3(n36429), 
            .O(n14558[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_10_lut (.I0(\PID_CONTROLLER.result [8]), 
            .I1(n49815), .I2(n60[8]), .I3(n36042), .O(n463)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3340_5 (.CI(n36429), .I0(n14910[2]), .I1(n326), .CO(n36430));
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_8  (.CI(n36956), .I0(\PID_CONTROLLER.err[6] ), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n36957));
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n36955), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_5 (.CI(n37209), .I0(n8104[2]), .I1(n404), .CO(n37210));
    SB_LUT4 add_3340_4_lut (.I0(GND_net), .I1(n14910[1]), .I2(n253), .I3(n36428), 
            .O(n14558[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_10 (.CI(n36042), .I0(n49815), .I1(n60[8]), 
            .CO(n36043));
    SB_CARRY add_3340_4 (.CI(n36428), .I0(n14910[1]), .I1(n253), .CO(n36429));
    SB_LUT4 add_3340_3_lut (.I0(GND_net), .I1(n14910[0]), .I2(n180), .I3(n36427), 
            .O(n14558[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_9_lut (.I0(\PID_CONTROLLER.result[7] ), .I1(n49815), 
            .I2(n60[7]), .I3(n36041), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3340_3 (.CI(n36427), .I0(n14910[0]), .I1(n180), .CO(n36428));
    SB_CARRY unary_minus_23_add_3_9 (.CI(n36041), .I0(n49815), .I1(n60[7]), 
            .CO(n36042));
    SB_LUT4 unary_minus_23_add_3_8_lut (.I0(\PID_CONTROLLER.result [6]), .I1(n49815), 
            .I2(n60[6]), .I3(n36040), .O(n465)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i32101_4_lut (.I0(n48461), .I1(\PID_CONTROLLER.result [28]), 
            .I2(deadband[23]), .I3(\PID_CONTROLLER.result [27]), .O(n47662));   // verilog/motorControl.v(44[10:27])
    defparam i32101_4_lut.LUT_INIT = 16'h8f0e;
    SB_CARRY mult_14_add_1216_16 (.CI(n37765), .I0(n1802[13]), .I1(GND_net), 
            .CO(n37766));
    SB_LUT4 mult_14_add_1216_15_lut (.I0(GND_net), .I1(n1802[12]), .I2(GND_net), 
            .I3(n37764), .O(n1801[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_15 (.CI(n37764), .I0(n1802[12]), .I1(GND_net), 
            .CO(n37765));
    SB_CARRY mult_14_add_1212_13 (.CI(n37670), .I0(n1798[10]), .I1(GND_net), 
            .CO(n37671));
    SB_LUT4 add_3487_7_lut (.I0(GND_net), .I1(n43968), .I2(n658), .I3(n37598), 
            .O(n16627[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3487_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_4 (.CI(n37518), .I0(n8470[1]), .I1(n253), .CO(n37519));
    SB_LUT4 add_3067_8_lut (.I0(GND_net), .I1(n8311[5]), .I2(n722), .I3(n37401), 
            .O(n8292[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_4_lut (.I0(GND_net), .I1(n8104[1]), .I2(n307), .I3(n37208), 
            .O(n8076[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_4 (.CI(n37208), .I0(n8104[1]), .I1(n307), .CO(n37209));
    SB_LUT4 add_3078_3_lut (.I0(GND_net), .I1(n8470[0]), .I2(n180), .I3(n37517), 
            .O(n8446[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_8 (.CI(n37401), .I0(n8311[5]), .I1(n722), .CO(n37402));
    SB_LUT4 add_3058_3_lut (.I0(GND_net), .I1(n8104[0]), .I2(n210), .I3(n37207), 
            .O(n8076[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_3 (.CI(n37207), .I0(n8104[0]), .I1(n210), .CO(n37208));
    SB_LUT4 add_3487_6_lut (.I0(GND_net), .I1(n16635[3]), .I2(n558), .I3(n37597), 
            .O(n16627[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3487_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_3 (.CI(n37517), .I0(n8470[0]), .I1(n180), .CO(n37518));
    SB_LUT4 add_3067_7_lut (.I0(GND_net), .I1(n8311[4]), .I2(n625), .I3(n37400), 
            .O(n8292[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_2_lut (.I0(GND_net), .I1(n20_adj_3384), .I2(n113), 
            .I3(GND_net), .O(n8076[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_2 (.CI(GND_net), .I0(n20_adj_3384), .I1(n113), .CO(n37207));
    SB_LUT4 add_3078_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n8446[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_7 (.CI(n37400), .I0(n8311[4]), .I1(n625), .CO(n37401));
    SB_LUT4 add_3057_28_lut (.I0(GND_net), .I1(n8076[25]), .I2(GND_net), 
            .I3(n37206), .O(n8047[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_27_lut (.I0(GND_net), .I1(n8076[24]), .I2(GND_net), 
            .I3(n37205), .O(n8047[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_12_lut (.I0(GND_net), .I1(n1798[9]), .I2(GND_net), 
            .I3(n37669), .O(n1797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3487_6 (.CI(n37597), .I0(n16635[3]), .I1(n558), .CO(n37598));
    SB_CARRY add_3078_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n37517));
    SB_LUT4 add_3067_6_lut (.I0(GND_net), .I1(n8311[3]), .I2(n528), .I3(n37399), 
            .O(n8292[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_27 (.CI(n37205), .I0(n8076[24]), .I1(GND_net), .CO(n37206));
    SB_LUT4 add_3057_26_lut (.I0(GND_net), .I1(n8076[23]), .I2(GND_net), 
            .I3(n37204), .O(n8047[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_8_lut (.I0(GND_net), .I1(n9317[5]), .I2(n752), .I3(n37516), 
            .O(n8437[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_12 (.CI(n37669), .I0(n1798[9]), .I1(GND_net), 
            .CO(n37670));
    SB_LUT4 sub_11_inv_0_i7_1_lut (.I0(\PID_CONTROLLER.err[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[6]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3067_6 (.CI(n37399), .I0(n8311[3]), .I1(n528), .CO(n37400));
    SB_CARRY add_3057_26 (.CI(n37204), .I0(n8076[23]), .I1(GND_net), .CO(n37205));
    SB_LUT4 add_3057_25_lut (.I0(GND_net), .I1(n8076[22]), .I2(GND_net), 
            .I3(n37203), .O(n8047[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3487_5_lut (.I0(GND_net), .I1(n16635[2]), .I2(n464), .I3(n37596), 
            .O(n16627[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3487_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_7_lut (.I0(GND_net), .I1(n9317[4]), .I2(n655), .I3(n37515), 
            .O(n8437[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3067_5_lut (.I0(GND_net), .I1(n8311[2]), .I2(n431), .I3(n37398), 
            .O(n8292[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_11_lut (.I0(GND_net), .I1(n1798[8]), .I2(GND_net), 
            .I3(n37668), .O(n1797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_25 (.CI(n37203), .I0(n8076[22]), .I1(GND_net), .CO(n37204));
    SB_LUT4 add_3057_24_lut (.I0(GND_net), .I1(n8076[21]), .I2(GND_net), 
            .I3(n37202), .O(n8047[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_7 (.CI(n37515), .I0(n9317[4]), .I1(n655), .CO(n37516));
    SB_LUT4 add_3077_6_lut (.I0(GND_net), .I1(n9317[3]), .I2(n558_adj_3386), 
            .I3(n37514), .O(n8437[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_5 (.CI(n37398), .I0(n8311[2]), .I1(n431), .CO(n37399));
    SB_CARRY add_3487_5 (.CI(n37596), .I0(n16635[2]), .I1(n464), .CO(n37597));
    SB_LUT4 add_13_add_1_21902_add_1_28_lut (.I0(GND_net), .I1(n7063[3]), 
            .I2(n58[26]), .I3(n35912), .O(n57[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_24 (.CI(n37202), .I0(n8076[21]), .I1(GND_net), .CO(n37203));
    SB_LUT4 i33319_3_lut (.I0(n48879), .I1(\PID_CONTROLLER.result [23]), 
            .I2(deadband[23]), .I3(GND_net), .O(n48880));   // verilog/motorControl.v(44[10:27])
    defparam i33319_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_14_add_1216_14_lut (.I0(GND_net), .I1(n1802[11]), .I2(GND_net), 
            .I3(n37763), .O(n1801[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_11 (.CI(n37668), .I0(n1798[8]), .I1(GND_net), 
            .CO(n37669));
    SB_LUT4 add_3487_4_lut (.I0(GND_net), .I1(n16635[1]), .I2(n370), .I3(n37595), 
            .O(n16627[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3487_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_6 (.CI(n37514), .I0(n9317[3]), .I1(n558_adj_3386), 
            .CO(n37515));
    SB_LUT4 add_3067_4_lut (.I0(GND_net), .I1(n8311[1]), .I2(n334), .I3(n37397), 
            .O(n8292[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33031_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [28]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(n47848), .O(n48592));
    defparam i33031_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 add_3077_5_lut (.I0(GND_net), .I1(n9317[2]), .I2(n461_adj_3387), 
            .I3(n37513), .O(n8437[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_4 (.CI(n37397), .I0(n8311[1]), .I1(n334), .CO(n37398));
    SB_CARRY add_3487_4 (.CI(n37595), .I0(n16635[1]), .I1(n370), .CO(n37596));
    SB_CARRY add_3077_5 (.CI(n37513), .I0(n9317[2]), .I1(n461_adj_3387), 
            .CO(n37514));
    SB_LUT4 add_3067_3_lut (.I0(GND_net), .I1(n8311[0]), .I2(n237), .I3(n37396), 
            .O(n8292[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_4_lut (.I0(GND_net), .I1(n9317[1]), .I2(n364), .I3(n37512), 
            .O(n8437[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_14 (.CI(n37763), .I0(n1802[11]), .I1(GND_net), 
            .CO(n37764));
    SB_LUT4 mult_14_add_1216_13_lut (.I0(GND_net), .I1(n1802[10]), .I2(GND_net), 
            .I3(n37762), .O(n1801[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_13 (.CI(n37762), .I0(n1802[10]), .I1(GND_net), 
            .CO(n37763));
    SB_CARRY add_3067_3 (.CI(n37396), .I0(n8311[0]), .I1(n237), .CO(n37397));
    SB_LUT4 mult_14_add_1212_10_lut (.I0(GND_net), .I1(n1798[7]), .I2(GND_net), 
            .I3(n37667), .O(n1797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3487_3_lut (.I0(GND_net), .I1(n16635[0]), .I2(n276), .I3(n37594), 
            .O(n16627[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3487_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_4 (.CI(n37512), .I0(n9317[1]), .I1(n364), .CO(n37513));
    SB_LUT4 add_3067_2_lut (.I0(GND_net), .I1(n47_adj_3388), .I2(n140), 
            .I3(GND_net), .O(n8292[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3067_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_3_lut (.I0(GND_net), .I1(n9317[0]), .I2(n267), .I3(n37511), 
            .O(n8437[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3067_2 (.CI(GND_net), .I0(n47_adj_3388), .I1(n140), .CO(n37396));
    SB_CARRY add_3487_3 (.CI(n37594), .I0(n16635[0]), .I1(n276), .CO(n37595));
    SB_CARRY add_3077_3 (.CI(n37511), .I0(n9317[0]), .I1(n267), .CO(n37512));
    SB_LUT4 add_3066_19_lut (.I0(GND_net), .I1(n8292[16]), .I2(GND_net), 
            .I3(n37395), .O(n8272[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_2_lut (.I0(GND_net), .I1(n86), .I2(n170), .I3(GND_net), 
            .O(n8437[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_18_lut (.I0(GND_net), .I1(n8292[15]), .I2(GND_net), 
            .I3(n37394), .O(n8272[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3487_2_lut (.I0(GND_net), .I1(n86_adj_3389), .I2(n182), 
            .I3(GND_net), .O(n16627[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3487_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_12_lut (.I0(GND_net), .I1(n1802[9]), .I2(GND_net), 
            .I3(n37761), .O(n1801[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_10 (.CI(n37667), .I0(n1798[7]), .I1(GND_net), 
            .CO(n37668));
    SB_CARRY add_3487_2 (.CI(GND_net), .I0(n86_adj_3389), .I1(n182), .CO(n37594));
    SB_CARRY add_3077_2 (.CI(GND_net), .I0(n86), .I1(n170), .CO(n37511));
    SB_CARRY add_3066_18 (.CI(n37394), .I0(n8292[15]), .I1(GND_net), .CO(n37395));
    SB_LUT4 add_3057_23_lut (.I0(GND_net), .I1(n8076[20]), .I2(GND_net), 
            .I3(n37201), .O(n8047[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_17_lut (.I0(GND_net), .I1(n8292[14]), .I2(GND_net), 
            .I3(n37393), .O(n8272[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33356_4_lut (.I0(n47662), .I1(n48487), .I2(n50234), .I3(n47091), 
            .O(n48917));   // verilog/motorControl.v(44[10:27])
    defparam i33356_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3057_23 (.CI(n37201), .I0(n8076[20]), .I1(GND_net), .CO(n37202));
    SB_LUT4 add_3402_16_lut (.I0(GND_net), .I1(n15848[13]), .I2(GND_net), 
            .I3(n37593), .O(n15638[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_9_lut (.I0(GND_net), .I1(n8437[6]), .I2(GND_net), 
            .I3(n37510), .O(n8427[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_7  (.CI(n36955), .I0(\PID_CONTROLLER.err[5] ), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n36956));
    SB_LUT4 add_3402_15_lut (.I0(GND_net), .I1(n15848[12]), .I2(GND_net), 
            .I3(n37592), .O(n15638[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_22_lut (.I0(GND_net), .I1(n8076[19]), .I2(GND_net), 
            .I3(n37200), .O(n8047[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n36954), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_8_lut (.I0(GND_net), .I1(n8437[5]), .I2(n749), .I3(n37509), 
            .O(n8427[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_8 (.CI(n36040), .I0(n49815), .I1(n60[6]), 
            .CO(n36041));
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_6  (.CI(n36954), .I0(\PID_CONTROLLER.err[4] ), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n36955));
    SB_LUT4 i32099_4_lut (.I0(n48880), .I1(\PID_CONTROLLER.result [25]), 
            .I2(deadband[23]), .I3(\PID_CONTROLLER.result [24]), .O(n47660));   // verilog/motorControl.v(44[10:27])
    defparam i32099_4_lut.LUT_INIT = 16'h8f0e;
    SB_CARRY add_3076_8 (.CI(n37509), .I0(n8437[5]), .I1(n749), .CO(n37510));
    SB_LUT4 i2_4_lut (.I0(\PID_CONTROLLER.result [29]), .I1(\PID_CONTROLLER.result [26]), 
            .I2(pwm_23__N_2960[24]), .I3(\PID_CONTROLLER.result [25]), .O(n43891));   // verilog/motorControl.v(44[31:51])
    defparam i2_4_lut.LUT_INIT = 16'h7ffe;
    SB_CARRY add_3066_17 (.CI(n37393), .I0(n8292[14]), .I1(GND_net), .CO(n37394));
    SB_CARRY add_3057_22 (.CI(n37200), .I0(n8076[19]), .I1(GND_net), .CO(n37201));
    SB_LUT4 add_3057_21_lut (.I0(GND_net), .I1(n8076[18]), .I2(GND_net), 
            .I3(n37199), .O(n8047[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_16_lut (.I0(GND_net), .I1(n8292[13]), .I2(GND_net), 
            .I3(n37392), .O(n8272[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_21 (.CI(n37199), .I0(n8076[18]), .I1(GND_net), .CO(n37200));
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n36953), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_5  (.CI(n36953), .I0(\PID_CONTROLLER.err[3] ), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n36954));
    SB_LUT4 add_3057_20_lut (.I0(GND_net), .I1(n8076[17]), .I2(GND_net), 
            .I3(n37198), .O(n8047[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n36952), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_4  (.CI(n36952), .I0(\PID_CONTROLLER.err[2] ), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n36953));
    SB_CARRY add_3402_15 (.CI(n37592), .I0(n15848[12]), .I1(GND_net), 
            .CO(n37593));
    SB_LUT4 add_3076_7_lut (.I0(GND_net), .I1(n8437[4]), .I2(n652), .I3(n37508), 
            .O(n8427[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_16 (.CI(n37392), .I0(n8292[13]), .I1(GND_net), .CO(n37393));
    SB_CARRY add_3057_20 (.CI(n37198), .I0(n8076[17]), .I1(GND_net), .CO(n37199));
    SB_LUT4 add_3057_19_lut (.I0(GND_net), .I1(n8076[16]), .I2(GND_net), 
            .I3(n37197), .O(n8047[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_15_lut (.I0(GND_net), .I1(n8292[12]), .I2(GND_net), 
            .I3(n37391), .O(n8272[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_15 (.CI(n37391), .I0(n8292[12]), .I1(GND_net), .CO(n37392));
    SB_CARRY add_3057_19 (.CI(n37197), .I0(n8076[16]), .I1(GND_net), .CO(n37198));
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n36951), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_3  (.CI(n36951), .I0(\PID_CONTROLLER.err[1] ), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n36952));
    SB_LUT4 add_3057_18_lut (.I0(GND_net), .I1(n8076[15]), .I2(GND_net), 
            .I3(n37196), .O(n8047[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1015_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1015_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1015_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err[0] ), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n36951));
    SB_CARRY add_3076_7 (.CI(n37508), .I0(n8437[4]), .I1(n652), .CO(n37509));
    SB_LUT4 add_3066_14_lut (.I0(GND_net), .I1(n8292[11]), .I2(GND_net), 
            .I3(n37390), .O(n8272[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_18 (.CI(n37196), .I0(n8076[15]), .I1(GND_net), .CO(n37197));
    SB_LUT4 add_3057_17_lut (.I0(GND_net), .I1(n8076[14]), .I2(GND_net), 
            .I3(n37195), .O(n8047[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_14 (.CI(n37390), .I0(n8292[11]), .I1(GND_net), .CO(n37391));
    SB_CARRY add_3057_17 (.CI(n37195), .I0(n8076[14]), .I1(GND_net), .CO(n37196));
    SB_LUT4 pwm_count_1014_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[8]), 
            .I3(n36950), .O(n64[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1014_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[7]), 
            .I3(n36949), .O(n64[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_16_lut (.I0(GND_net), .I1(n8076[13]), .I2(GND_net), 
            .I3(n37194), .O(n8047[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1014_add_4_9 (.CI(n36949), .I0(GND_net), .I1(pwm_count[7]), 
            .CO(n36950));
    SB_LUT4 pwm_count_1014_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[6]), 
            .I3(n36948), .O(n64[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_9_lut (.I0(GND_net), .I1(n1798[6]), .I2(GND_net), 
            .I3(n37666), .O(n1797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3402_14_lut (.I0(GND_net), .I1(n15848[11]), .I2(GND_net), 
            .I3(n37591), .O(n15638[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_6_lut (.I0(GND_net), .I1(n8437[3]), .I2(n555), .I3(n37507), 
            .O(n8427[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_13_lut (.I0(GND_net), .I1(n8292[10]), .I2(GND_net), 
            .I3(n37389), .O(n8272[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_16 (.CI(n37194), .I0(n8076[13]), .I1(GND_net), .CO(n37195));
    SB_LUT4 add_3057_15_lut (.I0(GND_net), .I1(n8076[12]), .I2(GND_net), 
            .I3(n37193), .O(n8047[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_13 (.CI(n37389), .I0(n8292[10]), .I1(GND_net), .CO(n37390));
    SB_CARRY add_3057_15 (.CI(n37193), .I0(n8076[12]), .I1(GND_net), .CO(n37194));
    SB_CARRY pwm_count_1014_add_4_8 (.CI(n36948), .I0(GND_net), .I1(pwm_count[6]), 
            .CO(n36949));
    SB_LUT4 pwm_count_1014_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[5]), 
            .I3(n36947), .O(n64[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_14_lut (.I0(GND_net), .I1(n8076[11]), .I2(GND_net), 
            .I3(n37192), .O(n8047[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1014_add_4_7 (.CI(n36947), .I0(GND_net), .I1(pwm_count[5]), 
            .CO(n36948));
    SB_LUT4 pwm_count_1014_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[4]), 
            .I3(n36946), .O(n64[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_6 (.CI(n37507), .I0(n8437[3]), .I1(n555), .CO(n37508));
    SB_LUT4 add_3066_12_lut (.I0(GND_net), .I1(n8292[9]), .I2(GND_net), 
            .I3(n37388), .O(n8272[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_14 (.CI(n37192), .I0(n8076[11]), .I1(GND_net), .CO(n37193));
    SB_LUT4 add_3057_13_lut (.I0(GND_net), .I1(n8076[10]), .I2(GND_net), 
            .I3(n37191), .O(n8047[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_12 (.CI(n37388), .I0(n8292[9]), .I1(GND_net), .CO(n37389));
    SB_CARRY add_3057_13 (.CI(n37191), .I0(n8076[10]), .I1(GND_net), .CO(n37192));
    SB_CARRY pwm_count_1014_add_4_6 (.CI(n36946), .I0(GND_net), .I1(pwm_count[4]), 
            .CO(n36947));
    SB_LUT4 pwm_count_1014_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[3]), 
            .I3(n36945), .O(n64[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_12_lut (.I0(GND_net), .I1(n8076[9]), .I2(GND_net), 
            .I3(n37190), .O(n8047[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1014_add_4_5 (.CI(n36945), .I0(GND_net), .I1(pwm_count[3]), 
            .CO(n36946));
    SB_LUT4 pwm_count_1014_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[2]), 
            .I3(n36944), .O(n64[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_14 (.CI(n37591), .I0(n15848[11]), .I1(GND_net), 
            .CO(n37592));
    SB_LUT4 add_3076_5_lut (.I0(GND_net), .I1(n8437[2]), .I2(n458), .I3(n37506), 
            .O(n8427[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_23__I_819_i4_3_lut (.I0(n46591), .I1(pwm_23__N_2960[1]), 
            .I2(\PID_CONTROLLER.result [1]), .I3(GND_net), .O(n4));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3066_11_lut (.I0(GND_net), .I1(n8292[8]), .I2(GND_net), 
            .I3(n37387), .O(n8272[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_12 (.CI(n37190), .I0(n8076[9]), .I1(GND_net), .CO(n37191));
    SB_LUT4 add_3057_11_lut (.I0(GND_net), .I1(n8076[8]), .I2(GND_net), 
            .I3(n37189), .O(n8047[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_11 (.CI(n37387), .I0(n8292[8]), .I1(GND_net), .CO(n37388));
    SB_CARRY add_3057_11 (.CI(n37189), .I0(n8076[8]), .I1(GND_net), .CO(n37190));
    SB_LUT4 i32896_3_lut (.I0(n4), .I1(\pwm_23__N_2960[13] ), .I2(\PID_CONTROLLER.result[13] ), 
            .I3(GND_net), .O(n48457));   // verilog/motorControl.v(44[31:51])
    defparam i32896_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY pwm_count_1014_add_4_4 (.CI(n36944), .I0(GND_net), .I1(pwm_count[2]), 
            .CO(n36945));
    SB_LUT4 pwm_count_1014_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[1]), 
            .I3(n36943), .O(n64[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_10_lut (.I0(GND_net), .I1(n8076[7]), .I2(GND_net), 
            .I3(n37188), .O(n8047[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1014_add_4_3 (.CI(n36943), .I0(GND_net), .I1(pwm_count[1]), 
            .CO(n36944));
    SB_LUT4 pwm_count_1014_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[0]), 
            .I3(VCC_net), .O(n64[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1014_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3076_5 (.CI(n37506), .I0(n8437[2]), .I1(n458), .CO(n37507));
    SB_LUT4 add_3066_10_lut (.I0(GND_net), .I1(n8292[7]), .I2(GND_net), 
            .I3(n37386), .O(n8272[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_10 (.CI(n37188), .I0(n8076[7]), .I1(GND_net), .CO(n37189));
    SB_LUT4 add_3057_9_lut (.I0(GND_net), .I1(n8076[6]), .I2(GND_net), 
            .I3(n37187), .O(n8047[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_10 (.CI(n37386), .I0(n8292[7]), .I1(GND_net), .CO(n37387));
    SB_CARRY add_3057_9 (.CI(n37187), .I0(n8076[6]), .I1(GND_net), .CO(n37188));
    SB_CARRY pwm_count_1014_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_count[0]), 
            .CO(n36943));
    SB_LUT4 add_3054_31_lut (.I0(GND_net), .I1(n7986[28]), .I2(GND_net), 
            .I3(n36942), .O(n7954[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3057_8_lut (.I0(GND_net), .I1(n8076[5]), .I2(n692), .I3(n37186), 
            .O(n8047[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3054_30_lut (.I0(GND_net), .I1(n7986[27]), .I2(GND_net), 
            .I3(n36941), .O(n7954[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_12 (.CI(n37761), .I0(n1802[9]), .I1(GND_net), 
            .CO(n37762));
    SB_CARRY mult_14_add_1212_9 (.CI(n37666), .I0(n1798[6]), .I1(GND_net), 
            .CO(n37667));
    SB_LUT4 add_3402_13_lut (.I0(GND_net), .I1(n15848[10]), .I2(GND_net), 
            .I3(n37590), .O(n15638[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_4_lut (.I0(GND_net), .I1(n8437[1]), .I2(n361), .I3(n37505), 
            .O(n8427[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_9_lut (.I0(GND_net), .I1(n8292[6]), .I2(GND_net), 
            .I3(n37385), .O(n8272[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_8 (.CI(n37186), .I0(n8076[5]), .I1(n692), .CO(n37187));
    SB_CARRY add_3066_9 (.CI(n37385), .I0(n8292[6]), .I1(GND_net), .CO(n37386));
    SB_LUT4 add_3057_7_lut (.I0(GND_net), .I1(n8076[4]), .I2(n595), .I3(n37185), 
            .O(n8047[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_30 (.CI(n36941), .I0(n7986[27]), .I1(GND_net), .CO(n36942));
    SB_LUT4 add_3340_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n14558[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3057_7 (.CI(n37185), .I0(n8076[4]), .I1(n595), .CO(n37186));
    SB_CARRY add_3340_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n36427));
    SB_LUT4 add_3195_26_lut (.I0(GND_net), .I1(n11990[23]), .I2(GND_net), 
            .I3(n36426), .O(n11356[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_25_lut (.I0(GND_net), .I1(n11990[22]), .I2(GND_net), 
            .I3(n36425), .O(n11356[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_25 (.CI(n36425), .I0(n11990[22]), .I1(GND_net), 
            .CO(n36426));
    SB_CARRY add_3076_4 (.CI(n37505), .I0(n8437[1]), .I1(n361), .CO(n37506));
    SB_LUT4 add_3066_8_lut (.I0(GND_net), .I1(n8292[5]), .I2(n719), .I3(n37384), 
            .O(n8272[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_8 (.CI(n37384), .I0(n8292[5]), .I1(n719), .CO(n37385));
    SB_LUT4 unary_minus_23_add_3_7_lut (.I0(\PID_CONTROLLER.result[5] ), .I1(n49815), 
            .I2(n60[5]), .I3(n36039), .O(n26834)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3057_6_lut (.I0(GND_net), .I1(n8076[3]), .I2(n498), .I3(n37184), 
            .O(n8047[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_24_lut (.I0(GND_net), .I1(n11990[21]), .I2(GND_net), 
            .I3(n36424), .O(n11356[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_24 (.CI(n36424), .I0(n11990[21]), .I1(GND_net), 
            .CO(n36425));
    SB_LUT4 i32897_3_lut (.I0(n48457), .I1(\pwm_23__N_2960[14] ), .I2(\PID_CONTROLLER.result[14] ), 
            .I3(GND_net), .O(n48458));   // verilog/motorControl.v(44[31:51])
    defparam i32897_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3057_6 (.CI(n37184), .I0(n8076[3]), .I1(n498), .CO(n37185));
    SB_LUT4 add_3195_23_lut (.I0(GND_net), .I1(n11990[20]), .I2(GND_net), 
            .I3(n36423), .O(n11356[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_23 (.CI(n36423), .I0(n11990[20]), .I1(GND_net), 
            .CO(n36424));
    SB_LUT4 add_3195_22_lut (.I0(GND_net), .I1(n11990[19]), .I2(GND_net), 
            .I3(n36422), .O(n11356[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_7 (.CI(n36039), .I0(n49815), .I1(n60[5]), 
            .CO(n36040));
    SB_CARRY add_3195_22 (.CI(n36422), .I0(n11990[19]), .I1(GND_net), 
            .CO(n36423));
    SB_LUT4 i31439_4_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n50255), 
            .I2(pwm_23__N_2960[16]), .I3(n47784), .O(n46999));
    defparam i31439_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_3402_13 (.CI(n37590), .I0(n15848[10]), .I1(GND_net), 
            .CO(n37591));
    SB_LUT4 add_3076_3_lut (.I0(GND_net), .I1(n8437[0]), .I2(n264), .I3(n37504), 
            .O(n8427[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_7_lut (.I0(GND_net), .I1(n8292[4]), .I2(n622), .I3(n37383), 
            .O(n8272[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_23__I_819_i35_rep_261_2_lut (.I0(\PID_CONTROLLER.result [17]), 
            .I1(pwm_23__N_2960[17]), .I2(GND_net), .I3(GND_net), .O(n50243));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i35_rep_261_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_add_1216_11_lut (.I0(GND_net), .I1(n1802[8]), .I2(GND_net), 
            .I3(n37760), .O(n1801[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_7 (.CI(n37383), .I0(n8292[4]), .I1(n622), .CO(n37384));
    SB_LUT4 add_3057_5_lut (.I0(GND_net), .I1(n8076[2]), .I2(n401), .I3(n37183), 
            .O(n8047[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_21_lut (.I0(GND_net), .I1(n11990[18]), .I2(GND_net), 
            .I3(n36421), .O(n11356[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_21 (.CI(n36421), .I0(n11990[18]), .I1(GND_net), 
            .CO(n36422));
    SB_CARRY add_3057_5 (.CI(n37183), .I0(n8076[2]), .I1(n401), .CO(n37184));
    SB_LUT4 add_3195_20_lut (.I0(GND_net), .I1(n11990[17]), .I2(GND_net), 
            .I3(n36420), .O(n11356[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33320_4_lut (.I0(n30_c), .I1(n10), .I2(n50243), .I3(n46995), 
            .O(n48881));   // verilog/motorControl.v(44[31:51])
    defparam i33320_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3195_20 (.CI(n36420), .I0(n11990[17]), .I1(GND_net), 
            .CO(n36421));
    SB_LUT4 add_3195_19_lut (.I0(GND_net), .I1(n11990[16]), .I2(GND_net), 
            .I3(n36419), .O(n11356[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_19 (.CI(n36419), .I0(n11990[16]), .I1(GND_net), 
            .CO(n36420));
    SB_CARRY add_3076_3 (.CI(n37504), .I0(n8437[0]), .I1(n264), .CO(n37505));
    SB_LUT4 add_3066_6_lut (.I0(GND_net), .I1(n8292[3]), .I2(n525), .I3(n37382), 
            .O(n8272[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_6 (.CI(n37382), .I0(n8292[3]), .I1(n525), .CO(n37383));
    SB_LUT4 add_3057_4_lut (.I0(GND_net), .I1(n8076[1]), .I2(n304), .I3(n37182), 
            .O(n8047[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_18_lut (.I0(GND_net), .I1(n11990[15]), .I2(GND_net), 
            .I3(n36418), .O(n11356[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_18 (.CI(n36418), .I0(n11990[15]), .I1(GND_net), 
            .CO(n36419));
    SB_CARRY add_3057_4 (.CI(n37182), .I0(n8076[1]), .I1(n304), .CO(n37183));
    SB_LUT4 add_3195_17_lut (.I0(GND_net), .I1(n11990[14]), .I2(GND_net), 
            .I3(n36417), .O(n11356[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_6_lut (.I0(\PID_CONTROLLER.result [4]), .I1(n49815), 
            .I2(n60[4]), .I3(n36038), .O(n467)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_23_add_3_6 (.CI(n36038), .I0(n49815), .I1(n60[4]), 
            .CO(n36039));
    SB_CARRY add_3195_17 (.CI(n36417), .I0(n11990[14]), .I1(GND_net), 
            .CO(n36418));
    SB_LUT4 add_3195_16_lut (.I0(GND_net), .I1(n11990[13]), .I2(GND_net), 
            .I3(n36416), .O(n11356[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_5_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n49815), 
            .I2(n60[3]), .I3(n36037), .O(n468)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_23_add_3_5 (.CI(n36037), .I0(n49815), .I1(n60[3]), 
            .CO(n36038));
    SB_CARRY add_3195_16 (.CI(n36416), .I0(n11990[13]), .I1(GND_net), 
            .CO(n36417));
    SB_LUT4 mult_14_add_1212_8_lut (.I0(GND_net), .I1(n1798[5]), .I2(n515), 
            .I3(n37665), .O(n1797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3402_12_lut (.I0(GND_net), .I1(n15848[9]), .I2(GND_net), 
            .I3(n37589), .O(n15638[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3076_2_lut (.I0(GND_net), .I1(n74), .I2(n167), .I3(GND_net), 
            .O(n8427[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3076_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_5_lut (.I0(GND_net), .I1(n8292[2]), .I2(n428), .I3(n37381), 
            .O(n8272[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_5 (.CI(n37381), .I0(n8292[2]), .I1(n428), .CO(n37382));
    SB_LUT4 add_3057_3_lut (.I0(GND_net), .I1(n8076[0]), .I2(n207), .I3(n37181), 
            .O(n8047[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_15_lut (.I0(GND_net), .I1(n11990[12]), .I2(GND_net), 
            .I3(n36415), .O(n11356[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_15 (.CI(n36415), .I0(n11990[12]), .I1(GND_net), 
            .CO(n36416));
    SB_CARRY add_3057_3 (.CI(n37181), .I0(n8076[0]), .I1(n207), .CO(n37182));
    SB_LUT4 add_3195_14_lut (.I0(GND_net), .I1(n11990[11]), .I2(GND_net), 
            .I3(n36414), .O(n11356[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_14 (.CI(n36414), .I0(n11990[11]), .I1(GND_net), 
            .CO(n36415));
    SB_LUT4 add_3195_13_lut (.I0(GND_net), .I1(n11990[10]), .I2(GND_net), 
            .I3(n36413), .O(n11356[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_13 (.CI(n36413), .I0(n11990[10]), .I1(GND_net), 
            .CO(n36414));
    SB_CARRY add_3076_2 (.CI(GND_net), .I0(n74), .I1(n167), .CO(n37504));
    SB_LUT4 add_3066_4_lut (.I0(GND_net), .I1(n8292[1]), .I2(n331), .I3(n37380), 
            .O(n8272[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32105_3_lut (.I0(n48458), .I1(pwm_23__N_2960[15]), .I2(\PID_CONTROLLER.result [15]), 
            .I3(GND_net), .O(n47666));   // verilog/motorControl.v(44[31:51])
    defparam i32105_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3066_4 (.CI(n37380), .I0(n8292[1]), .I1(n331), .CO(n37381));
    SB_LUT4 add_3057_2_lut (.I0(GND_net), .I1(n17), .I2(n110), .I3(GND_net), 
            .O(n8047[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3057_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_12_lut (.I0(GND_net), .I1(n11990[9]), .I2(GND_net), 
            .I3(n36412), .O(n11356[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_12 (.CI(n36412), .I0(n11990[9]), .I1(GND_net), .CO(n36413));
    SB_CARRY add_3057_2 (.CI(GND_net), .I0(n17), .I1(n110), .CO(n37181));
    SB_LUT4 add_3195_11_lut (.I0(GND_net), .I1(n11990[8]), .I2(GND_net), 
            .I3(n36411), .O(n11356[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_4_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n49815), 
            .I2(n60[2]), .I3(n36036), .O(n469)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3195_11 (.CI(n36411), .I0(n11990[8]), .I1(GND_net), .CO(n36412));
    SB_LUT4 add_3195_10_lut (.I0(GND_net), .I1(n11990[7]), .I2(GND_net), 
            .I3(n36410), .O(n11356[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_4 (.CI(n36036), .I0(n49815), .I1(n60[2]), 
            .CO(n36037));
    SB_CARRY add_3195_10 (.CI(n36410), .I0(n11990[7]), .I1(GND_net), .CO(n36411));
    SB_CARRY add_3402_12 (.CI(n37589), .I0(n15848[9]), .I1(GND_net), .CO(n37590));
    SB_LUT4 add_3075_10_lut (.I0(GND_net), .I1(n8427[7]), .I2(GND_net), 
            .I3(n37503), .O(n8416[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_3_lut (.I0(GND_net), .I1(n8292[0]), .I2(n234), .I3(n37379), 
            .O(n8272[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_3 (.CI(n37379), .I0(n8292[0]), .I1(n234), .CO(n37380));
    SB_LUT4 add_3056_29_lut (.I0(GND_net), .I1(n8047[26]), .I2(GND_net), 
            .I3(n37180), .O(n8017[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_9_lut (.I0(GND_net), .I1(n11990[6]), .I2(GND_net), 
            .I3(n36409), .O(n11356[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_9 (.CI(n36409), .I0(n11990[6]), .I1(GND_net), .CO(n36410));
    SB_LUT4 add_3056_28_lut (.I0(GND_net), .I1(n8047[25]), .I2(GND_net), 
            .I3(n37179), .O(n8017[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_8_lut (.I0(GND_net), .I1(n11990[5]), .I2(n698), .I3(n36408), 
            .O(n11356[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_8 (.CI(n36408), .I0(n11990[5]), .I1(n698), .CO(n36409));
    SB_LUT4 add_3195_7_lut (.I0(GND_net), .I1(n11990[4]), .I2(n601), .I3(n36407), 
            .O(n11356[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_7 (.CI(n36407), .I0(n11990[4]), .I1(n601), .CO(n36408));
    SB_LUT4 add_3075_9_lut (.I0(GND_net), .I1(n8427[6]), .I2(GND_net), 
            .I3(n37502), .O(n8416[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3066_2_lut (.I0(GND_net), .I1(n44_adj_3398), .I2(n137), 
            .I3(GND_net), .O(n8272[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3066_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3066_2 (.CI(GND_net), .I0(n44_adj_3398), .I1(n137), .CO(n37379));
    SB_CARRY add_3056_28 (.CI(n37179), .I0(n8047[25]), .I1(GND_net), .CO(n37180));
    SB_LUT4 add_3195_6_lut (.I0(GND_net), .I1(n11990[3]), .I2(n504), .I3(n36406), 
            .O(n11356[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_6 (.CI(n36406), .I0(n11990[3]), .I1(n504), .CO(n36407));
    SB_LUT4 add_3056_27_lut (.I0(GND_net), .I1(n8047[24]), .I2(GND_net), 
            .I3(n37178), .O(n8017[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_5_lut (.I0(GND_net), .I1(n11990[2]), .I2(n407_c), 
            .I3(n36405), .O(n11356[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_3_lut (.I0(\PID_CONTROLLER.result [1]), .I1(n49815), 
            .I2(n60[1]), .I3(n36035), .O(n470)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_23_add_3_3 (.CI(n36035), .I0(n49815), .I1(n60[1]), 
            .CO(n36036));
    SB_LUT4 i33492_4_lut (.I0(n47666), .I1(n48881), .I2(n50243), .I3(n46999), 
            .O(n49053));   // verilog/motorControl.v(44[31:51])
    defparam i33492_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3195_5 (.CI(n36405), .I0(n11990[2]), .I1(n407_c), .CO(n36406));
    SB_CARRY mult_14_add_1216_11 (.CI(n37760), .I0(n1802[8]), .I1(GND_net), 
            .CO(n37761));
    SB_LUT4 mult_14_add_1216_10_lut (.I0(GND_net), .I1(n1802[7]), .I2(GND_net), 
            .I3(n37759), .O(n1801[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_10 (.CI(n37759), .I0(n1802[7]), .I1(GND_net), 
            .CO(n37760));
    SB_CARRY mult_14_add_1212_8 (.CI(n37665), .I0(n1798[5]), .I1(n515), 
            .CO(n37666));
    SB_LUT4 add_3402_11_lut (.I0(GND_net), .I1(n15848[8]), .I2(GND_net), 
            .I3(n37588), .O(n15638[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_9 (.CI(n37502), .I0(n8427[6]), .I1(GND_net), .CO(n37503));
    SB_LUT4 add_3065_20_lut (.I0(GND_net), .I1(n8272[17]), .I2(GND_net), 
            .I3(n37378), .O(n8251[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33493_3_lut (.I0(n49053), .I1(pwm_23__N_2960[18]), .I2(\PID_CONTROLLER.result [18]), 
            .I3(GND_net), .O(n49054));   // verilog/motorControl.v(44[31:51])
    defparam i33493_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3056_27 (.CI(n37178), .I0(n8047[24]), .I1(GND_net), .CO(n37179));
    SB_LUT4 add_3056_26_lut (.I0(GND_net), .I1(n8047[23]), .I2(GND_net), 
            .I3(n37177), .O(n8017[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_19_lut (.I0(GND_net), .I1(n8272[16]), .I2(GND_net), 
            .I3(n37377), .O(n8251[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_26 (.CI(n37177), .I0(n8047[23]), .I1(GND_net), .CO(n37178));
    SB_LUT4 i33426_3_lut (.I0(n49054), .I1(pwm_23__N_2960[19]), .I2(\PID_CONTROLLER.result [19]), 
            .I3(GND_net), .O(n48987));   // verilog/motorControl.v(44[31:51])
    defparam i33426_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3056_25_lut (.I0(GND_net), .I1(n8047[22]), .I2(GND_net), 
            .I3(n37176), .O(n8017[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_11 (.CI(n37588), .I0(n15848[8]), .I1(GND_net), .CO(n37589));
    SB_LUT4 add_3075_8_lut (.I0(GND_net), .I1(n8427[5]), .I2(n746), .I3(n37501), 
            .O(n8416[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31398_4_lut (.I0(pwm_23__N_2960[21]), .I1(n50246), .I2(\PID_CONTROLLER.result[21] ), 
            .I3(n49004), .O(n46958));
    defparam i31398_4_lut.LUT_INIT = 16'h5a7b;
    SB_CARRY add_3065_19 (.CI(n37377), .I0(n8272[16]), .I1(GND_net), .CO(n37378));
    SB_CARRY add_3056_25 (.CI(n37176), .I0(n8047[22]), .I1(GND_net), .CO(n37177));
    SB_LUT4 add_3056_24_lut (.I0(GND_net), .I1(n8047[21]), .I2(GND_net), 
            .I3(n37175), .O(n8017[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_18_lut (.I0(GND_net), .I1(n8272[15]), .I2(GND_net), 
            .I3(n37376), .O(n8251[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_24 (.CI(n37175), .I0(n8047[21]), .I1(GND_net), .CO(n37176));
    SB_LUT4 add_3056_23_lut (.I0(GND_net), .I1(n8047[20]), .I2(GND_net), 
            .I3(n37174), .O(n8017[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_7_lut (.I0(GND_net), .I1(n1798[4]), .I2(n442), 
            .I3(n37664), .O(n1797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_23 (.CI(n37174), .I0(n8047[20]), .I1(GND_net), .CO(n37175));
    SB_LUT4 add_3402_10_lut (.I0(GND_net), .I1(n15848[7]), .I2(GND_net), 
            .I3(n37587), .O(n15638[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_8 (.CI(n37501), .I0(n8427[5]), .I1(n746), .CO(n37502));
    SB_CARRY add_3065_18 (.CI(n37376), .I0(n8272[15]), .I1(GND_net), .CO(n37377));
    SB_LUT4 add_3056_22_lut (.I0(GND_net), .I1(n8047[19]), .I2(GND_net), 
            .I3(n37173), .O(n8017[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_22 (.CI(n37173), .I0(n8047[19]), .I1(GND_net), .CO(n37174));
    SB_LUT4 add_3065_17_lut (.I0(GND_net), .I1(n8272[14]), .I2(GND_net), 
            .I3(n37375), .O(n8251[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_21_lut (.I0(GND_net), .I1(n8047[18]), .I2(GND_net), 
            .I3(n37172), .O(n8017[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_21 (.CI(n37172), .I0(n8047[18]), .I1(GND_net), .CO(n37173));
    SB_CARRY add_3402_10 (.CI(n37587), .I0(n15848[7]), .I1(GND_net), .CO(n37588));
    SB_LUT4 add_3075_7_lut (.I0(GND_net), .I1(n8427[4]), .I2(n649), .I3(n37500), 
            .O(n8416[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_17 (.CI(n37375), .I0(n8272[14]), .I1(GND_net), .CO(n37376));
    SB_LUT4 add_3056_20_lut (.I0(GND_net), .I1(n8047[17]), .I2(GND_net), 
            .I3(n37171), .O(n8017[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_20 (.CI(n37171), .I0(n8047[17]), .I1(GND_net), .CO(n37172));
    SB_LUT4 add_3065_16_lut (.I0(GND_net), .I1(n8272[13]), .I2(GND_net), 
            .I3(n37374), .O(n8251[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_19_lut (.I0(GND_net), .I1(n8047[16]), .I2(GND_net), 
            .I3(n37170), .O(n8017[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_9_lut (.I0(GND_net), .I1(n1802[6]), .I2(GND_net), 
            .I3(n37758), .O(n1801[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_7 (.CI(n37664), .I0(n1798[4]), .I1(n442), 
            .CO(n37665));
    SB_LUT4 add_3402_9_lut (.I0(GND_net), .I1(n15848[6]), .I2(GND_net), 
            .I3(n37586), .O(n15638[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_7 (.CI(n37500), .I0(n8427[4]), .I1(n649), .CO(n37501));
    SB_CARRY add_3065_16 (.CI(n37374), .I0(n8272[13]), .I1(GND_net), .CO(n37375));
    SB_LUT4 add_3065_15_lut (.I0(GND_net), .I1(n8272[12]), .I2(GND_net), 
            .I3(n37373), .O(n8251[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_9 (.CI(n37586), .I0(n15848[6]), .I1(GND_net), .CO(n37587));
    SB_LUT4 add_3075_6_lut (.I0(GND_net), .I1(n8427[3]), .I2(n552), .I3(n37499), 
            .O(n8416[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_15 (.CI(n37373), .I0(n8272[12]), .I1(GND_net), .CO(n37374));
    SB_LUT4 add_3065_14_lut (.I0(GND_net), .I1(n8272[11]), .I2(GND_net), 
            .I3(n37372), .O(n8251[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_6_lut (.I0(GND_net), .I1(n1798[3]), .I2(n369), 
            .I3(n37663), .O(n1797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3402_8_lut (.I0(GND_net), .I1(n15848[5]), .I2(n728), .I3(n37585), 
            .O(n15638[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33542_4_lut (.I0(n47664), .I1(n48954), .I2(n50239), .I3(n46953), 
            .O(n49103));   // verilog/motorControl.v(44[31:51])
    defparam i33542_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3075_6 (.CI(n37499), .I0(n8427[3]), .I1(n552), .CO(n37500));
    SB_CARRY add_3065_14 (.CI(n37372), .I0(n8272[11]), .I1(GND_net), .CO(n37373));
    SB_LUT4 add_3065_13_lut (.I0(GND_net), .I1(n8272[10]), .I2(GND_net), 
            .I3(n37371), .O(n8251[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_8 (.CI(n37585), .I0(n15848[5]), .I1(n728), .CO(n37586));
    SB_LUT4 add_3075_5_lut (.I0(GND_net), .I1(n8427[2]), .I2(n455_c), 
            .I3(n37498), .O(n8416[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_13 (.CI(n37371), .I0(n8272[10]), .I1(GND_net), .CO(n37372));
    SB_LUT4 add_3065_12_lut (.I0(GND_net), .I1(n8272[9]), .I2(GND_net), 
            .I3(n37370), .O(n8251[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32111_3_lut (.I0(n48987), .I1(\pwm_23__N_2960[20] ), .I2(\PID_CONTROLLER.result[20] ), 
            .I3(GND_net), .O(n47672));   // verilog/motorControl.v(44[31:51])
    defparam i32111_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY mult_14_add_1216_9 (.CI(n37758), .I0(n1802[6]), .I1(GND_net), 
            .CO(n37759));
    SB_CARRY mult_14_add_1212_6 (.CI(n37663), .I0(n1798[3]), .I1(n369), 
            .CO(n37664));
    SB_LUT4 add_3402_7_lut (.I0(GND_net), .I1(n15848[4]), .I2(n631), .I3(n37584), 
            .O(n15638[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_5 (.CI(n37498), .I0(n8427[2]), .I1(n455_c), .CO(n37499));
    SB_CARRY add_3065_12 (.CI(n37370), .I0(n8272[9]), .I1(GND_net), .CO(n37371));
    SB_CARRY add_3056_19 (.CI(n37170), .I0(n8047[16]), .I1(GND_net), .CO(n37171));
    SB_LUT4 add_3065_11_lut (.I0(GND_net), .I1(n8272[8]), .I2(GND_net), 
            .I3(n37369), .O(n8251[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_18_lut (.I0(GND_net), .I1(n8047[15]), .I2(GND_net), 
            .I3(n37169), .O(n8017[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_18 (.CI(n37169), .I0(n8047[15]), .I1(GND_net), .CO(n37170));
    SB_LUT4 add_3075_4_lut (.I0(GND_net), .I1(n8427[1]), .I2(n358), .I3(n37497), 
            .O(n8416[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_11 (.CI(n37369), .I0(n8272[8]), .I1(GND_net), .CO(n37370));
    SB_LUT4 add_3056_17_lut (.I0(GND_net), .I1(n8047[14]), .I2(GND_net), 
            .I3(n37168), .O(n8017[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3054_29_lut (.I0(GND_net), .I1(n7986[26]), .I2(GND_net), 
            .I3(n36940), .O(n7954[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_17 (.CI(n37168), .I0(n8047[14]), .I1(GND_net), .CO(n37169));
    SB_CARRY add_3054_29 (.CI(n36940), .I0(n7986[26]), .I1(GND_net), .CO(n36941));
    SB_LUT4 add_3054_28_lut (.I0(GND_net), .I1(n7986[25]), .I2(GND_net), 
            .I3(n36939), .O(n7954[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_10_lut (.I0(GND_net), .I1(n8272[7]), .I2(GND_net), 
            .I3(n37368), .O(n8251[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_16_lut (.I0(GND_net), .I1(n8047[13]), .I2(GND_net), 
            .I3(n37167), .O(n8017[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_28 (.CI(n36939), .I0(n7986[25]), .I1(GND_net), .CO(n36940));
    SB_LUT4 add_3054_27_lut (.I0(GND_net), .I1(n7986[24]), .I2(GND_net), 
            .I3(n36938), .O(n7954[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_16 (.CI(n37167), .I0(n8047[13]), .I1(GND_net), .CO(n37168));
    SB_LUT4 i33548_4_lut (.I0(n47672), .I1(n49103), .I2(n50239), .I3(n46958), 
            .O(n49109));   // verilog/motorControl.v(44[31:51])
    defparam i33548_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3054_27 (.CI(n36938), .I0(n7986[24]), .I1(GND_net), .CO(n36939));
    SB_LUT4 add_3054_26_lut (.I0(GND_net), .I1(n7986[23]), .I2(GND_net), 
            .I3(n36937), .O(n7954[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_7 (.CI(n37584), .I0(n15848[4]), .I1(n631), .CO(n37585));
    SB_CARRY add_3075_4 (.CI(n37497), .I0(n8427[1]), .I1(n358), .CO(n37498));
    SB_CARRY add_3065_10 (.CI(n37368), .I0(n8272[7]), .I1(GND_net), .CO(n37369));
    SB_LUT4 add_3056_15_lut (.I0(GND_net), .I1(n8047[12]), .I2(GND_net), 
            .I3(n37166), .O(n8017[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_15 (.CI(n37166), .I0(n8047[12]), .I1(GND_net), .CO(n37167));
    SB_LUT4 add_3065_9_lut (.I0(GND_net), .I1(n8272[6]), .I2(GND_net), 
            .I3(n37367), .O(n8251[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_14_lut (.I0(GND_net), .I1(n8047[11]), .I2(GND_net), 
            .I3(n37165), .O(n8017[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_14 (.CI(n37165), .I0(n8047[11]), .I1(GND_net), .CO(n37166));
    SB_LUT4 add_3075_3_lut (.I0(GND_net), .I1(n8427[0]), .I2(n261), .I3(n37496), 
            .O(n8416[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_9 (.CI(n37367), .I0(n8272[6]), .I1(GND_net), .CO(n37368));
    SB_LUT4 add_3056_13_lut (.I0(GND_net), .I1(n8047[10]), .I2(GND_net), 
            .I3(n37164), .O(n8017[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_26 (.CI(n36937), .I0(n7986[23]), .I1(GND_net), .CO(n36938));
    SB_LUT4 add_3054_25_lut (.I0(GND_net), .I1(n7986[22]), .I2(GND_net), 
            .I3(n36936), .O(n7954[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_13 (.CI(n37164), .I0(n8047[10]), .I1(GND_net), .CO(n37165));
    SB_CARRY add_3054_25 (.CI(n36936), .I0(n7986[22]), .I1(GND_net), .CO(n36937));
    SB_LUT4 add_3054_24_lut (.I0(GND_net), .I1(n7986[21]), .I2(GND_net), 
            .I3(n36935), .O(n7954[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_8_lut (.I0(GND_net), .I1(n8272[5]), .I2(n716), .I3(n37366), 
            .O(n8251[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_12_lut (.I0(GND_net), .I1(n8047[9]), .I2(GND_net), 
            .I3(n37163), .O(n8017[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_24 (.CI(n36935), .I0(n7986[21]), .I1(GND_net), .CO(n36936));
    SB_LUT4 add_3054_23_lut (.I0(GND_net), .I1(n7986[20]), .I2(GND_net), 
            .I3(n36934), .O(n7954[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_12 (.CI(n37163), .I0(n8047[9]), .I1(GND_net), .CO(n37164));
    SB_CARRY add_3054_23 (.CI(n36934), .I0(n7986[20]), .I1(GND_net), .CO(n36935));
    SB_LUT4 add_3054_22_lut (.I0(GND_net), .I1(n7986[19]), .I2(GND_net), 
            .I3(n36933), .O(n7954[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_5_lut (.I0(GND_net), .I1(n1798[2]), .I2(n296), 
            .I3(n37662), .O(n1797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3402_6_lut (.I0(GND_net), .I1(n15848[3]), .I2(n534), .I3(n37583), 
            .O(n15638[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_3 (.CI(n37496), .I0(n8427[0]), .I1(n261), .CO(n37497));
    SB_LUT4 i3_4_lut (.I0(\PID_CONTROLLER.result [27]), .I1(n43891), .I2(pwm_23__N_2960[24]), 
            .I3(\PID_CONTROLLER.result [24]), .O(n8_adj_3401));   // verilog/motorControl.v(44[31:51])
    defparam i3_4_lut.LUT_INIT = 16'hdffe;
    SB_CARRY add_3065_8 (.CI(n37366), .I0(n8272[5]), .I1(n716), .CO(n37367));
    SB_LUT4 add_3056_11_lut (.I0(GND_net), .I1(n8047[8]), .I2(GND_net), 
            .I3(n37162), .O(n8017[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_11 (.CI(n37162), .I0(n8047[8]), .I1(GND_net), .CO(n37163));
    SB_LUT4 add_3065_7_lut (.I0(GND_net), .I1(n8272[4]), .I2(n619), .I3(n37365), 
            .O(n8251[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_10_lut (.I0(GND_net), .I1(n8047[7]), .I2(GND_net), 
            .I3(n37161), .O(n8017[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_10 (.CI(n37161), .I0(n8047[7]), .I1(GND_net), .CO(n37162));
    SB_LUT4 add_3075_2_lut (.I0(GND_net), .I1(n71), .I2(n164), .I3(GND_net), 
            .O(n8416[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3075_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(\PID_CONTROLLER.result [28]), .I1(n8_adj_3401), 
            .I2(\PID_CONTROLLER.result [30]), .I3(pwm_23__N_2960[24]), .O(n44147));   // verilog/motorControl.v(44[31:51])
    defparam i4_4_lut.LUT_INIT = 16'hdffe;
    SB_CARRY add_3065_7 (.CI(n37365), .I0(n8272[4]), .I1(n619), .CO(n37366));
    SB_LUT4 add_3056_9_lut (.I0(GND_net), .I1(n8047[6]), .I2(GND_net), 
            .I3(n37160), .O(n8017[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_22 (.CI(n36933), .I0(n7986[19]), .I1(GND_net), .CO(n36934));
    SB_LUT4 add_3054_21_lut (.I0(GND_net), .I1(n7986[18]), .I2(GND_net), 
            .I3(n36932), .O(n7954[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_9 (.CI(n37160), .I0(n8047[6]), .I1(GND_net), .CO(n37161));
    SB_CARRY add_3054_21 (.CI(n36932), .I0(n7986[18]), .I1(GND_net), .CO(n36933));
    SB_LUT4 add_3054_20_lut (.I0(GND_net), .I1(n7986[17]), .I2(GND_net), 
            .I3(n36931), .O(n7954[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_20 (.CI(n36931), .I0(n7986[17]), .I1(GND_net), .CO(n36932));
    SB_LUT4 add_3054_19_lut (.I0(GND_net), .I1(n7986[16]), .I2(GND_net), 
            .I3(n36930), .O(n7954[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3075_2 (.CI(GND_net), .I0(n71), .I1(n164), .CO(n37496));
    SB_LUT4 add_3065_6_lut (.I0(GND_net), .I1(n8272[3]), .I2(n522), .I3(n37364), 
            .O(n8251[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33549_3_lut (.I0(n49109), .I1(pwm_23__N_2960[23]), .I2(\PID_CONTROLLER.result [23]), 
            .I3(GND_net), .O(n49110));   // verilog/motorControl.v(44[31:51])
    defparam i33549_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3065_6 (.CI(n37364), .I0(n8272[3]), .I1(n522), .CO(n37365));
    SB_LUT4 add_3056_8_lut (.I0(GND_net), .I1(n8047[5]), .I2(n689), .I3(n37159), 
            .O(n8017[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_19 (.CI(n36930), .I0(n7986[16]), .I1(GND_net), .CO(n36931));
    SB_LUT4 add_3054_18_lut (.I0(GND_net), .I1(n7986[15]), .I2(GND_net), 
            .I3(n36929), .O(n7954[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_8 (.CI(n37159), .I0(n8047[5]), .I1(n689), .CO(n37160));
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i4_4_lut  (.I0(deadband[0]), .I1(\PID_CONTROLLER.result [1]), 
            .I2(deadband[1]), .I3(\PID_CONTROLLER.result [0]), .O(n4_adj_3402));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i4_4_lut .LUT_INIT = 16'h4d0c;
    SB_CARRY add_3054_18 (.CI(n36929), .I0(n7986[15]), .I1(GND_net), .CO(n36930));
    SB_LUT4 add_3054_17_lut (.I0(GND_net), .I1(n7986[14]), .I2(GND_net), 
            .I3(n36928), .O(n7954[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32910_3_lut (.I0(n4_adj_3402), .I1(\PID_CONTROLLER.result[13] ), 
            .I2(n27), .I3(GND_net), .O(n48471));   // verilog/motorControl.v(44[10:27])
    defparam i32910_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3402_6 (.CI(n37583), .I0(n15848[3]), .I1(n534), .CO(n37584));
    SB_LUT4 add_3074_11_lut (.I0(GND_net), .I1(n8416[8]), .I2(GND_net), 
            .I3(n37495), .O(n8404[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_5_lut (.I0(GND_net), .I1(n8272[2]), .I2(n425), .I3(n37363), 
            .O(n8251[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_7_lut (.I0(GND_net), .I1(n8047[4]), .I2(n592_adj_3404), 
            .I3(n37158), .O(n8017[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_7 (.CI(n37158), .I0(n8047[4]), .I1(n592_adj_3404), 
            .CO(n37159));
    SB_CARRY add_3065_5 (.CI(n37363), .I0(n8272[2]), .I1(n425), .CO(n37364));
    SB_LUT4 i32911_3_lut (.I0(n48471), .I1(\PID_CONTROLLER.result[14] ), 
            .I2(n29), .I3(GND_net), .O(n48472));   // verilog/motorControl.v(44[10:27])
    defparam i32911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3056_6_lut (.I0(GND_net), .I1(n8047[3]), .I2(n495), .I3(n37157), 
            .O(n8017[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_6 (.CI(n37157), .I0(n8047[3]), .I1(n495), .CO(n37158));
    SB_LUT4 add_3074_10_lut (.I0(GND_net), .I1(n8416[7]), .I2(GND_net), 
            .I3(n37494), .O(n8404[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_4_lut (.I0(GND_net), .I1(n8272[1]), .I2(n328), .I3(n37362), 
            .O(n8251[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_5_lut (.I0(GND_net), .I1(n8047[2]), .I2(n398), .I3(n37156), 
            .O(n8017[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_17 (.CI(n36928), .I0(n7986[14]), .I1(GND_net), .CO(n36929));
    SB_LUT4 add_3054_16_lut (.I0(GND_net), .I1(n7986[13]), .I2(GND_net), 
            .I3(n36927), .O(n7954[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31610_4_lut (.I0(n33), .I1(n31_adj_3406), .I2(n29), .I3(n47187), 
            .O(n47171));
    defparam i31610_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3056_5 (.CI(n37156), .I0(n8047[2]), .I1(n398), .CO(n37157));
    SB_CARRY add_3054_16 (.CI(n36927), .I0(n7986[13]), .I1(GND_net), .CO(n36928));
    SB_LUT4 add_3054_15_lut (.I0(GND_net), .I1(n7986[12]), .I2(GND_net), 
            .I3(n36926), .O(n7954[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_4 (.CI(n37362), .I0(n8272[1]), .I1(n328), .CO(n37363));
    SB_LUT4 add_3056_4_lut (.I0(GND_net), .I1(n8047[1]), .I2(n301), .I3(n37155), 
            .O(n8017[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_15 (.CI(n36926), .I0(n7986[12]), .I1(GND_net), .CO(n36927));
    SB_LUT4 add_3054_14_lut (.I0(GND_net), .I1(n7986[11]), .I2(GND_net), 
            .I3(n36925), .O(n7954[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_4 (.CI(n37155), .I0(n8047[1]), .I1(n301), .CO(n37156));
    SB_CARRY add_3054_14 (.CI(n36925), .I0(n7986[11]), .I1(GND_net), .CO(n36926));
    SB_LUT4 mult_14_add_1216_8_lut (.I0(GND_net), .I1(n1802[5]), .I2(n527), 
            .I3(n37757), .O(n1801[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_5 (.CI(n37662), .I0(n1798[2]), .I1(n296), 
            .CO(n37663));
    SB_LUT4 add_3402_5_lut (.I0(GND_net), .I1(n15848[2]), .I2(n437), .I3(n37582), 
            .O(n15638[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_10 (.CI(n37494), .I0(n8416[7]), .I1(GND_net), .CO(n37495));
    SB_LUT4 add_3065_3_lut (.I0(GND_net), .I1(n8272[0]), .I2(n231), .I3(n37361), 
            .O(n8251[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_3_lut (.I0(GND_net), .I1(n8047[0]), .I2(n204), .I3(n37154), 
            .O(n8017[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_3 (.CI(n37361), .I0(n8272[0]), .I1(n231), .CO(n37362));
    SB_LUT4 add_3074_9_lut (.I0(GND_net), .I1(n8416[6]), .I2(GND_net), 
            .I3(n37493), .O(n8404[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3065_2_lut (.I0(GND_net), .I1(n41_c), .I2(n134), .I3(GND_net), 
            .O(n8251[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3065_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3056_3 (.CI(n37154), .I0(n8047[0]), .I1(n204), .CO(n37155));
    SB_LUT4 add_3054_13_lut (.I0(GND_net), .I1(n7986[10]), .I2(GND_net), 
            .I3(n36924), .O(n7954[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3195_4_lut (.I0(GND_net), .I1(n11990[1]), .I2(n310), .I3(n36404), 
            .O(n11356[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3056_2_lut (.I0(GND_net), .I1(n14), .I2(n107_adj_3409), 
            .I3(GND_net), .O(n8017[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3056_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_4 (.CI(n36404), .I0(n11990[1]), .I1(n310), .CO(n36405));
    SB_LUT4 add_3195_3_lut (.I0(GND_net), .I1(n11990[0]), .I2(n213), .I3(n36403), 
            .O(n11356[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3195_3 (.CI(n36403), .I0(n11990[0]), .I1(n213), .CO(n36404));
    SB_LUT4 add_3195_2_lut (.I0(GND_net), .I1(n23_adj_3410), .I2(n116), 
            .I3(GND_net), .O(n11356[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3195_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3065_2 (.CI(GND_net), .I0(n41_c), .I1(n134), .CO(n37361));
    SB_CARRY add_3056_2 (.CI(GND_net), .I0(n14), .I1(n107_adj_3409), .CO(n37154));
    SB_CARRY add_3195_2 (.CI(GND_net), .I0(n23_adj_3410), .I1(n116), .CO(n36403));
    SB_LUT4 add_3359_11_lut (.I0(GND_net), .I1(n15224[8]), .I2(GND_net), 
            .I3(n36402), .O(n14910[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_30_lut (.I0(GND_net), .I1(n8017[27]), .I2(GND_net), 
            .I3(n37153), .O(n7986[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3359_10_lut (.I0(GND_net), .I1(n15224[7]), .I2(GND_net), 
            .I3(n36401), .O(n14910[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3359_10 (.CI(n36401), .I0(n15224[7]), .I1(GND_net), .CO(n36402));
    SB_LUT4 add_3359_9_lut (.I0(GND_net), .I1(n15224[6]), .I2(GND_net), 
            .I3(n36400), .O(n14910[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_2_lut (.I0(\PID_CONTROLLER.result [0]), .I1(n49815), 
            .I2(n60[0]), .I3(VCC_net), .O(n471)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 state_23__I_0_add_2_26_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n66[23]), .I3(n36153), .O(\PID_CONTROLLER.err_31__N_2825 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3359_9 (.CI(n36400), .I0(n15224[6]), .I1(GND_net), .CO(n36401));
    SB_CARRY add_3402_5 (.CI(n37582), .I0(n15848[2]), .I1(n437), .CO(n37583));
    SB_CARRY add_3074_9 (.CI(n37493), .I0(n8416[6]), .I1(GND_net), .CO(n37494));
    SB_LUT4 add_3064_21_lut (.I0(GND_net), .I1(n8251[18]), .I2(GND_net), 
            .I3(n37360), .O(n8229[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_20_lut (.I0(GND_net), .I1(n8251[17]), .I2(GND_net), 
            .I3(n37359), .O(n8229[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_8_lut (.I0(GND_net), .I1(n8416[5]), .I2(n743), .I3(n37492), 
            .O(n8404[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_20 (.CI(n37359), .I0(n8251[17]), .I1(GND_net), .CO(n37360));
    SB_LUT4 add_3055_29_lut (.I0(GND_net), .I1(n8017[26]), .I2(GND_net), 
            .I3(n37152), .O(n7986[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3359_8_lut (.I0(GND_net), .I1(n15224[5]), .I2(n545), .I3(n36399), 
            .O(n14910[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3359_8 (.CI(n36399), .I0(n15224[5]), .I1(n545), .CO(n36400));
    SB_CARRY add_3055_29 (.CI(n37152), .I0(n8017[26]), .I1(GND_net), .CO(n37153));
    SB_LUT4 add_3359_7_lut (.I0(GND_net), .I1(n15224[4]), .I2(n472), .I3(n36398), 
            .O(n14910[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n66[23]), .I3(n36152), .O(\PID_CONTROLLER.err_31__N_2825 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3359_7 (.CI(n36398), .I0(n15224[4]), .I1(n472), .CO(n36399));
    SB_LUT4 add_3359_6_lut (.I0(GND_net), .I1(n15224[3]), .I2(n399_c), 
            .I3(n36397), .O(n14910[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_25 (.CI(n36152), .I0(\motor_state[23] ), 
            .I1(n66[23]), .CO(n36153));
    SB_CARRY add_3359_6 (.CI(n36397), .I0(n15224[3]), .I1(n399_c), .CO(n36398));
    SB_LUT4 add_3064_19_lut (.I0(GND_net), .I1(n8251[16]), .I2(GND_net), 
            .I3(n37358), .O(n8229[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_28_lut (.I0(GND_net), .I1(n8017[25]), .I2(GND_net), 
            .I3(n37151), .O(n7986[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3359_5_lut (.I0(GND_net), .I1(n15224[2]), .I2(n326), .I3(n36396), 
            .O(n14910[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3359_5 (.CI(n36396), .I0(n15224[2]), .I1(n326), .CO(n36397));
    SB_CARRY add_3055_28 (.CI(n37151), .I0(n8017[25]), .I1(GND_net), .CO(n37152));
    SB_LUT4 add_3359_4_lut (.I0(GND_net), .I1(n15224[1]), .I2(n253), .I3(n36395), 
            .O(n14910[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(\motor_state[22] ), 
            .I2(n66[22]), .I3(n36151), .O(\PID_CONTROLLER.err_31__N_2825 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_2 (.CI(VCC_net), .I0(n49815), .I1(n60[0]), 
            .CO(n36035));
    SB_LUT4 unary_minus_21_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(n60[31]), 
            .I3(n36034), .O(n67[24])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n36151), .I0(\motor_state[22] ), 
            .I1(n66[22]), .CO(n36152));
    SB_CARRY add_3359_4 (.CI(n36395), .I0(n15224[1]), .I1(n253), .CO(n36396));
    SB_LUT4 add_3359_3_lut (.I0(GND_net), .I1(n15224[0]), .I2(n180), .I3(n36394), 
            .O(n14910[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(\motor_state[21] ), 
            .I2(n66[21]), .I3(n36150), .O(\PID_CONTROLLER.err_31__N_2825 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n60[31]), 
            .I3(n36033), .O(n67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_25 (.CI(n36033), .I0(GND_net), .I1(n60[31]), 
            .CO(n36034));
    SB_CARRY state_23__I_0_add_2_23 (.CI(n36150), .I0(\motor_state[21] ), 
            .I1(n66[21]), .CO(n36151));
    SB_CARRY add_3359_3 (.CI(n36394), .I0(n15224[0]), .I1(n180), .CO(n36395));
    SB_LUT4 mult_14_add_1212_4_lut (.I0(GND_net), .I1(n1798[1]), .I2(n223), 
            .I3(n37661), .O(n1797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3402_4_lut (.I0(GND_net), .I1(n15848[1]), .I2(n340), .I3(n37581), 
            .O(n15638[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_8 (.CI(n37492), .I0(n8416[5]), .I1(n743), .CO(n37493));
    SB_CARRY add_3064_19 (.CI(n37358), .I0(n8251[16]), .I1(GND_net), .CO(n37359));
    SB_LUT4 add_3064_18_lut (.I0(GND_net), .I1(n8251[15]), .I2(GND_net), 
            .I3(n37357), .O(n8229[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33316_4_lut (.I0(n30_adj_3414), .I1(n10_adj_3415), .I2(n35_adj_3416), 
            .I3(n47167), .O(n48877));   // verilog/motorControl.v(44[10:27])
    defparam i33316_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3064_18 (.CI(n37357), .I0(n8251[15]), .I1(GND_net), .CO(n37358));
    SB_CARRY mult_14_add_1216_8 (.CI(n37757), .I0(n1802[5]), .I1(n527), 
            .CO(n37758));
    SB_CARRY add_3402_4 (.CI(n37581), .I0(n15848[1]), .I1(n340), .CO(n37582));
    SB_LUT4 add_3074_7_lut (.I0(GND_net), .I1(n8416[4]), .I2(n646), .I3(n37491), 
            .O(n8404[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_7 (.CI(n37491), .I0(n8416[4]), .I1(n646), .CO(n37492));
    SB_LUT4 add_3064_17_lut (.I0(GND_net), .I1(n8251[14]), .I2(GND_net), 
            .I3(n37356), .O(n8229[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_27_lut (.I0(GND_net), .I1(n8017[24]), .I2(GND_net), 
            .I3(n37150), .O(n7986[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_17 (.CI(n37356), .I0(n8251[14]), .I1(GND_net), .CO(n37357));
    SB_CARRY add_3055_27 (.CI(n37150), .I0(n8017[24]), .I1(GND_net), .CO(n37151));
    SB_CARRY mult_14_add_1212_4 (.CI(n37661), .I0(n1798[1]), .I1(n223), 
            .CO(n37662));
    SB_LUT4 add_3055_26_lut (.I0(GND_net), .I1(n8017[23]), .I2(GND_net), 
            .I3(n37149), .O(n7986[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3359_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n14910[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3359_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3359_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n36394));
    SB_CARRY add_3055_26 (.CI(n37149), .I0(n8017[23]), .I1(GND_net), .CO(n37150));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(\motor_state[20] ), 
            .I2(n66[20]), .I3(n36149), .O(\PID_CONTROLLER.err_31__N_2825 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32089_3_lut (.I0(n48472), .I1(\PID_CONTROLLER.result [15]), 
            .I2(n31_adj_3406), .I3(GND_net), .O(n47650));   // verilog/motorControl.v(44[10:27])
    defparam i32089_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n36149), .I0(\motor_state[20] ), 
            .I1(n66[20]), .CO(n36150));
    SB_LUT4 add_3064_16_lut (.I0(GND_net), .I1(n8251[13]), .I2(GND_net), 
            .I3(n37355), .O(n8229[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_25_lut (.I0(GND_net), .I1(n8017[22]), .I2(GND_net), 
            .I3(n37148), .O(n7986[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33490_4_lut (.I0(n47650), .I1(n48877), .I2(n35_adj_3416), 
            .I3(n47171), .O(n49051));   // verilog/motorControl.v(44[10:27])
    defparam i33490_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3055_25 (.CI(n37148), .I0(n8017[22]), .I1(GND_net), .CO(n37149));
    SB_LUT4 i33491_3_lut (.I0(n49051), .I1(\PID_CONTROLLER.result [18]), 
            .I2(n37), .I3(GND_net), .O(n49052));   // verilog/motorControl.v(44[10:27])
    defparam i33491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(\motor_state[19] ), 
            .I2(n66[19]), .I3(n36148), .O(\PID_CONTROLLER.err_31__N_2825 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n60[22]), 
            .I3(n36032), .O(n67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n36148), .I0(\motor_state[19] ), 
            .I1(n66[19]), .CO(n36149));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(\motor_state[18] ), 
            .I2(n66[18]), .I3(n36147), .O(\PID_CONTROLLER.err_31__N_2825 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_24 (.CI(n36032), .I0(GND_net), .I1(n60[22]), 
            .CO(n36033));
    SB_CARRY state_23__I_0_add_2_20 (.CI(n36147), .I0(\motor_state[18] ), 
            .I1(n66[18]), .CO(n36148));
    SB_LUT4 add_3402_3_lut (.I0(GND_net), .I1(n15848[0]), .I2(n243), .I3(n37580), 
            .O(n15638[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_6_lut (.I0(GND_net), .I1(n8416[3]), .I2(n549), .I3(n37490), 
            .O(n8404[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_16 (.CI(n37355), .I0(n8251[13]), .I1(GND_net), .CO(n37356));
    SB_LUT4 add_3064_15_lut (.I0(GND_net), .I1(n8251[12]), .I2(GND_net), 
            .I3(n37354), .O(n8229[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_6 (.CI(n37490), .I0(n8416[3]), .I1(n549), .CO(n37491));
    SB_CARRY add_3064_15 (.CI(n37354), .I0(n8251[12]), .I1(GND_net), .CO(n37355));
    SB_LUT4 add_3055_24_lut (.I0(GND_net), .I1(n8017[21]), .I2(GND_net), 
            .I3(n37147), .O(n7986[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_24 (.CI(n37147), .I0(n8017[21]), .I1(GND_net), .CO(n37148));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(\motor_state[17] ), 
            .I2(n66[17]), .I3(n36146), .O(\PID_CONTROLLER.err_31__N_2825 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_25_lut (.I0(GND_net), .I1(n12573[22]), .I2(GND_net), 
            .I3(n36387), .O(n11990[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_24_lut (.I0(GND_net), .I1(n12573[21]), .I2(GND_net), 
            .I3(n36386), .O(n11990[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n36146), .I0(\motor_state[17] ), 
            .I1(n66[17]), .CO(n36147));
    SB_CARRY add_3221_24 (.CI(n36386), .I0(n12573[21]), .I1(GND_net), 
            .CO(n36387));
    SB_LUT4 add_3064_14_lut (.I0(GND_net), .I1(n8251[11]), .I2(GND_net), 
            .I3(n37353), .O(n8229[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_23_lut (.I0(GND_net), .I1(n8017[20]), .I2(GND_net), 
            .I3(n37146), .O(n7986[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_23_lut (.I0(GND_net), .I1(n12573[20]), .I2(GND_net), 
            .I3(n36385), .O(n11990[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_23 (.CI(n36385), .I0(n12573[20]), .I1(GND_net), 
            .CO(n36386));
    SB_CARRY add_3055_23 (.CI(n37146), .I0(n8017[20]), .I1(GND_net), .CO(n37147));
    SB_LUT4 add_3221_22_lut (.I0(GND_net), .I1(n12573[19]), .I2(GND_net), 
            .I3(n36384), .O(n11990[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_22 (.CI(n36384), .I0(n12573[19]), .I1(GND_net), 
            .CO(n36385));
    SB_LUT4 i33430_3_lut (.I0(n49052), .I1(\PID_CONTROLLER.result [19]), 
            .I2(n39), .I3(GND_net), .O(n48991));   // verilog/motorControl.v(44[10:27])
    defparam i33430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33562_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [29]), 
            .I2(\PID_CONTROLLER.result [30]), .I3(n49081), .O(n49123));
    defparam i33562_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33358_4_lut (.I0(n47660), .I1(n48917), .I2(n50234), .I3(n48592), 
            .O(n48919));   // verilog/motorControl.v(44[10:27])
    defparam i33358_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32095_3_lut (.I0(n48991), .I1(\PID_CONTROLLER.result[20] ), 
            .I2(n41), .I3(GND_net), .O(n47656));   // verilog/motorControl.v(44[10:27])
    defparam i32095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33511_4_lut (.I0(n49110), .I1(\PID_CONTROLLER.result [31]), 
            .I2(pwm_23__N_2960[24]), .I3(n44147), .O(pwm_23__N_2959));   // verilog/motorControl.v(44[31:51])
    defparam i33511_4_lut.LUT_INIT = 16'hcc8e;
    SB_LUT4 i33360_3_lut (.I0(n47656), .I1(n48919), .I2(n49123), .I3(GND_net), 
            .O(n48921));   // verilog/motorControl.v(44[10:27])
    defparam i33360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_23__I_818_4_lut (.I0(n48921), .I1(pwm_23__N_2959), .I2(deadband[23]), 
            .I3(\PID_CONTROLLER.result [31]), .O(pwm_23__N_2957));   // verilog/motorControl.v(44[10:51])
    defparam pwm_23__I_818_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(\motor_state[16] ), 
            .I2(n66[16]), .I3(n36145), .O(\PID_CONTROLLER.err_31__N_2825 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n60[21]), 
            .I3(n36031), .O(n399)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_23 (.CI(n36031), .I0(GND_net), .I1(n60[21]), 
            .CO(n36032));
    SB_CARRY state_23__I_0_add_2_18 (.CI(n36145), .I0(\motor_state[16] ), 
            .I1(n66[16]), .CO(n36146));
    SB_LUT4 add_3074_5_lut (.I0(GND_net), .I1(n8416[2]), .I2(n452_c), 
            .I3(n37489), .O(n8404[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3402_3 (.CI(n37580), .I0(n15848[0]), .I1(n243), .CO(n37581));
    SB_DFF pwm__i23 (.Q(pwm[23]), .C(clk32MHz), .D(n24225));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i22 (.Q(pwm[22]), .C(clk32MHz), .D(n24224));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i21 (.Q(pwm[21]), .C(clk32MHz), .D(n24223));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i20 (.Q(pwm[20]), .C(clk32MHz), .D(n24222));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i19 (.Q(pwm[19]), .C(clk32MHz), .D(n24221));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i18 (.Q(pwm[18]), .C(clk32MHz), .D(n24220));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i17 (.Q(pwm[17]), .C(clk32MHz), .D(n24219));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i16 (.Q(pwm[16]), .C(clk32MHz), .D(n24218));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i15 (.Q(pwm[15]), .C(clk32MHz), .D(n24217));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i14 (.Q(pwm[14]), .C(clk32MHz), .D(n24216));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i13 (.Q(pwm[13]), .C(clk32MHz), .D(n24215));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i12 (.Q(pwm[12]), .C(clk32MHz), .D(n24214));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i11 (.Q(pwm[11]), .C(clk32MHz), .D(n24213));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i10 (.Q(pwm[10]), .C(clk32MHz), .D(n24212));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i9 (.Q(pwm[9]), .C(clk32MHz), .D(n24211));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i8 (.Q(pwm[8]), .C(clk32MHz), .D(n24210));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i7 (.Q(pwm[7]), .C(clk32MHz), .D(n24209));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i6 (.Q(pwm[6]), .C(clk32MHz), .D(n24208));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i5 (.Q(pwm[5]), .C(clk32MHz), .D(n24207));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i4 (.Q(pwm[4]), .C(clk32MHz), .D(n24206));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3055_22_lut (.I0(GND_net), .I1(n8017[19]), .I2(GND_net), 
            .I3(n37145), .O(n7986[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_22_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm__i3 (.Q(pwm[3]), .C(clk32MHz), .D(n24205));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i2 (.Q(pwm[2]), .C(clk32MHz), .D(n24204));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i1 (.Q(pwm[1]), .C(clk32MHz), .D(n24203));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF pwm__i0 (.Q(pwm[0]), .C(clk32MHz), .D(n24172));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_14_add_1216_7_lut (.I0(GND_net), .I1(n1802[4]), .I2(n454_c), 
            .I3(n37756), .O(n1801[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_3_lut (.I0(GND_net), .I1(n1798[0]), .I2(n150), 
            .I3(n37660), .O(n1797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n60[20]), 
            .I3(n36030), .O(n400)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_13 (.CI(n36924), .I0(n7986[10]), .I1(GND_net), .CO(n36925));
    SB_CARRY mult_14_add_1216_7 (.CI(n37756), .I0(n1802[4]), .I1(n454_c), 
            .CO(n37757));
    SB_CARRY add_13_add_1_21902_add_1_28 (.CI(n35912), .I0(n7063[3]), .I1(n58[26]), 
            .CO(n35913));
    SB_CARRY add_3064_14 (.CI(n37353), .I0(n8251[11]), .I1(GND_net), .CO(n37354));
    SB_CARRY add_3055_22 (.CI(n37145), .I0(n8017[19]), .I1(GND_net), .CO(n37146));
    SB_LUT4 add_3064_13_lut (.I0(GND_net), .I1(n8251[10]), .I2(GND_net), 
            .I3(n37352), .O(n8229[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_6_lut (.I0(GND_net), .I1(n1802[3]), .I2(n381), 
            .I3(n37755), .O(n1801[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3054_12_lut (.I0(GND_net), .I1(n7986[9]), .I2(GND_net), 
            .I3(n36923), .O(n7954[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_21_lut (.I0(GND_net), .I1(n8017[18]), .I2(GND_net), 
            .I3(n37144), .O(n7986[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_21 (.CI(n37144), .I0(n8017[18]), .I1(GND_net), .CO(n37145));
    SB_CARRY mult_14_add_1216_6 (.CI(n37755), .I0(n1802[3]), .I1(n381), 
            .CO(n37756));
    SB_LUT4 mult_14_add_1216_5_lut (.I0(GND_net), .I1(n1802[2]), .I2(n308), 
            .I3(n37754), .O(n1801[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_5 (.CI(n37754), .I0(n1802[2]), .I1(n308), 
            .CO(n37755));
    SB_LUT4 add_3055_20_lut (.I0(GND_net), .I1(n8017[17]), .I2(GND_net), 
            .I3(n37143), .O(n7986[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_12 (.CI(n36923), .I0(n7986[9]), .I1(GND_net), .CO(n36924));
    SB_LUT4 add_3221_21_lut (.I0(GND_net), .I1(n12573[18]), .I2(GND_net), 
            .I3(n36383), .O(n11990[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_20 (.CI(n37143), .I0(n8017[17]), .I1(GND_net), .CO(n37144));
    SB_CARRY add_3064_13 (.CI(n37352), .I0(n8251[10]), .I1(GND_net), .CO(n37353));
    SB_LUT4 add_13_add_1_21902_add_1_27_lut (.I0(GND_net), .I1(n7063[2]), 
            .I2(n58[25]), .I3(n35911), .O(n57[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_19_lut (.I0(GND_net), .I1(n8017[16]), .I2(GND_net), 
            .I3(n37142), .O(n7986[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_22 (.CI(n36030), .I0(GND_net), .I1(n60[20]), 
            .CO(n36031));
    SB_LUT4 add_3054_11_lut (.I0(GND_net), .I1(n7986[8]), .I2(GND_net), 
            .I3(n36922), .O(n7954[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_11 (.CI(n36922), .I0(n7986[8]), .I1(GND_net), .CO(n36923));
    SB_CARRY add_3055_19 (.CI(n37142), .I0(n8017[16]), .I1(GND_net), .CO(n37143));
    SB_LUT4 add_3054_10_lut (.I0(GND_net), .I1(n7986[7]), .I2(GND_net), 
            .I3(n36921), .O(n7954[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_10 (.CI(n36921), .I0(n7986[7]), .I1(GND_net), .CO(n36922));
    SB_LUT4 add_3402_2_lut (.I0(GND_net), .I1(n53_adj_3424), .I2(n146), 
            .I3(GND_net), .O(n15638[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3402_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3074_5 (.CI(n37489), .I0(n8416[2]), .I1(n452_c), .CO(n37490));
    SB_LUT4 add_3064_12_lut (.I0(GND_net), .I1(n8251[9]), .I2(GND_net), 
            .I3(n37351), .O(n8229[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_18_lut (.I0(GND_net), .I1(n8017[15]), .I2(GND_net), 
            .I3(n37141), .O(n7986[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_18 (.CI(n37141), .I0(n8017[15]), .I1(GND_net), .CO(n37142));
    SB_CARRY add_3064_12 (.CI(n37351), .I0(n8251[9]), .I1(GND_net), .CO(n37352));
    SB_LUT4 add_3055_17_lut (.I0(GND_net), .I1(n8017[14]), .I2(GND_net), 
            .I3(n37140), .O(n7986[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3054_9_lut (.I0(GND_net), .I1(n7986[6]), .I2(GND_net), 
            .I3(n36920), .O(n7954[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_9 (.CI(n36920), .I0(n7986[6]), .I1(GND_net), .CO(n36921));
    SB_CARRY add_3055_17 (.CI(n37140), .I0(n8017[14]), .I1(GND_net), .CO(n37141));
    SB_LUT4 add_3054_8_lut (.I0(GND_net), .I1(n7986[5]), .I2(n683), .I3(n36919), 
            .O(n7954[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_8 (.CI(n36919), .I0(n7986[5]), .I1(n683), .CO(n36920));
    SB_LUT4 add_3074_4_lut (.I0(GND_net), .I1(n8416[1]), .I2(n355), .I3(n37488), 
            .O(n8404[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_11_lut (.I0(GND_net), .I1(n8251[8]), .I2(GND_net), 
            .I3(n37350), .O(n8229[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_16_lut (.I0(GND_net), .I1(n8017[13]), .I2(GND_net), 
            .I3(n37139), .O(n7986[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_16 (.CI(n37139), .I0(n8017[13]), .I1(GND_net), .CO(n37140));
    SB_CARRY add_3064_11 (.CI(n37350), .I0(n8251[8]), .I1(GND_net), .CO(n37351));
    SB_LUT4 add_3055_15_lut (.I0(GND_net), .I1(n8017[12]), .I2(GND_net), 
            .I3(n37138), .O(n7986[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3054_7_lut (.I0(GND_net), .I1(n7986[4]), .I2(n586), .I3(n36918), 
            .O(n7954[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_7 (.CI(n36918), .I0(n7986[4]), .I1(n586), .CO(n36919));
    SB_CARRY add_3055_15 (.CI(n37138), .I0(n8017[12]), .I1(GND_net), .CO(n37139));
    SB_LUT4 add_3054_6_lut (.I0(GND_net), .I1(n7986[3]), .I2(n489), .I3(n36917), 
            .O(n7954[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_4_lut (.I0(GND_net), .I1(n1802[1]), .I2(n235), 
            .I3(n37753), .O(n1801[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_10_lut (.I0(GND_net), .I1(n8251[7]), .I2(GND_net), 
            .I3(n37349), .O(n8229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_3 (.CI(n37660), .I0(n1798[0]), .I1(n150), 
            .CO(n37661));
    SB_CARRY add_13_add_1_21902_add_1_27 (.CI(n35911), .I0(n7063[2]), .I1(n58[25]), 
            .CO(n35912));
    SB_CARRY add_3402_2 (.CI(GND_net), .I0(n53_adj_3424), .I1(n146), .CO(n37580));
    SB_CARRY add_3074_4 (.CI(n37488), .I0(n8416[1]), .I1(n355), .CO(n37489));
    SB_CARRY add_3054_6 (.CI(n36917), .I0(n7986[3]), .I1(n489), .CO(n36918));
    SB_CARRY add_3064_10 (.CI(n37349), .I0(n8251[7]), .I1(GND_net), .CO(n37350));
    SB_LUT4 add_3055_14_lut (.I0(GND_net), .I1(n8017[11]), .I2(GND_net), 
            .I3(n37137), .O(n7986[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_9_lut (.I0(GND_net), .I1(n8251[6]), .I2(GND_net), 
            .I3(n37348), .O(n8229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_14 (.CI(n37137), .I0(n8017[11]), .I1(GND_net), .CO(n37138));
    SB_CARRY add_3064_9 (.CI(n37348), .I0(n8251[6]), .I1(GND_net), .CO(n37349));
    SB_LUT4 add_3054_5_lut (.I0(GND_net), .I1(n7986[2]), .I2(n392), .I3(n36916), 
            .O(n7954[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(\motor_state[15] ), 
            .I2(n66[15]), .I3(n36144), .O(\PID_CONTROLLER.err_31__N_2825 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_3_lut (.I0(GND_net), .I1(n8416[0]), .I2(n258), .I3(n37487), 
            .O(n8404[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_21 (.CI(n36383), .I0(n12573[18]), .I1(GND_net), 
            .CO(n36384));
    SB_DFF \PID_CONTROLLER.result_i0  (.Q(\PID_CONTROLLER.result [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [0]));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY state_23__I_0_add_2_17 (.CI(n36144), .I0(\motor_state[15] ), 
            .I1(n66[15]), .CO(n36145));
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err[0] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [0]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF GATES_i2 (.Q(PIN_7_c_1), .C(clk32MHz), .D(GATES_5__N_2788[1]));   // verilog/motorControl.v(64[10] 111[6])
    SB_LUT4 add_3055_13_lut (.I0(GND_net), .I1(n8017[10]), .I2(GND_net), 
            .I3(n37136), .O(n7986[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n60[19]), 
            .I3(n36029), .O(n67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(\motor_state[14] ), 
            .I2(n66[14]), .I3(n36143), .O(\PID_CONTROLLER.err_31__N_2825 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_20_lut (.I0(GND_net), .I1(n12573[17]), .I2(GND_net), 
            .I3(n36382), .O(n11990[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_20 (.CI(n36382), .I0(n12573[17]), .I1(GND_net), 
            .CO(n36383));
    SB_LUT4 add_3221_19_lut (.I0(GND_net), .I1(n12573[16]), .I2(GND_net), 
            .I3(n36381), .O(n11990[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n36143), .I0(\motor_state[14] ), 
            .I1(n66[14]), .CO(n36144));
    SB_CARRY add_3221_19 (.CI(n36381), .I0(n12573[16]), .I1(GND_net), 
            .CO(n36382));
    SB_CARRY add_3074_3 (.CI(n37487), .I0(n8416[0]), .I1(n258), .CO(n37488));
    SB_LUT4 add_3064_8_lut (.I0(GND_net), .I1(n8251[5]), .I2(n713), .I3(n37347), 
            .O(n8229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_8 (.CI(n37347), .I0(n8251[5]), .I1(n713), .CO(n37348));
    SB_CARRY add_3055_13 (.CI(n37136), .I0(n8017[10]), .I1(GND_net), .CO(n37137));
    SB_LUT4 add_3221_18_lut (.I0(GND_net), .I1(n12573[15]), .I2(GND_net), 
            .I3(n36380), .O(n11990[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_18 (.CI(n36380), .I0(n12573[15]), .I1(GND_net), 
            .CO(n36381));
    SB_LUT4 add_3055_12_lut (.I0(GND_net), .I1(n8017[9]), .I2(GND_net), 
            .I3(n37135), .O(n7986[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_17_lut (.I0(GND_net), .I1(n12573[14]), .I2(GND_net), 
            .I3(n36379), .O(n11990[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_4 (.CI(n37753), .I0(n1802[1]), .I1(n235), 
            .CO(n37754));
    SB_DFF GATES_i1 (.Q(PIN_6_c_0), .C(clk32MHz), .D(GATES_5__N_2788[0]));   // verilog/motorControl.v(64[10] 111[6])
    SB_CARRY unary_minus_21_add_3_21 (.CI(n36029), .I0(GND_net), .I1(n60[19]), 
            .CO(n36030));
    SB_CARRY add_3221_17 (.CI(n36379), .I0(n12573[14]), .I1(GND_net), 
            .CO(n36380));
    SB_LUT4 add_3064_7_lut (.I0(GND_net), .I1(n8251[4]), .I2(n616), .I3(n37346), 
            .O(n8229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(\motor_state[13] ), 
            .I2(n66[13]), .I3(n36142), .O(\PID_CONTROLLER.err_31__N_2825 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n36142), .I0(\motor_state[13] ), 
            .I1(n66[13]), .CO(n36143));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(\motor_state[12] ), 
            .I2(n66[12]), .I3(n36141), .O(\PID_CONTROLLER.err_31__N_2825 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_12 (.CI(n37135), .I0(n8017[9]), .I1(GND_net), .CO(n37136));
    SB_CARRY add_3054_5 (.CI(n36916), .I0(n7986[2]), .I1(n392), .CO(n36917));
    SB_LUT4 add_3486_8_lut (.I0(GND_net), .I1(n16627[5]), .I2(n752_adj_3431), 
            .I3(n37579), .O(n16618[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3486_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_16_lut (.I0(GND_net), .I1(n12573[13]), .I2(GND_net), 
            .I3(n36378), .O(n11990[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3054_4_lut (.I0(GND_net), .I1(n7986[1]), .I2(n295), .I3(n36915), 
            .O(n7954[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_16 (.CI(n36378), .I0(n12573[13]), .I1(GND_net), 
            .CO(n36379));
    SB_LUT4 add_3055_11_lut (.I0(GND_net), .I1(n8017[8]), .I2(GND_net), 
            .I3(n37134), .O(n7986[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_4 (.CI(n36915), .I0(n7986[1]), .I1(n295), .CO(n36916));
    SB_LUT4 add_3054_3_lut (.I0(GND_net), .I1(n7986[0]), .I2(n198), .I3(n36914), 
            .O(n7954[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_3 (.CI(n36914), .I0(n7986[0]), .I1(n198), .CO(n36915));
    SB_CARRY state_23__I_0_add_2_14 (.CI(n36141), .I0(\motor_state[12] ), 
            .I1(n66[12]), .CO(n36142));
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(\motor_state[11] ), 
            .I2(n66[11]), .I3(n36140), .O(\PID_CONTROLLER.err_31__N_2825 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n60[18]), 
            .I3(n36028), .O(n67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n36140), .I0(\motor_state[11] ), 
            .I1(n66[11]), .CO(n36141));
    SB_LUT4 add_3054_2_lut (.I0(GND_net), .I1(n8_adj_3433), .I2(n101), 
            .I3(GND_net), .O(n7954[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3054_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_15_lut (.I0(GND_net), .I1(n12573[12]), .I2(GND_net), 
            .I3(n36377), .O(n11990[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3486_7_lut (.I0(GND_net), .I1(n16627[4]), .I2(n658), .I3(n37578), 
            .O(n16618[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3486_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3074_2_lut (.I0(GND_net), .I1(n68), .I2(n161), .I3(GND_net), 
            .O(n8404[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3074_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_7 (.CI(n37346), .I0(n8251[4]), .I1(n616), .CO(n37347));
    SB_LUT4 add_3064_6_lut (.I0(GND_net), .I1(n8251[3]), .I2(n519_adj_3434), 
            .I3(n37345), .O(n8229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_11 (.CI(n37134), .I0(n8017[8]), .I1(GND_net), .CO(n37135));
    SB_CARRY add_3221_15 (.CI(n36377), .I0(n12573[12]), .I1(GND_net), 
            .CO(n36378));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(\motor_state[10] ), 
            .I2(n66[10]), .I3(n36139), .O(\PID_CONTROLLER.err_31__N_2825 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_14_lut (.I0(GND_net), .I1(n12573[11]), .I2(GND_net), 
            .I3(n36376), .O(n11990[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_10_lut (.I0(GND_net), .I1(n8017[7]), .I2(GND_net), 
            .I3(n37133), .O(n7986[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_3_lut (.I0(GND_net), .I1(n1802[0]), .I2(n162), 
            .I3(n37752), .O(n1801[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_14 (.CI(n36376), .I0(n12573[11]), .I1(GND_net), 
            .CO(n36377));
    SB_CARRY state_23__I_0_add_2_12 (.CI(n36139), .I0(\motor_state[10] ), 
            .I1(n66[10]), .CO(n36140));
    SB_LUT4 add_3221_13_lut (.I0(GND_net), .I1(n12573[10]), .I2(GND_net), 
            .I3(n36375), .O(n11990[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_13 (.CI(n36375), .I0(n12573[10]), .I1(GND_net), 
            .CO(n36376));
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(\motor_state[9] ), 
            .I2(n66[9]), .I3(n36138), .O(\PID_CONTROLLER.err_31__N_2825 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_12_lut (.I0(GND_net), .I1(n12573[9]), .I2(GND_net), 
            .I3(n36374), .O(n11990[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_3 (.CI(n37752), .I0(n1802[0]), .I1(n162), 
            .CO(n37753));
    SB_CARRY add_3074_2 (.CI(GND_net), .I0(n68), .I1(n161), .CO(n37487));
    SB_CARRY add_3064_6 (.CI(n37345), .I0(n8251[3]), .I1(n519_adj_3434), 
            .CO(n37346));
    SB_LUT4 add_3064_5_lut (.I0(GND_net), .I1(n8251[2]), .I2(n422), .I3(n37344), 
            .O(n8229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_10 (.CI(n37133), .I0(n8017[7]), .I1(GND_net), .CO(n37134));
    SB_CARRY add_3221_12 (.CI(n36374), .I0(n12573[9]), .I1(GND_net), .CO(n36375));
    SB_LUT4 add_3221_11_lut (.I0(GND_net), .I1(n12573[8]), .I2(GND_net), 
            .I3(n36373), .O(n11990[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_9_lut (.I0(GND_net), .I1(n8017[6]), .I2(GND_net), 
            .I3(n37132), .O(n7986[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_11 (.CI(n36373), .I0(n12573[8]), .I1(GND_net), .CO(n36374));
    SB_CARRY state_23__I_0_add_2_11 (.CI(n36138), .I0(\motor_state[9] ), 
            .I1(n66[9]), .CO(n36139));
    SB_CARRY unary_minus_21_add_3_20 (.CI(n36028), .I0(GND_net), .I1(n60[18]), 
            .CO(n36029));
    SB_LUT4 unary_minus_21_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n60[17]), 
            .I3(n36027), .O(n67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(\motor_state[8] ), 
            .I2(n66[8]), .I3(n36137), .O(\PID_CONTROLLER.err_31__N_2825 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_10_lut (.I0(GND_net), .I1(n12573[7]), .I2(GND_net), 
            .I3(n36372), .O(n11990[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_10 (.CI(n36372), .I0(n12573[7]), .I1(GND_net), .CO(n36373));
    SB_LUT4 mult_14_add_1216_2_lut (.I0(GND_net), .I1(n20_adj_3439), .I2(n89), 
            .I3(GND_net), .O(n1801[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n36137), .I0(\motor_state[8] ), 
            .I1(n66[8]), .CO(n36138));
    SB_CARRY unary_minus_21_add_3_19 (.CI(n36027), .I0(GND_net), .I1(n60[17]), 
            .CO(n36028));
    SB_LUT4 unary_minus_21_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n60[16]), 
            .I3(n36026), .O(n67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(\motor_state[7] ), 
            .I2(n66[7]), .I3(n36136), .O(\PID_CONTROLLER.err_31__N_2825 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_9_lut (.I0(GND_net), .I1(n12573[6]), .I2(GND_net), 
            .I3(n36371), .O(n11990[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_2_lut (.I0(GND_net), .I1(n8_adj_3443), .I2(n77), 
            .I3(GND_net), .O(n1797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3486_7 (.CI(n37578), .I0(n16627[4]), .I1(n658), .CO(n37579));
    SB_LUT4 add_3073_12_lut (.I0(GND_net), .I1(n8404[9]), .I2(GND_net), 
            .I3(n37486), .O(n8391[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_5 (.CI(n37344), .I0(n8251[2]), .I1(n422), .CO(n37345));
    SB_LUT4 add_3064_4_lut (.I0(GND_net), .I1(n8251[1]), .I2(n325), .I3(n37343), 
            .O(n8229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_9 (.CI(n37132), .I0(n8017[6]), .I1(GND_net), .CO(n37133));
    SB_CARRY mult_14_add_1212_2 (.CI(GND_net), .I0(n8_adj_3443), .I1(n77), 
            .CO(n37660));
    SB_CARRY add_3221_9 (.CI(n36371), .I0(n12573[6]), .I1(GND_net), .CO(n36372));
    SB_LUT4 add_3486_6_lut (.I0(GND_net), .I1(n16627[3]), .I2(n558), .I3(n37577), 
            .O(n16618[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3486_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_8_lut (.I0(GND_net), .I1(n12573[5]), .I2(n701), .I3(n36370), 
            .O(n11990[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_8_lut (.I0(GND_net), .I1(n8017[5]), .I2(n686), .I3(n37131), 
            .O(n7986[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_8 (.CI(n36370), .I0(n12573[5]), .I1(n701), .CO(n36371));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n36136), .I0(\motor_state[7] ), 
            .I1(n66[7]), .CO(n36137));
    SB_LUT4 add_3221_7_lut (.I0(GND_net), .I1(n12573[4]), .I2(n604_adj_3444), 
            .I3(n36369), .O(n11990[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_7 (.CI(n36369), .I0(n12573[4]), .I1(n604_adj_3444), 
            .CO(n36370));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(\motor_state[6] ), 
            .I2(n66[6]), .I3(n36135), .O(\PID_CONTROLLER.err_31__N_2825 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3221_6_lut (.I0(GND_net), .I1(n12573[3]), .I2(n507), .I3(n36368), 
            .O(n11990[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_11_lut (.I0(GND_net), .I1(n8404[8]), .I2(GND_net), 
            .I3(n37485), .O(n8391[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_4 (.CI(n37343), .I0(n8251[1]), .I1(n325), .CO(n37344));
    SB_LUT4 add_3064_3_lut (.I0(GND_net), .I1(n8251[0]), .I2(n228), .I3(n37342), 
            .O(n8229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_8 (.CI(n37131), .I0(n8017[5]), .I1(n686), .CO(n37132));
    SB_CARRY add_3221_6 (.CI(n36368), .I0(n12573[3]), .I1(n507), .CO(n36369));
    SB_LUT4 add_3221_5_lut (.I0(GND_net), .I1(n12573[2]), .I2(n410), .I3(n36367), 
            .O(n11990[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_11 (.CI(n37485), .I0(n8404[8]), .I1(GND_net), .CO(n37486));
    SB_LUT4 add_3055_7_lut (.I0(GND_net), .I1(n8017[4]), .I2(n589_adj_3446), 
            .I3(n37130), .O(n7986[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n36135), .I0(\motor_state[6] ), 
            .I1(n66[6]), .CO(n36136));
    SB_CARRY add_3221_5 (.CI(n36367), .I0(n12573[2]), .I1(n410), .CO(n36368));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(\motor_state[5] ), 
            .I2(n66[5]), .I3(n36134), .O(\PID_CONTROLLER.err_31__N_2825 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3064_3 (.CI(n37342), .I0(n8251[0]), .I1(n228), .CO(n37343));
    SB_CARRY unary_minus_21_add_3_18 (.CI(n36026), .I0(GND_net), .I1(n60[16]), 
            .CO(n36027));
    SB_CARRY state_23__I_0_add_2_7 (.CI(n36134), .I0(\motor_state[5] ), 
            .I1(n66[5]), .CO(n36135));
    SB_LUT4 add_3221_4_lut (.I0(GND_net), .I1(n12573[1]), .I2(n313), .I3(n36366), 
            .O(n11990[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_4 (.CI(n36366), .I0(n12573[1]), .I1(n313), .CO(n36367));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(\motor_state[4] ), 
            .I2(n66[4]), .I3(n36133), .O(\PID_CONTROLLER.err_31__N_2825 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n60[15]), 
            .I3(n36025), .O(n67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n36133), .I0(\motor_state[4] ), 
            .I1(n66[4]), .CO(n36134));
    SB_CARRY add_3055_7 (.CI(n37130), .I0(n8017[4]), .I1(n589_adj_3446), 
            .CO(n37131));
    SB_LUT4 add_3221_3_lut (.I0(GND_net), .I1(n12573[0]), .I2(n216), .I3(n36365), 
            .O(n11990[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3486_6 (.CI(n37577), .I0(n16627[3]), .I1(n558), .CO(n37578));
    SB_CARRY unary_minus_21_add_3_17 (.CI(n36025), .I0(GND_net), .I1(n60[15]), 
            .CO(n36026));
    SB_LUT4 add_3073_10_lut (.I0(GND_net), .I1(n8404[7]), .I2(GND_net), 
            .I3(n37484), .O(n8391[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3064_2_lut (.I0(GND_net), .I1(n38), .I2(n131_adj_3450), 
            .I3(GND_net), .O(n8229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3064_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3054_2 (.CI(GND_net), .I0(n8_adj_3433), .I1(n101), .CO(n36914));
    SB_CARRY add_3064_2 (.CI(GND_net), .I0(n38), .I1(n131_adj_3450), .CO(n37342));
    SB_LUT4 add_3055_6_lut (.I0(GND_net), .I1(n8017[3]), .I2(n492), .I3(n37129), 
            .O(n7986[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3221_3 (.CI(n36365), .I0(n12573[0]), .I1(n216), .CO(n36366));
    SB_LUT4 add_3221_2_lut (.I0(GND_net), .I1(n26_adj_3451), .I2(n119), 
            .I3(GND_net), .O(n11990[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_6 (.CI(n37129), .I0(n8017[3]), .I1(n492), .CO(n37130));
    SB_CARRY add_3221_2 (.CI(GND_net), .I0(n26_adj_3451), .I1(n119), .CO(n36365));
    SB_LUT4 add_3377_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(n36364), .O(n15224[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(\motor_state[3] ), 
            .I2(n66[3]), .I3(n36132), .O(\PID_CONTROLLER.err_31__N_2825 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_9_lut (.I0(GND_net), .I1(n583), .I2(GND_net), .I3(n36363), 
            .O(n15224[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_9 (.CI(n36363), .I0(n583), .I1(GND_net), .CO(n36364));
    SB_CARRY state_23__I_0_add_2_5 (.CI(n36132), .I0(\motor_state[3] ), 
            .I1(n66[3]), .CO(n36133));
    SB_LUT4 add_3377_8_lut (.I0(GND_net), .I1(n510), .I2(n545), .I3(n36362), 
            .O(n15224[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_10 (.CI(n37484), .I0(n8404[7]), .I1(GND_net), .CO(n37485));
    SB_LUT4 add_3063_22_lut (.I0(GND_net), .I1(n8229[19]), .I2(GND_net), 
            .I3(n37341), .O(n8206[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_21_lut (.I0(GND_net), .I1(n8229[18]), .I2(GND_net), 
            .I3(n37340), .O(n8206[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_26_lut (.I0(GND_net), .I1(n7063[1]), 
            .I2(n58[24]), .I3(n35910), .O(n57[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_5_lut (.I0(GND_net), .I1(n8017[2]), .I2(n395), .I3(n37128), 
            .O(n7986[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_8 (.CI(n36362), .I0(n510), .I1(n545), .CO(n36363));
    SB_LUT4 add_3377_7_lut (.I0(GND_net), .I1(n437_adj_3453), .I2(n472), 
            .I3(n36361), .O(n15224[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_5 (.CI(n37128), .I0(n8017[2]), .I1(n395), .CO(n37129));
    SB_CARRY add_3377_7 (.CI(n36361), .I0(n437_adj_3453), .I1(n472), .CO(n36362));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(\motor_state[2] ), 
            .I2(n66[2]), .I3(n36131), .O(\PID_CONTROLLER.err_31__N_2825 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n60[14]), 
            .I3(n36024), .O(n406)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_16 (.CI(n36024), .I0(GND_net), .I1(n60[14]), 
            .CO(n36025));
    SB_CARRY state_23__I_0_add_2_4 (.CI(n36131), .I0(\motor_state[2] ), 
            .I1(n66[2]), .CO(n36132));
    SB_LUT4 add_3377_6_lut (.I0(GND_net), .I1(n364_adj_3455), .I2(n399_c), 
            .I3(n36360), .O(n15224[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_2 (.CI(GND_net), .I0(n20_adj_3439), .I1(n89), 
            .CO(n37752));
    SB_LUT4 add_3254_16_lut (.I0(GND_net), .I1(n13254[13]), .I2(GND_net), 
            .I3(n36913), .O(n12730[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_26 (.CI(n35910), .I0(n7063[1]), .I1(n58[24]), 
            .CO(n35911));
    SB_LUT4 add_13_add_1_21902_add_1_25_lut (.I0(GND_net), .I1(n7063[0]), 
            .I2(n58[23]), .I3(n35909), .O(n57[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3254_15_lut (.I0(GND_net), .I1(n13254[12]), .I2(GND_net), 
            .I3(n36912), .O(n12730[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_6 (.CI(n36360), .I0(n364_adj_3455), .I1(n399_c), 
            .CO(n36361));
    SB_LUT4 add_3377_5_lut (.I0(GND_net), .I1(n291), .I2(n326), .I3(n36359), 
            .O(n15224[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_15 (.CI(n36912), .I0(n13254[12]), .I1(GND_net), 
            .CO(n36913));
    SB_CARRY add_3377_5 (.CI(n36359), .I0(n291), .I1(n326), .CO(n36360));
    SB_LUT4 mult_14_add_1215_24_lut (.I0(GND_net), .I1(n1801[21]), .I2(GND_net), 
            .I3(n37750), .O(n1800[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_24 (.CI(n37750), .I0(n1801[21]), .I1(GND_net), 
            .CO(n1699));
    SB_LUT4 mult_14_add_1215_23_lut (.I0(GND_net), .I1(n1801[20]), .I2(GND_net), 
            .I3(n37749), .O(n1800[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_24_lut (.I0(GND_net), .I1(n1797[21]), .I2(GND_net), 
            .I3(n37658), .O(n1796[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3486_5_lut (.I0(GND_net), .I1(n16627[2]), .I2(n464), .I3(n37576), 
            .O(n16618[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3486_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_9_lut (.I0(GND_net), .I1(n8404[6]), .I2(GND_net), 
            .I3(n37483), .O(n8391[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_21 (.CI(n37340), .I0(n8229[18]), .I1(GND_net), .CO(n37341));
    SB_LUT4 add_3055_4_lut (.I0(GND_net), .I1(n8017[1]), .I2(n298), .I3(n37127), 
            .O(n7986[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_4 (.CI(n37127), .I0(n8017[1]), .I1(n298), .CO(n37128));
    SB_LUT4 add_3063_20_lut (.I0(GND_net), .I1(n8229[17]), .I2(GND_net), 
            .I3(n37339), .O(n8206[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3055_3_lut (.I0(GND_net), .I1(n8017[0]), .I2(n201), .I3(n37126), 
            .O(n7986[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_3 (.CI(n37126), .I0(n8017[0]), .I1(n201), .CO(n37127));
    SB_CARRY add_3486_5 (.CI(n37576), .I0(n16627[2]), .I1(n464), .CO(n37577));
    SB_CARRY add_3073_9 (.CI(n37483), .I0(n8404[6]), .I1(GND_net), .CO(n37484));
    SB_CARRY add_3063_20 (.CI(n37339), .I0(n8229[17]), .I1(GND_net), .CO(n37340));
    SB_LUT4 add_3055_2_lut (.I0(GND_net), .I1(n11_adj_3457), .I2(n104), 
            .I3(GND_net), .O(n7986[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3055_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3055_2 (.CI(GND_net), .I0(n11_adj_3457), .I1(n104), .CO(n37126));
    SB_LUT4 add_3063_19_lut (.I0(GND_net), .I1(n8229[16]), .I2(GND_net), 
            .I3(n37338), .O(n8206[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_32_lut (.I0(n69[25]), .I1(n7954[29]), .I2(GND_net), 
            .I3(n37125), .O(n7059[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_12_add_2137_31_lut (.I0(GND_net), .I1(n7954[28]), .I2(GND_net), 
            .I3(n37124), .O(n191[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_24 (.CI(n37658), .I0(n1797[21]), .I1(GND_net), 
            .CO(n1683));
    SB_LUT4 add_3486_4_lut (.I0(GND_net), .I1(n16627[1]), .I2(n370), .I3(n37575), 
            .O(n16618[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3486_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_8_lut (.I0(GND_net), .I1(n8404[5]), .I2(n740), .I3(n37482), 
            .O(n8391[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_19 (.CI(n37338), .I0(n8229[16]), .I1(GND_net), .CO(n37339));
    SB_CARRY mult_12_add_2137_31 (.CI(n37124), .I0(n7954[28]), .I1(GND_net), 
            .CO(n37125));
    SB_LUT4 mult_12_add_2137_30_lut (.I0(GND_net), .I1(n7954[27]), .I2(GND_net), 
            .I3(n37123), .O(n191[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_18_lut (.I0(GND_net), .I1(n8229[15]), .I2(GND_net), 
            .I3(n37337), .O(n8206[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_30 (.CI(n37123), .I0(n7954[27]), .I1(GND_net), 
            .CO(n37124));
    SB_LUT4 mult_12_add_2137_29_lut (.I0(GND_net), .I1(n7954[26]), .I2(GND_net), 
            .I3(n37122), .O(n191[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3486_4 (.CI(n37575), .I0(n16627[1]), .I1(n370), .CO(n37576));
    SB_CARRY add_3073_8 (.CI(n37482), .I0(n8404[5]), .I1(n740), .CO(n37483));
    SB_CARRY add_3063_18 (.CI(n37337), .I0(n8229[15]), .I1(GND_net), .CO(n37338));
    SB_CARRY mult_12_add_2137_29 (.CI(n37122), .I0(n7954[26]), .I1(GND_net), 
            .CO(n37123));
    SB_LUT4 mult_12_add_2137_28_lut (.I0(GND_net), .I1(n7954[25]), .I2(GND_net), 
            .I3(n37121), .O(n191[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_17_lut (.I0(GND_net), .I1(n8229[14]), .I2(GND_net), 
            .I3(n37336), .O(n8206[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_28 (.CI(n37121), .I0(n7954[25]), .I1(GND_net), 
            .CO(n37122));
    SB_CARRY mult_14_add_1215_23 (.CI(n37749), .I0(n1801[20]), .I1(GND_net), 
            .CO(n37750));
    SB_LUT4 mult_14_add_1211_23_lut (.I0(GND_net), .I1(n1797[20]), .I2(GND_net), 
            .I3(n37657), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3486_3_lut (.I0(GND_net), .I1(n16627[0]), .I2(n276), .I3(n37574), 
            .O(n16618[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3486_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_7_lut (.I0(GND_net), .I1(n8404[4]), .I2(n643), .I3(n37481), 
            .O(n8391[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_17 (.CI(n37336), .I0(n8229[14]), .I1(GND_net), .CO(n37337));
    SB_LUT4 add_3063_16_lut (.I0(GND_net), .I1(n8229[13]), .I2(GND_net), 
            .I3(n37335), .O(n8206[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3486_3 (.CI(n37574), .I0(n16627[0]), .I1(n276), .CO(n37575));
    SB_CARRY add_3073_7 (.CI(n37481), .I0(n8404[4]), .I1(n643), .CO(n37482));
    SB_CARRY add_3063_16 (.CI(n37335), .I0(n8229[13]), .I1(GND_net), .CO(n37336));
    SB_LUT4 add_3063_15_lut (.I0(GND_net), .I1(n8229[12]), .I2(GND_net), 
            .I3(n37334), .O(n8206[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_23 (.CI(n37657), .I0(n1797[20]), .I1(GND_net), 
            .CO(n37658));
    SB_LUT4 add_3486_2_lut (.I0(GND_net), .I1(n86_adj_3389), .I2(n182), 
            .I3(GND_net), .O(n16618[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3486_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_6_lut (.I0(GND_net), .I1(n8404[3]), .I2(n546), .I3(n37480), 
            .O(n8391[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_15 (.CI(n37334), .I0(n8229[12]), .I1(GND_net), .CO(n37335));
    SB_LUT4 add_3063_14_lut (.I0(GND_net), .I1(n8229[11]), .I2(GND_net), 
            .I3(n37333), .O(n8206[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3486_2 (.CI(GND_net), .I0(n86_adj_3389), .I1(n182), .CO(n37574));
    SB_CARRY add_3073_6 (.CI(n37480), .I0(n8404[3]), .I1(n546), .CO(n37481));
    SB_CARRY add_3063_14 (.CI(n37333), .I0(n8229[11]), .I1(GND_net), .CO(n37334));
    SB_LUT4 add_3063_13_lut (.I0(GND_net), .I1(n8229[10]), .I2(GND_net), 
            .I3(n37332), .O(n8206[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_22_lut (.I0(GND_net), .I1(n1801[19]), .I2(GND_net), 
            .I3(n37748), .O(n1800[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_22_lut (.I0(GND_net), .I1(n1797[19]), .I2(GND_net), 
            .I3(n37656), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_15_lut (.I0(GND_net), .I1(n16029[12]), .I2(GND_net), 
            .I3(n37573), .O(n15848[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_5_lut (.I0(GND_net), .I1(n8404[2]), .I2(n449_c), 
            .I3(n37479), .O(n8391[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_13 (.CI(n37332), .I0(n8229[10]), .I1(GND_net), .CO(n37333));
    SB_LUT4 mult_12_add_2137_27_lut (.I0(GND_net), .I1(n7954[24]), .I2(GND_net), 
            .I3(n37120), .O(n191[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_12_lut (.I0(GND_net), .I1(n8229[9]), .I2(GND_net), 
            .I3(n37331), .O(n8206[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_27 (.CI(n37120), .I0(n7954[24]), .I1(GND_net), 
            .CO(n37121));
    SB_LUT4 mult_12_add_2137_26_lut (.I0(GND_net), .I1(n7954[23]), .I2(GND_net), 
            .I3(n37119), .O(n191[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3073_5 (.CI(n37479), .I0(n8404[2]), .I1(n449_c), .CO(n37480));
    SB_CARRY add_3063_12 (.CI(n37331), .I0(n8229[9]), .I1(GND_net), .CO(n37332));
    SB_CARRY mult_12_add_2137_26 (.CI(n37119), .I0(n7954[23]), .I1(GND_net), 
            .CO(n37120));
    SB_LUT4 add_3254_14_lut (.I0(GND_net), .I1(n13254[11]), .I2(GND_net), 
            .I3(n36911), .O(n12730[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_25_lut (.I0(GND_net), .I1(n7954[22]), .I2(GND_net), 
            .I3(n37118), .O(n191[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_14 (.CI(n36911), .I0(n13254[11]), .I1(GND_net), 
            .CO(n36912));
    SB_LUT4 add_3254_13_lut (.I0(GND_net), .I1(n13254[10]), .I2(GND_net), 
            .I3(n36910), .O(n12730[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_11_lut (.I0(GND_net), .I1(n8229[8]), .I2(GND_net), 
            .I3(n37330), .O(n8206[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_25 (.CI(n37118), .I0(n7954[22]), .I1(GND_net), 
            .CO(n37119));
    SB_CARRY add_3254_13 (.CI(n36910), .I0(n13254[10]), .I1(GND_net), 
            .CO(n36911));
    SB_LUT4 add_3254_12_lut (.I0(GND_net), .I1(n13254[9]), .I2(GND_net), 
            .I3(n36909), .O(n12730[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_24_lut (.I0(GND_net), .I1(n7954[21]), .I2(GND_net), 
            .I3(n37117), .O(n191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_12 (.CI(n36909), .I0(n13254[9]), .I1(GND_net), .CO(n36910));
    SB_LUT4 add_3254_11_lut (.I0(GND_net), .I1(n13254[8]), .I2(GND_net), 
            .I3(n36908), .O(n12730[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_14_lut (.I0(GND_net), .I1(n16029[11]), .I2(GND_net), 
            .I3(n37572), .O(n15848[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_4_lut (.I0(GND_net), .I1(n8404[1]), .I2(n352), .I3(n37478), 
            .O(n8391[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_11 (.CI(n37330), .I0(n8229[8]), .I1(GND_net), .CO(n37331));
    SB_LUT4 add_3063_10_lut (.I0(GND_net), .I1(n8229[7]), .I2(GND_net), 
            .I3(n37329), .O(n8206[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_11 (.CI(n36908), .I0(n13254[8]), .I1(GND_net), .CO(n36909));
    SB_CARRY mult_12_add_2137_24 (.CI(n37117), .I0(n7954[21]), .I1(GND_net), 
            .CO(n37118));
    SB_LUT4 mult_12_add_2137_23_lut (.I0(GND_net), .I1(n7954[20]), .I2(GND_net), 
            .I3(n37116), .O(n191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_10 (.CI(n37329), .I0(n8229[7]), .I1(GND_net), .CO(n37330));
    SB_CARRY mult_12_add_2137_23 (.CI(n37116), .I0(n7954[20]), .I1(GND_net), 
            .CO(n37117));
    SB_LUT4 mult_12_add_2137_22_lut (.I0(GND_net), .I1(n7954[19]), .I2(GND_net), 
            .I3(n37115), .O(n191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_22 (.CI(n37748), .I0(n1801[19]), .I1(GND_net), 
            .CO(n37749));
    SB_CARRY mult_12_add_2137_22 (.CI(n37115), .I0(n7954[19]), .I1(GND_net), 
            .CO(n37116));
    SB_CARRY add_3073_4 (.CI(n37478), .I0(n8404[1]), .I1(n352), .CO(n37479));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(\motor_state[1] ), 
            .I2(n66[1]), .I3(n36130), .O(\PID_CONTROLLER.err_31__N_2825 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_9_lut (.I0(GND_net), .I1(n8229[6]), .I2(GND_net), 
            .I3(n37328), .O(n8206[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_21_lut (.I0(GND_net), .I1(n7954[18]), .I2(GND_net), 
            .I3(n37114), .O(n191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3254_10_lut (.I0(GND_net), .I1(n13254[7]), .I2(GND_net), 
            .I3(n36907), .O(n12730[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_10 (.CI(n36907), .I0(n13254[7]), .I1(GND_net), .CO(n36908));
    SB_CARRY mult_12_add_2137_21 (.CI(n37114), .I0(n7954[18]), .I1(GND_net), 
            .CO(n37115));
    SB_LUT4 add_3254_9_lut (.I0(GND_net), .I1(n13254[6]), .I2(GND_net), 
            .I3(n36906), .O(n12730[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_9 (.CI(n36906), .I0(n13254[6]), .I1(GND_net), .CO(n36907));
    SB_LUT4 add_3377_4_lut (.I0(GND_net), .I1(n218_adj_3463), .I2(n253), 
            .I3(n36358), .O(n15224[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_9 (.CI(n37328), .I0(n8229[6]), .I1(GND_net), .CO(n37329));
    SB_LUT4 mult_12_add_2137_20_lut (.I0(GND_net), .I1(n7954[17]), .I2(GND_net), 
            .I3(n37113), .O(n191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3254_8_lut (.I0(GND_net), .I1(n13254[5]), .I2(n545), .I3(n36905), 
            .O(n12730[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_8 (.CI(n36905), .I0(n13254[5]), .I1(n545), .CO(n36906));
    SB_CARRY mult_12_add_2137_20 (.CI(n37113), .I0(n7954[17]), .I1(GND_net), 
            .CO(n37114));
    SB_LUT4 add_3254_7_lut (.I0(GND_net), .I1(n13254[4]), .I2(n472), .I3(n36904), 
            .O(n12730[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_7 (.CI(n36904), .I0(n13254[4]), .I1(n472), .CO(n36905));
    SB_CARRY mult_14_add_1211_22 (.CI(n37656), .I0(n1797[19]), .I1(GND_net), 
            .CO(n37657));
    SB_CARRY add_3416_14 (.CI(n37572), .I0(n16029[11]), .I1(GND_net), 
            .CO(n37573));
    SB_LUT4 mult_12_add_2137_19_lut (.I0(GND_net), .I1(n7954[16]), .I2(GND_net), 
            .I3(n37112), .O(n191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_3_lut (.I0(GND_net), .I1(n8404[0]), .I2(n255), .I3(n37477), 
            .O(n8391[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_8_lut (.I0(GND_net), .I1(n8229[5]), .I2(n710), .I3(n37327), 
            .O(n8206[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_19 (.CI(n37112), .I0(n7954[16]), .I1(GND_net), 
            .CO(n37113));
    SB_LUT4 mult_12_add_2137_18_lut (.I0(GND_net), .I1(n7954[15]), .I2(GND_net), 
            .I3(n37111), .O(n191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_21_lut (.I0(GND_net), .I1(n1801[18]), .I2(GND_net), 
            .I3(n37747), .O(n1800[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n60[13]), 
            .I3(n36023), .O(n407)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_18 (.CI(n37111), .I0(n7954[15]), .I1(GND_net), 
            .CO(n37112));
    SB_LUT4 add_3254_6_lut (.I0(GND_net), .I1(n13254[3]), .I2(n399_c), 
            .I3(n36903), .O(n12730[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_4 (.CI(n36358), .I0(n218_adj_3463), .I1(n253), .CO(n36359));
    SB_CARRY add_3254_6 (.CI(n36903), .I0(n13254[3]), .I1(n399_c), .CO(n36904));
    SB_LUT4 add_3377_3_lut (.I0(GND_net), .I1(n145), .I2(n180), .I3(n36357), 
            .O(n15224[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_3 (.CI(n36357), .I0(n145), .I1(n180), .CO(n36358));
    SB_CARRY add_3063_8 (.CI(n37327), .I0(n8229[5]), .I1(n710), .CO(n37328));
    SB_CARRY state_23__I_0_add_2_3 (.CI(n36130), .I0(\motor_state[1] ), 
            .I1(n66[1]), .CO(n36131));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(\motor_state[0] ), 
            .I2(n66[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_31__N_2825 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3254_5_lut (.I0(GND_net), .I1(n13254[2]), .I2(n326), .I3(n36902), 
            .O(n12730[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_5 (.CI(n36902), .I0(n13254[2]), .I1(n326), .CO(n36903));
    SB_LUT4 add_3254_4_lut (.I0(GND_net), .I1(n13254[1]), .I2(n253), .I3(n36901), 
            .O(n12730[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_17_lut (.I0(GND_net), .I1(n7954[14]), .I2(GND_net), 
            .I3(n37110), .O(n191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_17 (.CI(n37110), .I0(n7954[14]), .I1(GND_net), 
            .CO(n37111));
    SB_CARRY unary_minus_21_add_3_15 (.CI(n36023), .I0(GND_net), .I1(n60[13]), 
            .CO(n36024));
    SB_LUT4 unary_minus_21_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n60[12]), 
            .I3(n36022), .O(n67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_16_lut (.I0(GND_net), .I1(n7954[13]), .I2(GND_net), 
            .I3(n37109), .O(n191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3377_2_lut (.I0(GND_net), .I1(n72), .I2(n107), .I3(GND_net), 
            .O(n15224[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3377_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_4 (.CI(n36901), .I0(n13254[1]), .I1(n253), .CO(n36902));
    SB_CARRY mult_12_add_2137_16 (.CI(n37109), .I0(n7954[13]), .I1(GND_net), 
            .CO(n37110));
    SB_CARRY mult_14_add_1215_21 (.CI(n37747), .I0(n1801[18]), .I1(GND_net), 
            .CO(n37748));
    SB_CARRY add_3073_3 (.CI(n37477), .I0(n8404[0]), .I1(n255), .CO(n37478));
    SB_LUT4 add_3063_7_lut (.I0(GND_net), .I1(n8229[4]), .I2(n613), .I3(n37326), 
            .O(n8206[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3254_3_lut (.I0(GND_net), .I1(n13254[0]), .I2(n180), .I3(n36900), 
            .O(n12730[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3377_2 (.CI(GND_net), .I0(n72), .I1(n107), .CO(n36357));
    SB_CARRY add_3254_3 (.CI(n36900), .I0(n13254[0]), .I1(n180), .CO(n36901));
    SB_LUT4 add_3246_24_lut (.I0(GND_net), .I1(n13107[21]), .I2(GND_net), 
            .I3(n36356), .O(n12573[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_15_lut (.I0(GND_net), .I1(n7954[12]), .I2(GND_net), 
            .I3(n37108), .O(n191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(\motor_state[0] ), 
            .I1(n66[0]), .CO(n36130));
    SB_LUT4 add_3254_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n12730[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3254_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3254_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n36900));
    SB_CARRY mult_12_add_2137_15 (.CI(n37108), .I0(n7954[12]), .I1(GND_net), 
            .CO(n37109));
    SB_LUT4 Kd_delay_counter_1013_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[6]), .I3(n36899), .O(n70[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1013_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1013_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[5]), .I3(n36898), .O(n70[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1013_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_7 (.CI(n37326), .I0(n8229[4]), .I1(n613), .CO(n37327));
    SB_LUT4 mult_12_add_2137_14_lut (.I0(GND_net), .I1(n7954[11]), .I2(GND_net), 
            .I3(n37107), .O(n191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1013_add_4_7 (.CI(n36898), .I0(GND_net), .I1(Kd_delay_counter[5]), 
            .CO(n36899));
    SB_LUT4 Kd_delay_counter_1013_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[4]), .I3(n36897), .O(n70[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1013_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_14 (.CI(n37107), .I0(n7954[11]), .I1(GND_net), 
            .CO(n37108));
    SB_CARRY unary_minus_21_add_3_14 (.CI(n36022), .I0(GND_net), .I1(n60[12]), 
            .CO(n36023));
    SB_CARRY Kd_delay_counter_1013_add_4_6 (.CI(n36897), .I0(GND_net), .I1(Kd_delay_counter[4]), 
            .CO(n36898));
    SB_LUT4 mult_12_add_2137_13_lut (.I0(GND_net), .I1(n7954[10]), .I2(GND_net), 
            .I3(n37106), .O(n191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_6_lut (.I0(GND_net), .I1(n8229[3]), .I2(n516_adj_3471), 
            .I3(n37325), .O(n8206[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_13 (.CI(n37106), .I0(n7954[10]), .I1(GND_net), 
            .CO(n37107));
    SB_LUT4 sub_11_add_2_27_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n63[26]), .I3(n36129), .O(n69[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1013_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[3]), .I3(n36896), .O(n70[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1013_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n60[11]), 
            .I3(n36021), .O(n67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1013_add_4_5 (.CI(n36896), .I0(GND_net), .I1(Kd_delay_counter[3]), 
            .CO(n36897));
    SB_LUT4 add_3416_13_lut (.I0(GND_net), .I1(n16029[10]), .I2(GND_net), 
            .I3(n37571), .O(n15848[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1013_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[2]), .I3(n36895), .O(n70[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1013_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3073_2_lut (.I0(GND_net), .I1(n65), .I2(n158), .I3(GND_net), 
            .O(n8391[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3073_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_6 (.CI(n37325), .I0(n8229[3]), .I1(n516_adj_3471), 
            .CO(n37326));
    SB_LUT4 mult_12_add_2137_12_lut (.I0(GND_net), .I1(n7954[9]), .I2(GND_net), 
            .I3(n37105), .O(n191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_26_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n63[26]), .I3(n36128), .O(n69[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_12 (.CI(n37105), .I0(n7954[9]), .I1(GND_net), 
            .CO(n37106));
    SB_CARRY unary_minus_21_add_3_13 (.CI(n36021), .I0(GND_net), .I1(n60[11]), 
            .CO(n36022));
    SB_LUT4 add_3246_23_lut (.I0(GND_net), .I1(n13107[20]), .I2(GND_net), 
            .I3(n36355), .O(n12573[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_5_lut (.I0(GND_net), .I1(n8229[2]), .I2(n419), .I3(n37324), 
            .O(n8206[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_11_lut (.I0(GND_net), .I1(n7954[8]), .I2(GND_net), 
            .I3(n37104), .O(n191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_23 (.CI(n36355), .I0(n13107[20]), .I1(GND_net), 
            .CO(n36356));
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n60[10]), 
            .I3(n36020), .O(n67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1013_add_4_4 (.CI(n36895), .I0(GND_net), .I1(Kd_delay_counter[2]), 
            .CO(n36896));
    SB_CARRY mult_12_add_2137_11 (.CI(n37104), .I0(n7954[8]), .I1(GND_net), 
            .CO(n37105));
    SB_CARRY add_3073_2 (.CI(GND_net), .I0(n65), .I1(n158), .CO(n37477));
    SB_CARRY sub_11_add_2_26 (.CI(n36128), .I0(\PID_CONTROLLER.err_prev[31] ), 
            .I1(n63[26]), .CO(n36129));
    SB_LUT4 sub_11_add_2_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[23] ), 
            .I2(n63[23]), .I3(n36127), .O(n69[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_13 (.CI(n37571), .I0(n16029[10]), .I1(GND_net), 
            .CO(n37572));
    SB_CARRY add_3063_5 (.CI(n37324), .I0(n8229[2]), .I1(n419), .CO(n37325));
    SB_LUT4 mult_12_add_2137_10_lut (.I0(GND_net), .I1(n7954[7]), .I2(GND_net), 
            .I3(n37103), .O(n191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1013_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[1]), .I3(n36894), .O(n70[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1013_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1013_add_4_3 (.CI(n36894), .I0(GND_net), .I1(Kd_delay_counter[1]), 
            .CO(n36895));
    SB_CARRY mult_12_add_2137_10 (.CI(n37103), .I0(n7954[7]), .I1(GND_net), 
            .CO(n37104));
    SB_LUT4 Kd_delay_counter_1013_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[0]), .I3(VCC_net), .O(n70[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1013_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1013_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(Kd_delay_counter[0]), .CO(n36894));
    SB_LUT4 add_3063_4_lut (.I0(GND_net), .I1(n8229[1]), .I2(n322), .I3(n37323), 
            .O(n8206[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_9_lut (.I0(GND_net), .I1(n7954[6]), .I2(GND_net), 
            .I3(n37102), .O(n191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_9 (.CI(n37102), .I0(n7954[6]), .I1(GND_net), 
            .CO(n37103));
    SB_LUT4 mult_14_add_1215_20_lut (.I0(GND_net), .I1(n1801[17]), .I2(GND_net), 
            .I3(n37746), .O(n1800[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_21_lut (.I0(GND_net), .I1(n1797[18]), .I2(GND_net), 
            .I3(n37655), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_12_lut (.I0(GND_net), .I1(n16029[9]), .I2(GND_net), 
            .I3(n37570), .O(n15848[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_13_lut (.I0(GND_net), .I1(n8391[10]), .I2(GND_net), 
            .I3(n37476), .O(n8377[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_4 (.CI(n37323), .I0(n8229[1]), .I1(n322), .CO(n37324));
    SB_LUT4 mult_12_add_2137_8_lut (.I0(GND_net), .I1(n7954[5]), .I2(n680), 
            .I3(n37101), .O(n191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_3_lut (.I0(GND_net), .I1(n8229[0]), .I2(n225_adj_3485), 
            .I3(n37322), .O(n8206[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_12_lut (.I0(GND_net), .I1(n8391[9]), .I2(GND_net), 
            .I3(n37475), .O(n8377[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3063_3 (.CI(n37322), .I0(n8229[0]), .I1(n225_adj_3485), 
            .CO(n37323));
    SB_CARRY mult_12_add_2137_8 (.CI(n37101), .I0(n7954[5]), .I1(n680), 
            .CO(n37102));
    SB_LUT4 add_3246_22_lut (.I0(GND_net), .I1(n13107[19]), .I2(GND_net), 
            .I3(n36354), .O(n12573[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_7_lut (.I0(GND_net), .I1(n7954[4]), .I2(n583_adj_3486), 
            .I3(n37100), .O(n191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_22 (.CI(n36354), .I0(n13107[19]), .I1(GND_net), 
            .CO(n36355));
    SB_LUT4 add_3246_21_lut (.I0(GND_net), .I1(n13107[18]), .I2(GND_net), 
            .I3(n36353), .O(n12573[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_21 (.CI(n36353), .I0(n13107[18]), .I1(GND_net), 
            .CO(n36354));
    SB_CARRY sub_11_add_2_25 (.CI(n36127), .I0(\PID_CONTROLLER.err_prev[23] ), 
            .I1(n63[23]), .CO(n36128));
    SB_LUT4 add_3246_20_lut (.I0(GND_net), .I1(n13107[17]), .I2(GND_net), 
            .I3(n36352), .O(n12573[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3063_2_lut (.I0(GND_net), .I1(n35_adj_3487), .I2(n128), 
            .I3(GND_net), .O(n8206[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3063_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_7 (.CI(n37100), .I0(n7954[4]), .I1(n583_adj_3486), 
            .CO(n37101));
    SB_CARRY add_3246_20 (.CI(n36352), .I0(n13107[17]), .I1(GND_net), 
            .CO(n36353));
    SB_LUT4 add_3246_19_lut (.I0(GND_net), .I1(n13107[16]), .I2(GND_net), 
            .I3(n36351), .O(n12573[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_6_lut (.I0(GND_net), .I1(n7954[3]), .I2(n486), 
            .I3(n37099), .O(n191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_19 (.CI(n36351), .I0(n13107[16]), .I1(GND_net), 
            .CO(n36352));
    SB_LUT4 sub_11_add_2_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[22] ), 
            .I2(n63[22]), .I3(n36126), .O(n69[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_24 (.CI(n36126), .I0(\PID_CONTROLLER.err_prev[22] ), 
            .I1(n63[22]), .CO(n36127));
    SB_LUT4 add_3246_18_lut (.I0(GND_net), .I1(n13107[15]), .I2(GND_net), 
            .I3(n36350), .O(n12573[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_18 (.CI(n36350), .I0(n13107[15]), .I1(GND_net), 
            .CO(n36351));
    SB_LUT4 sub_11_add_2_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[21] ), 
            .I2(n63[21]), .I3(n36125), .O(n69[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_12 (.CI(n36020), .I0(GND_net), .I1(n60[10]), 
            .CO(n36021));
    SB_CARRY sub_11_add_2_23 (.CI(n36125), .I0(\PID_CONTROLLER.err_prev[21] ), 
            .I1(n63[21]), .CO(n36126));
    SB_LUT4 add_3246_17_lut (.I0(GND_net), .I1(n13107[14]), .I2(GND_net), 
            .I3(n36349), .O(n12573[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_12 (.CI(n37570), .I0(n16029[9]), .I1(GND_net), .CO(n37571));
    SB_CARRY add_3072_12 (.CI(n37475), .I0(n8391[9]), .I1(GND_net), .CO(n37476));
    SB_CARRY add_3063_2 (.CI(GND_net), .I0(n35_adj_3487), .I1(n128), .CO(n37322));
    SB_LUT4 add_3062_23_lut (.I0(GND_net), .I1(n8206[20]), .I2(GND_net), 
            .I3(n37321), .O(n8182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3072_11_lut (.I0(GND_net), .I1(n8391[8]), .I2(GND_net), 
            .I3(n37474), .O(n8377[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_22_lut (.I0(GND_net), .I1(n8206[19]), .I2(GND_net), 
            .I3(n37320), .O(n8182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_6 (.CI(n37099), .I0(n7954[3]), .I1(n486), 
            .CO(n37100));
    SB_CARRY add_3246_17 (.CI(n36349), .I0(n13107[14]), .I1(GND_net), 
            .CO(n36350));
    SB_LUT4 add_3246_16_lut (.I0(GND_net), .I1(n13107[13]), .I2(GND_net), 
            .I3(n36348), .O(n12573[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_5_lut (.I0(GND_net), .I1(n7954[2]), .I2(n389), 
            .I3(n37098), .O(n191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_16 (.CI(n36348), .I0(n13107[13]), .I1(GND_net), 
            .CO(n36349));
    SB_LUT4 sub_11_add_2_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[20] ), 
            .I2(n63[20]), .I3(n36124), .O(n69[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3246_15_lut (.I0(GND_net), .I1(n13107[12]), .I2(GND_net), 
            .I3(n36347), .O(n12573[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_15 (.CI(n36347), .I0(n13107[12]), .I1(GND_net), 
            .CO(n36348));
    SB_CARRY sub_11_add_2_22 (.CI(n36124), .I0(\PID_CONTROLLER.err_prev[20] ), 
            .I1(n63[20]), .CO(n36125));
    SB_LUT4 add_3246_14_lut (.I0(GND_net), .I1(n13107[11]), .I2(GND_net), 
            .I3(n36346), .O(n12573[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_22 (.CI(n37320), .I0(n8206[19]), .I1(GND_net), .CO(n37321));
    SB_CARRY mult_12_add_2137_5 (.CI(n37098), .I0(n7954[2]), .I1(n389), 
            .CO(n37099));
    SB_CARRY add_3246_14 (.CI(n36346), .I0(n13107[11]), .I1(GND_net), 
            .CO(n36347));
    SB_LUT4 add_3246_13_lut (.I0(GND_net), .I1(n13107[10]), .I2(GND_net), 
            .I3(n36345), .O(n12573[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_4_lut (.I0(GND_net), .I1(n7954[1]), .I2(n292), 
            .I3(n37097), .O(n191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_13 (.CI(n36345), .I0(n13107[10]), .I1(GND_net), 
            .CO(n36346));
    SB_LUT4 sub_11_add_2_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[19] ), 
            .I2(n63[19]), .I3(n36123), .O(n69[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n60[9]), 
            .I3(n36019), .O(n67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n36019), .I0(GND_net), .I1(n60[9]), 
            .CO(n36020));
    SB_CARRY sub_11_add_2_21 (.CI(n36123), .I0(\PID_CONTROLLER.err_prev[19] ), 
            .I1(n63[19]), .CO(n36124));
    SB_LUT4 add_3246_12_lut (.I0(GND_net), .I1(n13107[9]), .I2(GND_net), 
            .I3(n36344), .O(n12573[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_12 (.CI(n36344), .I0(n13107[9]), .I1(GND_net), .CO(n36345));
    SB_LUT4 sub_11_add_2_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[18] ), 
            .I2(n63[18]), .I3(n36122), .O(n69[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n60[8]), 
            .I3(n36018), .O(n67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_10 (.CI(n36018), .I0(GND_net), .I1(n60[8]), 
            .CO(n36019));
    SB_CARRY sub_11_add_2_20 (.CI(n36122), .I0(\PID_CONTROLLER.err_prev[18] ), 
            .I1(n63[18]), .CO(n36123));
    SB_LUT4 add_3246_11_lut (.I0(GND_net), .I1(n13107[8]), .I2(GND_net), 
            .I3(n36343), .O(n12573[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_21 (.CI(n37655), .I0(n1797[18]), .I1(GND_net), 
            .CO(n37656));
    SB_LUT4 add_3416_11_lut (.I0(GND_net), .I1(n16029[8]), .I2(GND_net), 
            .I3(n37569), .O(n15848[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_11 (.CI(n37474), .I0(n8391[8]), .I1(GND_net), .CO(n37475));
    SB_LUT4 add_3062_21_lut (.I0(GND_net), .I1(n8206[18]), .I2(GND_net), 
            .I3(n37319), .O(n8182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_21 (.CI(n37319), .I0(n8206[18]), .I1(GND_net), .CO(n37320));
    SB_LUT4 add_3072_10_lut (.I0(GND_net), .I1(n8391[7]), .I2(GND_net), 
            .I3(n37473), .O(n8377[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_20_lut (.I0(GND_net), .I1(n8206[17]), .I2(GND_net), 
            .I3(n37318), .O(n8182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_4 (.CI(n37097), .I0(n7954[1]), .I1(n292), 
            .CO(n37098));
    SB_CARRY add_3246_11 (.CI(n36343), .I0(n13107[8]), .I1(GND_net), .CO(n36344));
    SB_LUT4 add_3246_10_lut (.I0(GND_net), .I1(n13107[7]), .I2(GND_net), 
            .I3(n36342), .O(n12573[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_3_lut (.I0(GND_net), .I1(n7954[0]), .I2(n195), 
            .I3(n37096), .O(n191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_10 (.CI(n36342), .I0(n13107[7]), .I1(GND_net), .CO(n36343));
    SB_LUT4 sub_11_add_2_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[17] ), 
            .I2(n63[17]), .I3(n36121), .O(n69[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3246_9_lut (.I0(GND_net), .I1(n13107[6]), .I2(GND_net), 
            .I3(n36341), .O(n12573[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_9 (.CI(n36341), .I0(n13107[6]), .I1(GND_net), .CO(n36342));
    SB_CARRY sub_11_add_2_19 (.CI(n36121), .I0(\PID_CONTROLLER.err_prev[17] ), 
            .I1(n63[17]), .CO(n36122));
    SB_LUT4 add_3246_8_lut (.I0(GND_net), .I1(n13107[5]), .I2(n704), .I3(n36340), 
            .O(n12573[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_20 (.CI(n37318), .I0(n8206[17]), .I1(GND_net), .CO(n37319));
    SB_CARRY mult_12_add_2137_3 (.CI(n37096), .I0(n7954[0]), .I1(n195), 
            .CO(n37097));
    SB_CARRY add_3246_8 (.CI(n36340), .I0(n13107[5]), .I1(n704), .CO(n36341));
    SB_LUT4 add_3246_7_lut (.I0(GND_net), .I1(n13107[4]), .I2(n607), .I3(n36339), 
            .O(n12573[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3496), .I2(n98), 
            .I3(GND_net), .O(n191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_7 (.CI(n36339), .I0(n13107[4]), .I1(n607), .CO(n36340));
    SB_LUT4 sub_11_add_2_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[16] ), 
            .I2(n63[16]), .I3(n36120), .O(n69[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n60[7]), 
            .I3(n36017), .O(n413)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_18 (.CI(n36120), .I0(\PID_CONTROLLER.err_prev[16] ), 
            .I1(n63[16]), .CO(n36121));
    SB_LUT4 add_3246_6_lut (.I0(GND_net), .I1(n13107[3]), .I2(n510_adj_3498), 
            .I3(n36338), .O(n12573[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_6 (.CI(n36338), .I0(n13107[3]), .I1(n510_adj_3498), 
            .CO(n36339));
    SB_LUT4 sub_11_add_2_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[15] ), 
            .I2(n63[15]), .I3(n36119), .O(n69[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_9 (.CI(n36017), .I0(GND_net), .I1(n60[7]), 
            .CO(n36018));
    SB_CARRY sub_11_add_2_17 (.CI(n36119), .I0(\PID_CONTROLLER.err_prev[15] ), 
            .I1(n63[15]), .CO(n36120));
    SB_LUT4 add_3246_5_lut (.I0(GND_net), .I1(n13107[2]), .I2(n413_adj_3500), 
            .I3(n36337), .O(n12573[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_11 (.CI(n37569), .I0(n16029[8]), .I1(GND_net), .CO(n37570));
    SB_CARRY add_3072_10 (.CI(n37473), .I0(n8391[7]), .I1(GND_net), .CO(n37474));
    SB_LUT4 add_3062_19_lut (.I0(GND_net), .I1(n8206[16]), .I2(GND_net), 
            .I3(n37317), .O(n8182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_19 (.CI(n37317), .I0(n8206[16]), .I1(GND_net), .CO(n37318));
    SB_LUT4 add_3072_9_lut (.I0(GND_net), .I1(n8391[6]), .I2(GND_net), 
            .I3(n37472), .O(n8377[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_18_lut (.I0(GND_net), .I1(n8206[15]), .I2(GND_net), 
            .I3(n37316), .O(n8182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_2 (.CI(GND_net), .I0(n5_adj_3496), .I1(n98), 
            .CO(n37096));
    SB_CARRY add_3246_5 (.CI(n36337), .I0(n13107[2]), .I1(n413_adj_3500), 
            .CO(n36338));
    SB_LUT4 add_3246_4_lut (.I0(GND_net), .I1(n13107[1]), .I2(n316), .I3(n36336), 
            .O(n12573[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_21_lut (.I0(GND_net), .I1(n10116[18]), .I2(GND_net), 
            .I3(n37095), .O(n9325[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_4 (.CI(n36336), .I0(n13107[1]), .I1(n316), .CO(n36337));
    SB_LUT4 sub_11_add_2_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[14] ), 
            .I2(n63[14]), .I3(n36118), .O(n69[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3246_3_lut (.I0(GND_net), .I1(n13107[0]), .I2(n219_adj_3502), 
            .I3(n36335), .O(n12573[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3246_3 (.CI(n36335), .I0(n13107[0]), .I1(n219_adj_3502), 
            .CO(n36336));
    SB_LUT4 mult_14_add_1211_20_lut (.I0(GND_net), .I1(n1797[17]), .I2(GND_net), 
            .I3(n37654), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_20 (.CI(n37654), .I0(n1797[17]), .I1(GND_net), 
            .CO(n37655));
    SB_CARRY add_13_add_1_21902_add_1_25 (.CI(n35909), .I0(n7063[0]), .I1(n58[23]), 
            .CO(n35910));
    SB_LUT4 add_13_add_1_21902_add_1_24_lut (.I0(GND_net), .I1(n282[22]), 
            .I2(n58[22]), .I3(n35908), .O(n57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_19_lut (.I0(GND_net), .I1(n1797[16]), .I2(GND_net), 
            .I3(n37653), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_10_lut (.I0(GND_net), .I1(n16029[7]), .I2(GND_net), 
            .I3(n37568), .O(n15848[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_18 (.CI(n37316), .I0(n8206[15]), .I1(GND_net), .CO(n37317));
    SB_CARRY sub_11_add_2_16 (.CI(n36118), .I0(\PID_CONTROLLER.err_prev[14] ), 
            .I1(n63[14]), .CO(n36119));
    SB_LUT4 add_3246_2_lut (.I0(GND_net), .I1(n29_adj_3505), .I2(n122), 
            .I3(GND_net), .O(n12573[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3246_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_9 (.CI(n37472), .I0(n8391[6]), .I1(GND_net), .CO(n37473));
    SB_LUT4 add_3072_8_lut (.I0(GND_net), .I1(n8391[5]), .I2(n737), .I3(n37471), 
            .O(n8377[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_19 (.CI(n37653), .I0(n1797[16]), .I1(GND_net), 
            .CO(n37654));
    SB_CARRY add_3246_2 (.CI(GND_net), .I0(n29_adj_3505), .I1(n122), .CO(n36335));
    SB_LUT4 sub_11_add_2_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[13] ), 
            .I2(n63[13]), .I3(n36117), .O(n69[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3452_12_lut (.I0(GND_net), .I1(n16418[9]), .I2(GND_net), 
            .I3(n36334), .O(n16312[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3452_11_lut (.I0(GND_net), .I1(n16418[8]), .I2(GND_net), 
            .I3(n36333), .O(n16312[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_8 (.CI(n37471), .I0(n8391[5]), .I1(n737), .CO(n37472));
    SB_LUT4 add_3072_7_lut (.I0(GND_net), .I1(n8391[4]), .I2(n640), .I3(n37470), 
            .O(n8377[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_20 (.CI(n37746), .I0(n1801[17]), .I1(GND_net), 
            .CO(n37747));
    SB_CARRY add_3416_10 (.CI(n37568), .I0(n16029[7]), .I1(GND_net), .CO(n37569));
    SB_LUT4 mult_14_add_1211_18_lut (.I0(GND_net), .I1(n1797[15]), .I2(GND_net), 
            .I3(n37652), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_18 (.CI(n37652), .I0(n1797[15]), .I1(GND_net), 
            .CO(n37653));
    SB_LUT4 mult_14_add_1211_17_lut (.I0(GND_net), .I1(n1797[14]), .I2(GND_net), 
            .I3(n37651), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_20_lut (.I0(GND_net), .I1(n10116[17]), .I2(GND_net), 
            .I3(n37094), .O(n9325[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_15 (.CI(n36117), .I0(\PID_CONTROLLER.err_prev[13] ), 
            .I1(n63[13]), .CO(n36118));
    SB_LUT4 mult_14_add_1215_19_lut (.I0(GND_net), .I1(n1801[16]), .I2(GND_net), 
            .I3(n37745), .O(n1800[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_11 (.CI(n36333), .I0(n16418[8]), .I1(GND_net), .CO(n36334));
    SB_LUT4 add_3452_10_lut (.I0(GND_net), .I1(n16418[7]), .I2(GND_net), 
            .I3(n36332), .O(n16312[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_10 (.CI(n36332), .I0(n16418[7]), .I1(GND_net), .CO(n36333));
    SB_CARRY add_13_add_1_21902_add_1_24 (.CI(n35908), .I0(n282[22]), .I1(n58[22]), 
            .CO(n35909));
    SB_LUT4 sub_11_add_2_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[12] ), 
            .I2(n63[12]), .I3(n36116), .O(n69[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_20 (.CI(n37094), .I0(n10116[17]), .I1(GND_net), 
            .CO(n37095));
    SB_CARRY mult_14_add_1215_19 (.CI(n37745), .I0(n1801[16]), .I1(GND_net), 
            .CO(n37746));
    SB_LUT4 mult_14_add_1215_18_lut (.I0(GND_net), .I1(n1801[15]), .I2(GND_net), 
            .I3(n37744), .O(n1800[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_14 (.CI(n36116), .I0(\PID_CONTROLLER.err_prev[12] ), 
            .I1(n63[12]), .CO(n36117));
    SB_CARRY mult_14_add_1211_17 (.CI(n37651), .I0(n1797[14]), .I1(GND_net), 
            .CO(n37652));
    SB_CARRY mult_14_add_1215_18 (.CI(n37744), .I0(n1801[15]), .I1(GND_net), 
            .CO(n37745));
    SB_LUT4 add_3119_19_lut (.I0(GND_net), .I1(n10116[16]), .I2(GND_net), 
            .I3(n37093), .O(n9325[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n60[6]), 
            .I3(n36016), .O(n67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_16_lut (.I0(GND_net), .I1(n1797[13]), .I2(GND_net), 
            .I3(n37650), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_16 (.CI(n37650), .I0(n1797[13]), .I1(GND_net), 
            .CO(n37651));
    SB_LUT4 add_3062_17_lut (.I0(GND_net), .I1(n8206[14]), .I2(GND_net), 
            .I3(n37315), .O(n8182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3452_9_lut (.I0(GND_net), .I1(n16418[6]), .I2(GND_net), 
            .I3(n36331), .O(n16312[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_17_lut (.I0(GND_net), .I1(n1801[14]), .I2(GND_net), 
            .I3(n37743), .O(n1800[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_7 (.CI(n37470), .I0(n8391[4]), .I1(n640), .CO(n37471));
    SB_LUT4 mult_14_add_1211_15_lut (.I0(GND_net), .I1(n1797[12]), .I2(GND_net), 
            .I3(n37649), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_23_lut (.I0(GND_net), .I1(n282[21]), 
            .I2(n58[21]), .I3(n35907), .O(n57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_8 (.CI(n36016), .I0(GND_net), .I1(n60[6]), 
            .CO(n36017));
    SB_CARRY add_3062_17 (.CI(n37315), .I0(n8206[14]), .I1(GND_net), .CO(n37316));
    SB_CARRY add_3119_19 (.CI(n37093), .I0(n10116[16]), .I1(GND_net), 
            .CO(n37094));
    SB_CARRY mult_14_add_1215_17 (.CI(n37743), .I0(n1801[14]), .I1(GND_net), 
            .CO(n37744));
    SB_LUT4 sub_11_add_2_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[11] ), 
            .I2(n63[11]), .I3(n36115), .O(n69[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3452_9 (.CI(n36331), .I0(n16418[6]), .I1(GND_net), .CO(n36332));
    SB_LUT4 add_3452_8_lut (.I0(GND_net), .I1(n16418[5]), .I2(n740_adj_3511), 
            .I3(n36330), .O(n16312[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i300_2_lut (.I0(\Kd[4] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n446_adj_3512));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i300_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3452_8 (.CI(n36330), .I0(n16418[5]), .I1(n740_adj_3511), 
            .CO(n36331));
    SB_LUT4 mult_14_add_1215_16_lut (.I0(GND_net), .I1(n1801[13]), .I2(GND_net), 
            .I3(n37742), .O(n1800[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_16 (.CI(n37742), .I0(n1801[13]), .I1(GND_net), 
            .CO(n37743));
    SB_LUT4 mult_10_i491_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i491_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_13_add_1_21902_add_1_23 (.CI(n35907), .I0(n282[21]), .I1(n58[21]), 
            .CO(n35908));
    SB_LUT4 mult_14_add_1215_15_lut (.I0(GND_net), .I1(n1801[12]), .I2(GND_net), 
            .I3(n37741), .O(n1800[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3452_7_lut (.I0(GND_net), .I1(n16418[4]), .I2(n643_adj_3513), 
            .I3(n36329), .O(n16312[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_15 (.CI(n37649), .I0(n1797[12]), .I1(GND_net), 
            .CO(n37650));
    SB_LUT4 add_3119_18_lut (.I0(GND_net), .I1(n10116[15]), .I2(GND_net), 
            .I3(n37092), .O(n9325[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_18 (.CI(n37092), .I0(n10116[15]), .I1(GND_net), 
            .CO(n37093));
    SB_CARRY mult_14_add_1215_15 (.CI(n37741), .I0(n1801[12]), .I1(GND_net), 
            .CO(n37742));
    SB_CARRY add_3452_7 (.CI(n36329), .I0(n16418[4]), .I1(n643_adj_3513), 
            .CO(n36330));
    SB_LUT4 add_3452_6_lut (.I0(GND_net), .I1(n16418[3]), .I2(n546_adj_3514), 
            .I3(n36328), .O(n16312[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_17_lut (.I0(GND_net), .I1(n10116[14]), .I2(GND_net), 
            .I3(n37091), .O(n9325[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n60[5]), 
            .I3(n36015), .O(n415)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_14_lut (.I0(GND_net), .I1(n1797[11]), .I2(GND_net), 
            .I3(n37648), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_13 (.CI(n36115), .I0(\PID_CONTROLLER.err_prev[11] ), 
            .I1(n63[11]), .CO(n36116));
    SB_CARRY unary_minus_21_add_3_7 (.CI(n36015), .I0(GND_net), .I1(n60[5]), 
            .CO(n36016));
    SB_CARRY add_3119_17 (.CI(n37091), .I0(n10116[14]), .I1(GND_net), 
            .CO(n37092));
    SB_LUT4 mult_14_add_1215_14_lut (.I0(GND_net), .I1(n1801[11]), .I2(GND_net), 
            .I3(n37740), .O(n1800[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_22_lut (.I0(GND_net), .I1(n282[20]), 
            .I2(n58[20]), .I3(n35906), .O(n57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[10] ), 
            .I2(n63[10]), .I3(n36114), .O(n69[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_22 (.CI(n35906), .I0(n282[20]), .I1(n58[20]), 
            .CO(n35907));
    SB_CARRY add_3452_6 (.CI(n36328), .I0(n16418[3]), .I1(n546_adj_3514), 
            .CO(n36329));
    SB_CARRY mult_14_add_1215_14 (.CI(n37740), .I0(n1801[11]), .I1(GND_net), 
            .CO(n37741));
    SB_LUT4 add_3452_5_lut (.I0(GND_net), .I1(n16418[2]), .I2(n449_adj_3518), 
            .I3(n36327), .O(n16312[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_12 (.CI(n36114), .I0(\PID_CONTROLLER.err_prev[10] ), 
            .I1(n63[10]), .CO(n36115));
    SB_CARRY add_3452_5 (.CI(n36327), .I0(n16418[2]), .I1(n449_adj_3518), 
            .CO(n36328));
    SB_LUT4 mult_14_add_1215_13_lut (.I0(GND_net), .I1(n1801[10]), .I2(GND_net), 
            .I3(n37739), .O(n1800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[9] ), 
            .I2(n63[9]), .I3(n36113), .O(n69[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3452_4_lut (.I0(GND_net), .I1(n16418[1]), .I2(n352_adj_3520), 
            .I3(n36326), .O(n16312[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_11 (.CI(n36113), .I0(\PID_CONTROLLER.err_prev[9] ), 
            .I1(n63[9]), .CO(n36114));
    SB_CARRY add_3452_4 (.CI(n36326), .I0(n16418[1]), .I1(n352_adj_3520), 
            .CO(n36327));
    SB_LUT4 add_3072_6_lut (.I0(GND_net), .I1(n8391[3]), .I2(n543), .I3(n37469), 
            .O(n8377[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n60[4]), 
            .I3(n36014), .O(n67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[8] ), 
            .I2(n63[8]), .I3(n36112), .O(n69[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_16_lut (.I0(GND_net), .I1(n8206[13]), .I2(GND_net), 
            .I3(n37314), .O(n8182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_6 (.CI(n36014), .I0(GND_net), .I1(n60[4]), 
            .CO(n36015));
    SB_LUT4 add_3119_16_lut (.I0(GND_net), .I1(n10116[13]), .I2(GND_net), 
            .I3(n37090), .O(n9325[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n60[3]), 
            .I3(n36013), .O(n67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3452_3_lut (.I0(GND_net), .I1(n16418[0]), .I2(n255_adj_3523), 
            .I3(n36325), .O(n16312[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_16 (.CI(n37314), .I0(n8206[13]), .I1(GND_net), .CO(n37315));
    SB_CARRY add_3452_3 (.CI(n36325), .I0(n16418[0]), .I1(n255_adj_3523), 
            .CO(n36326));
    SB_CARRY add_3119_16 (.CI(n37090), .I0(n10116[13]), .I1(GND_net), 
            .CO(n37091));
    SB_LUT4 add_13_add_1_21902_add_1_21_lut (.I0(GND_net), .I1(n282[19]), 
            .I2(n58[19]), .I3(n35905), .O(n57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_5 (.CI(n36013), .I0(GND_net), .I1(n60[3]), 
            .CO(n36014));
    SB_LUT4 add_3416_9_lut (.I0(GND_net), .I1(n16029[6]), .I2(GND_net), 
            .I3(n37567), .O(n15848[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_10 (.CI(n36112), .I0(\PID_CONTROLLER.err_prev[8] ), 
            .I1(n63[8]), .CO(n36113));
    SB_LUT4 add_3452_2_lut (.I0(GND_net), .I1(n65_adj_3524), .I2(n158_adj_3525), 
            .I3(GND_net), .O(n16312[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3452_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_15_lut (.I0(GND_net), .I1(n10116[12]), .I2(GND_net), 
            .I3(n37089), .O(n9325[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[7] ), 
            .I2(n63[7]), .I3(n36111), .O(n69[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n60[2]), 
            .I3(n36012), .O(n67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_32_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n6540[29]), 
            .I2(GND_net), .I3(n36644), .O(n5784[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3416_9 (.CI(n37567), .I0(n16029[6]), .I1(GND_net), .CO(n37568));
    SB_CARRY add_3452_2 (.CI(GND_net), .I0(n65_adj_3524), .I1(n158_adj_3525), 
            .CO(n36325));
    SB_CARRY unary_minus_21_add_3_4 (.CI(n36012), .I0(GND_net), .I1(n60[2]), 
            .CO(n36013));
    SB_LUT4 mult_10_add_2137_31_lut (.I0(GND_net), .I1(n6540[28]), .I2(GND_net), 
            .I3(n36643), .O(n58[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_31 (.CI(n36643), .I0(n6540[28]), .I1(GND_net), 
            .CO(n36644));
    SB_CARRY add_13_add_1_21902_add_1_21 (.CI(n35905), .I0(n282[19]), .I1(n58[19]), 
            .CO(n35906));
    SB_LUT4 add_3062_15_lut (.I0(GND_net), .I1(n8206[12]), .I2(GND_net), 
            .I3(n37313), .O(n8182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_30_lut (.I0(GND_net), .I1(n6540[27]), .I2(GND_net), 
            .I3(n36642), .O(n58[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_15 (.CI(n37089), .I0(n10116[12]), .I1(GND_net), 
            .CO(n37090));
    SB_LUT4 add_3270_23_lut (.I0(GND_net), .I1(n13592[20]), .I2(GND_net), 
            .I3(n36324), .O(n13107[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_22_lut (.I0(GND_net), .I1(n13592[19]), .I2(GND_net), 
            .I3(n36323), .O(n13107[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_30 (.CI(n36642), .I0(n6540[27]), .I1(GND_net), 
            .CO(n36643));
    SB_CARRY mult_14_add_1215_13 (.CI(n37739), .I0(n1801[10]), .I1(GND_net), 
            .CO(n37740));
    SB_CARRY add_3072_6 (.CI(n37469), .I0(n8391[3]), .I1(n543), .CO(n37470));
    SB_LUT4 add_3119_14_lut (.I0(GND_net), .I1(n10116[11]), .I2(GND_net), 
            .I3(n37088), .O(n9325[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_15 (.CI(n37313), .I0(n8206[12]), .I1(GND_net), .CO(n37314));
    SB_LUT4 mult_10_add_2137_29_lut (.I0(GND_net), .I1(n6540[26]), .I2(GND_net), 
            .I3(n36641), .O(n58[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_29 (.CI(n36641), .I0(n6540[26]), .I1(GND_net), 
            .CO(n36642));
    SB_CARRY add_3270_22 (.CI(n36323), .I0(n13592[19]), .I1(GND_net), 
            .CO(n36324));
    SB_LUT4 add_3270_21_lut (.I0(GND_net), .I1(n13592[18]), .I2(GND_net), 
            .I3(n36322), .O(n13107[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_28_lut (.I0(GND_net), .I1(n6540[25]), .I2(GND_net), 
            .I3(n36640), .O(n58[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_28 (.CI(n36640), .I0(n6540[25]), .I1(GND_net), 
            .CO(n36641));
    SB_CARRY add_3270_21 (.CI(n36322), .I0(n13592[18]), .I1(GND_net), 
            .CO(n36323));
    SB_LUT4 add_3270_20_lut (.I0(GND_net), .I1(n13592[17]), .I2(GND_net), 
            .I3(n36321), .O(n13107[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3270_20 (.CI(n36321), .I0(n13592[17]), .I1(GND_net), 
            .CO(n36322));
    SB_DFF Kd_delay_counter_1013__i0 (.Q(Kd_delay_counter[0]), .C(clk32MHz), 
           .D(n70[0]));   // verilog/motorControl.v(55[27:47])
    SB_LUT4 add_3270_19_lut (.I0(GND_net), .I1(n13592[16]), .I2(GND_net), 
            .I3(n36320), .O(n13107[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_8_lut (.I0(GND_net), .I1(n16029[5]), .I2(n731), .I3(n37566), 
            .O(n15848[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_27_lut (.I0(GND_net), .I1(n6540[24]), .I2(GND_net), 
            .I3(n36639), .O(n58[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_8 (.CI(n37566), .I0(n16029[5]), .I1(n731), .CO(n37567));
    SB_LUT4 add_3072_5_lut (.I0(GND_net), .I1(n8391[2]), .I2(n446_adj_3512), 
            .I3(n37468), .O(n8377[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_14_lut (.I0(GND_net), .I1(n8206[11]), .I2(GND_net), 
            .I3(n37312), .O(n8182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_14 (.CI(n37088), .I0(n10116[11]), .I1(GND_net), 
            .CO(n37089));
    SB_CARRY mult_10_add_2137_27 (.CI(n36639), .I0(n6540[24]), .I1(GND_net), 
            .CO(n36640));
    SB_CARRY add_3270_19 (.CI(n36320), .I0(n13592[16]), .I1(GND_net), 
            .CO(n36321));
    SB_LUT4 mult_10_add_2137_26_lut (.I0(GND_net), .I1(n6540[23]), .I2(GND_net), 
            .I3(n36638), .O(n58[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_26 (.CI(n36638), .I0(n6540[23]), .I1(GND_net), 
            .CO(n36639));
    SB_LUT4 add_3270_18_lut (.I0(GND_net), .I1(n13592[15]), .I2(GND_net), 
            .I3(n36319), .O(n13107[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3270_18 (.CI(n36319), .I0(n13592[15]), .I1(GND_net), 
            .CO(n36320));
    SB_LUT4 mult_10_add_2137_25_lut (.I0(GND_net), .I1(n6540[22]), .I2(GND_net), 
            .I3(n36637), .O(n58[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_9 (.CI(n36111), .I0(\PID_CONTROLLER.err_prev[7] ), 
            .I1(n63[7]), .CO(n36112));
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n60[1]), 
            .I3(n36011), .O(n67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i8_1_lut (.I0(\PID_CONTROLLER.err[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[7]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_2137_25 (.CI(n36637), .I0(n6540[22]), .I1(GND_net), 
            .CO(n36638));
    SB_LUT4 mult_14_add_1215_12_lut (.I0(GND_net), .I1(n1801[9]), .I2(GND_net), 
            .I3(n37738), .O(n1800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_13_lut (.I0(GND_net), .I1(n10116[10]), .I2(GND_net), 
            .I3(n37087), .O(n9325[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_24_lut (.I0(GND_net), .I1(n6540[21]), .I2(GND_net), 
            .I3(n36636), .O(n58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_17_lut (.I0(GND_net), .I1(n13592[14]), .I2(GND_net), 
            .I3(n36318), .O(n13107[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_24 (.CI(n36636), .I0(n6540[21]), .I1(GND_net), 
            .CO(n36637));
    SB_LUT4 mult_10_add_2137_23_lut (.I0(GND_net), .I1(n6540[20]), .I2(GND_net), 
            .I3(n36635), .O(n58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3270_17 (.CI(n36318), .I0(n13592[14]), .I1(GND_net), 
            .CO(n36319));
    SB_LUT4 add_3270_16_lut (.I0(GND_net), .I1(n13592[13]), .I2(GND_net), 
            .I3(n36317), .O(n13107[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_23 (.CI(n36635), .I0(n6540[20]), .I1(GND_net), 
            .CO(n36636));
    SB_LUT4 sub_11_add_2_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[6] ), 
            .I2(n63[6]), .I3(n36110), .O(n69[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_8 (.CI(n36110), .I0(\PID_CONTROLLER.err_prev[6] ), 
            .I1(n63[6]), .CO(n36111));
    SB_CARRY add_3119_13 (.CI(n37087), .I0(n10116[10]), .I1(GND_net), 
            .CO(n37088));
    SB_CARRY add_3072_5 (.CI(n37468), .I0(n8391[2]), .I1(n446_adj_3512), 
            .CO(n37469));
    SB_CARRY unary_minus_21_add_3_3 (.CI(n36011), .I0(GND_net), .I1(n60[1]), 
            .CO(n36012));
    SB_LUT4 mult_10_add_2137_22_lut (.I0(GND_net), .I1(n6540[19]), .I2(GND_net), 
            .I3(n36634), .O(n58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(n28894), .I1(GND_net), .I2(n60[0]), 
            .I3(VCC_net), .O(n46593)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3062_14 (.CI(n37312), .I0(n8206[11]), .I1(GND_net), .CO(n37313));
    SB_LUT4 add_3119_12_lut (.I0(GND_net), .I1(n10116[9]), .I2(GND_net), 
            .I3(n37086), .O(n9325[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_13_lut (.I0(GND_net), .I1(n8206[10]), .I2(GND_net), 
            .I3(n37311), .O(n8182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_22 (.CI(n36634), .I0(n6540[19]), .I1(GND_net), 
            .CO(n36635));
    SB_CARRY add_3119_12 (.CI(n37086), .I0(n10116[9]), .I1(GND_net), .CO(n37087));
    SB_LUT4 mult_10_add_2137_21_lut (.I0(GND_net), .I1(n6540[18]), .I2(GND_net), 
            .I3(n36633), .O(n58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_21 (.CI(n36633), .I0(n6540[18]), .I1(GND_net), 
            .CO(n36634));
    SB_CARRY mult_14_add_1211_14 (.CI(n37648), .I0(n1797[11]), .I1(GND_net), 
            .CO(n37649));
    SB_LUT4 mult_10_i107_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n158_adj_3525));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i107_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3270_16 (.CI(n36317), .I0(n13592[13]), .I1(GND_net), 
            .CO(n36318));
    SB_LUT4 mult_14_add_1211_13_lut (.I0(GND_net), .I1(n1797[10]), .I2(GND_net), 
            .I3(n37647), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_12 (.CI(n37738), .I0(n1801[9]), .I1(GND_net), 
            .CO(n37739));
    SB_LUT4 mult_10_i44_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n65_adj_3524));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_2137_20_lut (.I0(GND_net), .I1(n6540[17]), .I2(GND_net), 
            .I3(n36632), .O(n58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_11_lut (.I0(GND_net), .I1(n1801[8]), .I2(GND_net), 
            .I3(n37737), .O(n1800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_11 (.CI(n37737), .I0(n1801[8]), .I1(GND_net), 
            .CO(n37738));
    SB_LUT4 mult_14_add_1215_10_lut (.I0(GND_net), .I1(n1801[7]), .I2(GND_net), 
            .I3(n37736), .O(n1800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_15_lut (.I0(GND_net), .I1(n13592[12]), .I2(GND_net), 
            .I3(n36316), .O(n13107[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_10 (.CI(n37736), .I0(n1801[7]), .I1(GND_net), 
            .CO(n37737));
    SB_CARRY add_3270_15 (.CI(n36316), .I0(n13592[12]), .I1(GND_net), 
            .CO(n36317));
    SB_CARRY mult_10_add_2137_20 (.CI(n36632), .I0(n6540[17]), .I1(GND_net), 
            .CO(n36633));
    SB_LUT4 sub_11_add_2_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[5] ), 
            .I2(n63[5]), .I3(n36109), .O(n69[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_14_lut (.I0(GND_net), .I1(n13592[11]), .I2(GND_net), 
            .I3(n36315), .O(n13107[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_19_lut (.I0(GND_net), .I1(n6540[16]), .I2(GND_net), 
            .I3(n36631), .O(n58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_13 (.CI(n37311), .I0(n8206[10]), .I1(GND_net), .CO(n37312));
    SB_LUT4 add_3119_11_lut (.I0(GND_net), .I1(n10116[8]), .I2(GND_net), 
            .I3(n37085), .O(n9325[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_7 (.CI(n36109), .I0(\PID_CONTROLLER.err_prev[5] ), 
            .I1(n63[5]), .CO(n36110));
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n60[0]), 
            .CO(n36011));
    SB_LUT4 i22217_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(n69[25]), 
            .I3(GND_net), .O(n10109[0]));   // verilog/motorControl.v(43[26:45])
    defparam i22217_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i22185_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(\Kd[2] ), 
            .I3(GND_net), .O(n35704));   // verilog/motorControl.v(43[26:45])
    defparam i22185_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 add_3022_10_lut (.I0(GND_net), .I1(n1804[22]), .I2(n1711), 
            .I3(n37870), .O(n7063[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3270_14 (.CI(n36315), .I0(n13592[11]), .I1(GND_net), 
            .CO(n36316));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n75[23]), 
            .I3(n36010), .O(n73[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_19 (.CI(n36631), .I0(n6540[16]), .I1(GND_net), 
            .CO(n36632));
    SB_LUT4 add_3270_13_lut (.I0(GND_net), .I1(n13592[10]), .I2(GND_net), 
            .I3(n36314), .O(n13107[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3270_13 (.CI(n36314), .I0(n13592[10]), .I1(GND_net), 
            .CO(n36315));
    SB_LUT4 add_3270_12_lut (.I0(GND_net), .I1(n13592[9]), .I2(GND_net), 
            .I3(n36313), .O(n13107[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3022_9_lut (.I0(GND_net), .I1(n1803[22]), .I2(n1707), 
            .I3(n37869), .O(n7063[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_18_lut (.I0(GND_net), .I1(n6540[15]), .I2(GND_net), 
            .I3(n36630), .O(n58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3022_9 (.CI(n37869), .I0(n1803[22]), .I1(n1707), .CO(n37870));
    SB_LUT4 mult_14_add_1215_9_lut (.I0(GND_net), .I1(n1801[6]), .I2(GND_net), 
            .I3(n37735), .O(n1800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_9 (.CI(n37735), .I0(n1801[6]), .I1(GND_net), 
            .CO(n37736));
    SB_LUT4 mult_14_add_1215_8_lut (.I0(GND_net), .I1(n1801[5]), .I2(n524), 
            .I3(n37734), .O(n1800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3022_8_lut (.I0(GND_net), .I1(n1802[22]), .I2(n1703), 
            .I3(n37868), .O(n7063[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_13 (.CI(n37647), .I0(n1797[10]), .I1(GND_net), 
            .CO(n37648));
    SB_LUT4 sub_11_add_2_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[4] ), 
            .I2(n63[4]), .I3(n36108), .O(n69[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_8 (.CI(n37734), .I0(n1801[5]), .I1(n524), 
            .CO(n37735));
    SB_LUT4 mult_14_add_1215_7_lut (.I0(GND_net), .I1(n1801[4]), .I2(n451), 
            .I3(n37733), .O(n1800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_18 (.CI(n36630), .I0(n6540[15]), .I1(GND_net), 
            .CO(n36631));
    SB_CARRY add_3022_8 (.CI(n37868), .I0(n1802[22]), .I1(n1703), .CO(n37869));
    SB_CARRY mult_14_add_1215_7 (.CI(n37733), .I0(n1801[4]), .I1(n451), 
            .CO(n37734));
    SB_CARRY sub_11_add_2_6 (.CI(n36108), .I0(\PID_CONTROLLER.err_prev[4] ), 
            .I1(n63[4]), .CO(n36109));
    SB_LUT4 mult_14_add_1215_6_lut (.I0(GND_net), .I1(n1801[3]), .I2(n378), 
            .I3(n37732), .O(n1800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3022_7_lut (.I0(GND_net), .I1(n1801[22]), .I2(n1699), 
            .I3(n37867), .O(n7063[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_6 (.CI(n37732), .I0(n1801[3]), .I1(n378), 
            .CO(n37733));
    SB_LUT4 mult_14_add_1211_12_lut (.I0(GND_net), .I1(n1797[9]), .I2(GND_net), 
            .I3(n37646), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_5_lut (.I0(GND_net), .I1(n1801[2]), .I2(n305_adj_3538), 
            .I3(n37731), .O(n1800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3022_7 (.CI(n37867), .I0(n1801[22]), .I1(n1699), .CO(n37868));
    SB_CARRY add_3119_11 (.CI(n37085), .I0(n10116[8]), .I1(GND_net), .CO(n37086));
    SB_LUT4 add_3022_6_lut (.I0(GND_net), .I1(n1800[22]), .I2(n1695), 
            .I3(n37866), .O(n7063[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_17_lut (.I0(GND_net), .I1(n6540[14]), .I2(GND_net), 
            .I3(n36629), .O(n58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_5 (.CI(n37731), .I0(n1801[2]), .I1(n305_adj_3538), 
            .CO(n37732));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[22]), .I3(n36009), .O(n45_adj_3539)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_10_add_2137_17 (.CI(n36629), .I0(n6540[14]), .I1(GND_net), 
            .CO(n36630));
    SB_CARRY add_3022_6 (.CI(n37866), .I0(n1800[22]), .I1(n1695), .CO(n37867));
    SB_CARRY add_3270_12 (.CI(n36313), .I0(n13592[9]), .I1(GND_net), .CO(n36314));
    SB_LUT4 add_3022_5_lut (.I0(GND_net), .I1(n1799[22]), .I2(n1691), 
            .I3(n37865), .O(n7063[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[3] ), 
            .I2(n63[3]), .I3(n36107), .O(n69[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_11_lut (.I0(GND_net), .I1(n13592[8]), .I2(GND_net), 
            .I3(n36312), .O(n13107[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3022_5 (.CI(n37865), .I0(n1799[22]), .I1(n1691), .CO(n37866));
    SB_LUT4 mult_10_add_2137_16_lut (.I0(GND_net), .I1(n6540[13]), .I2(GND_net), 
            .I3(n36628), .O(n58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3022_4_lut (.I0(GND_net), .I1(n1798[22]), .I2(n1687), 
            .I3(n37864), .O(n7063[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_20_lut (.I0(GND_net), .I1(n282[18]), 
            .I2(n58[18]), .I3(n35904), .O(n57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3022_4 (.CI(n37864), .I0(n1798[22]), .I1(n1687), .CO(n37865));
    SB_LUT4 add_3022_3_lut (.I0(GND_net), .I1(n1797[22]), .I2(n1683), 
            .I3(n37863), .O(n7063[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_12 (.CI(n37646), .I0(n1797[9]), .I1(GND_net), 
            .CO(n37647));
    SB_LUT4 mult_10_i172_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n255_adj_3523));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3119_10_lut (.I0(GND_net), .I1(n10116[7]), .I2(GND_net), 
            .I3(n37084), .O(n9325[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i9_1_lut (.I0(\PID_CONTROLLER.err[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[8]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i365_2_lut (.I0(\Kd[5] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n543));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i365_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_13_add_1_21902_add_1_20 (.CI(n35904), .I0(n282[18]), .I1(n58[18]), 
            .CO(n35905));
    SB_CARRY mult_10_add_2137_16 (.CI(n36628), .I0(n6540[13]), .I1(GND_net), 
            .CO(n36629));
    SB_CARRY add_3270_11 (.CI(n36312), .I0(n13592[8]), .I1(GND_net), .CO(n36313));
    SB_CARRY add_3022_3 (.CI(n37863), .I0(n1797[22]), .I1(n1683), .CO(n37864));
    SB_LUT4 mult_14_add_1215_4_lut (.I0(GND_net), .I1(n1801[1]), .I2(n232_adj_3543), 
            .I3(n37730), .O(n1800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut (.I0(n370_adj_3544), .I1(n4_adj_3545), .I2(n35704), 
            .I3(n69[25]), .O(n7_adj_3546));   // verilog/motorControl.v(43[26:45])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6966;
    SB_LUT4 add_3270_10_lut (.I0(GND_net), .I1(n13592[7]), .I2(GND_net), 
            .I3(n36311), .O(n13107[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_19_lut (.I0(GND_net), .I1(n282[17]), 
            .I2(n58[17]), .I3(n35903), .O(n57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n36009), .I0(GND_net), .I1(n75[22]), 
            .CO(n36010));
    SB_CARRY sub_11_add_2_5 (.CI(n36107), .I0(\PID_CONTROLLER.err_prev[3] ), 
            .I1(n63[3]), .CO(n36108));
    SB_CARRY add_3270_10 (.CI(n36311), .I0(n13592[7]), .I1(GND_net), .CO(n36312));
    SB_LUT4 mult_10_add_2137_15_lut (.I0(GND_net), .I1(n6540[12]), .I2(GND_net), 
            .I3(n36627), .O(n58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_10 (.CI(n37084), .I0(n10116[7]), .I1(GND_net), .CO(n37085));
    SB_LUT4 add_3270_9_lut (.I0(GND_net), .I1(n13592[6]), .I2(GND_net), 
            .I3(n36310), .O(n13107[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_15 (.CI(n36627), .I0(n6540[12]), .I1(GND_net), 
            .CO(n36628));
    SB_CARRY add_3270_9 (.CI(n36310), .I0(n13592[6]), .I1(GND_net), .CO(n36311));
    SB_LUT4 mult_10_add_2137_14_lut (.I0(GND_net), .I1(n6540[11]), .I2(GND_net), 
            .I3(n36626), .O(n58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3022_2_lut (.I0(GND_net), .I1(n1796[22]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n7063[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3022_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3022_2 (.CI(GND_net), .I0(n1796[22]), .I1(\PID_CONTROLLER.integral [9]), 
            .CO(n37863));
    SB_LUT4 add_3079_22_lut (.I0(GND_net), .I1(n9325[19]), .I2(GND_net), 
            .I3(n37862), .O(n8470[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_19 (.CI(n35903), .I0(n282[17]), .I1(n58[17]), 
            .CO(n35904));
    SB_LUT4 add_3079_21_lut (.I0(GND_net), .I1(n9325[18]), .I2(GND_net), 
            .I3(n37861), .O(n8470[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i237_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n352_adj_3520));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i237_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3079_21 (.CI(n37861), .I0(n9325[18]), .I1(GND_net), .CO(n37862));
    SB_CARRY mult_14_add_1215_4 (.CI(n37730), .I0(n1801[1]), .I1(n232_adj_3543), 
            .CO(n37731));
    SB_LUT4 mult_14_add_1215_3_lut (.I0(GND_net), .I1(n1801[0]), .I2(n159), 
            .I3(n37729), .O(n1800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_20_lut (.I0(GND_net), .I1(n9325[17]), .I2(GND_net), 
            .I3(n37860), .O(n8470[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_20 (.CI(n37860), .I0(n9325[17]), .I1(GND_net), .CO(n37861));
    SB_LUT4 add_3416_7_lut (.I0(GND_net), .I1(n16029[4]), .I2(n634), .I3(n37565), 
            .O(n15848[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_3 (.CI(n37729), .I0(n1801[0]), .I1(n159), 
            .CO(n37730));
    SB_LUT4 mult_14_add_1211_11_lut (.I0(GND_net), .I1(n1797[8]), .I2(GND_net), 
            .I3(n37645), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_7 (.CI(n37565), .I0(n16029[4]), .I1(n634), .CO(n37566));
    SB_LUT4 add_3072_4_lut (.I0(GND_net), .I1(n8391[1]), .I2(n349), .I3(n37467), 
            .O(n8377[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_12_lut (.I0(GND_net), .I1(n8206[9]), .I2(GND_net), 
            .I3(n37310), .O(n8182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_12 (.CI(n37310), .I0(n8206[9]), .I1(GND_net), .CO(n37311));
    SB_LUT4 add_3119_9_lut (.I0(GND_net), .I1(n10116[6]), .I2(GND_net), 
            .I3(n37083), .O(n9325[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_9 (.CI(n37083), .I0(n10116[6]), .I1(GND_net), .CO(n37084));
    SB_CARRY add_3072_4 (.CI(n37467), .I0(n8391[1]), .I1(n349), .CO(n37468));
    SB_LUT4 add_3079_19_lut (.I0(GND_net), .I1(n9325[16]), .I2(GND_net), 
            .I3(n37859), .O(n8470[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_11_lut (.I0(GND_net), .I1(n8206[8]), .I2(GND_net), 
            .I3(n37309), .O(n8182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_19 (.CI(n37859), .I0(n9325[16]), .I1(GND_net), .CO(n37860));
    SB_LUT4 add_3119_8_lut (.I0(GND_net), .I1(n10116[5]), .I2(n545), .I3(n37082), 
            .O(n9325[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i10_1_lut (.I0(\PID_CONTROLLER.err[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[9]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3119_8 (.CI(n37082), .I0(n10116[5]), .I1(n545), .CO(n37083));
    SB_LUT4 add_3416_6_lut (.I0(GND_net), .I1(n16029[3]), .I2(n537), .I3(n37564), 
            .O(n15848[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_11 (.CI(n37309), .I0(n8206[8]), .I1(GND_net), .CO(n37310));
    SB_LUT4 i1_4_lut_4_lut (.I0(pwm[23]), .I1(hall1), .I2(hall2), .I3(GATES_5__N_3048[5]), 
            .O(n5_adj_3549));   // verilog/motorControl.v(86[38:44])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h55fd;
    SB_LUT4 add_3072_3_lut (.I0(GND_net), .I1(n8391[0]), .I2(n252), .I3(n37466), 
            .O(n8377[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3072_3 (.CI(n37466), .I0(n8391[0]), .I1(n252), .CO(n37467));
    SB_LUT4 add_3062_10_lut (.I0(GND_net), .I1(n8206[7]), .I2(GND_net), 
            .I3(n37308), .O(n8182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_7_lut (.I0(GND_net), .I1(n10116[4]), .I2(n472), .I3(n37081), 
            .O(n9325[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_18_lut (.I0(GND_net), .I1(n9325[15]), .I2(GND_net), 
            .I3(n37858), .O(n8470[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_7 (.CI(n37081), .I0(n10116[4]), .I1(n472), .CO(n37082));
    SB_LUT4 add_3072_2_lut (.I0(GND_net), .I1(n62), .I2(n155), .I3(GND_net), 
            .O(n8377[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3072_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_10 (.CI(n37308), .I0(n8206[7]), .I1(GND_net), .CO(n37309));
    SB_LUT4 add_3119_6_lut (.I0(GND_net), .I1(n10116[3]), .I2(n399_c), 
            .I3(n37080), .O(n9325[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_6 (.CI(n37080), .I0(n10116[3]), .I1(n399_c), .CO(n37081));
    SB_CARRY mult_14_add_1211_11 (.CI(n37645), .I0(n1797[8]), .I1(GND_net), 
            .CO(n37646));
    SB_CARRY add_3072_2 (.CI(GND_net), .I0(n62), .I1(n155), .CO(n37466));
    SB_CARRY add_3416_6 (.CI(n37564), .I0(n16029[3]), .I1(n537), .CO(n37565));
    SB_LUT4 add_3071_14_lut (.I0(GND_net), .I1(n8377[11]), .I2(GND_net), 
            .I3(n37465), .O(n8362[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_5_lut (.I0(GND_net), .I1(n10116[2]), .I2(n326), .I3(n37079), 
            .O(n9325[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_9_lut (.I0(GND_net), .I1(n8206[6]), .I2(GND_net), 
            .I3(n37307), .O(n8182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_5 (.CI(n37079), .I0(n10116[2]), .I1(n326), .CO(n37080));
    SB_LUT4 add_3119_4_lut (.I0(GND_net), .I1(n10116[1]), .I2(n253), .I3(n37078), 
            .O(n9325[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_13_lut (.I0(GND_net), .I1(n8377[10]), .I2(GND_net), 
            .I3(n37464), .O(n8362[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_14 (.CI(n36626), .I0(n6540[11]), .I1(GND_net), 
            .CO(n36627));
    SB_CARRY add_3062_9 (.CI(n37307), .I0(n8206[6]), .I1(GND_net), .CO(n37308));
    SB_LUT4 mult_10_add_2137_13_lut (.I0(GND_net), .I1(n6540[10]), .I2(GND_net), 
            .I3(n36625), .O(n58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_4 (.CI(n37078), .I0(n10116[1]), .I1(n253), .CO(n37079));
    SB_LUT4 add_3062_8_lut (.I0(GND_net), .I1(n8206[5]), .I2(n707), .I3(n37306), 
            .O(n8182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_13 (.CI(n37464), .I0(n8377[10]), .I1(GND_net), .CO(n37465));
    SB_LUT4 add_3119_3_lut (.I0(GND_net), .I1(n10116[0]), .I2(n180), .I3(n37077), 
            .O(n9325[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_8 (.CI(n37306), .I0(n8206[5]), .I1(n707), .CO(n37307));
    SB_LUT4 add_3416_5_lut (.I0(GND_net), .I1(n16029[2]), .I2(n440), .I3(n37563), 
            .O(n15848[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_13 (.CI(n36625), .I0(n6540[10]), .I1(GND_net), 
            .CO(n36626));
    SB_CARRY add_3119_3 (.CI(n37077), .I0(n10116[0]), .I1(n180), .CO(n37078));
    SB_LUT4 add_3071_12_lut (.I0(GND_net), .I1(n8377[9]), .I2(GND_net), 
            .I3(n37463), .O(n8362[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n449_adj_3518));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3062_7_lut (.I0(GND_net), .I1(n8206[4]), .I2(n610), .I3(n37305), 
            .O(n8182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3119_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n9325[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3119_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_12_lut (.I0(GND_net), .I1(n6540[9]), .I2(GND_net), 
            .I3(n36624), .O(n58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_8_lut (.I0(GND_net), .I1(n13592[5]), .I2(n707_adj_3552), 
            .I3(n36309), .O(n13107[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3119_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n37077));
    SB_LUT4 add_3118_7_lut (.I0(GND_net), .I1(n43988), .I2(n658_adj_3553), 
            .I3(n37076), .O(n9317[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3118_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_5 (.CI(n37563), .I0(n16029[2]), .I1(n440), .CO(n37564));
    SB_CARRY add_3071_12 (.CI(n37463), .I0(n8377[9]), .I1(GND_net), .CO(n37464));
    SB_CARRY add_3062_7 (.CI(n37305), .I0(n8206[4]), .I1(n610), .CO(n37306));
    SB_LUT4 add_3118_6_lut (.I0(GND_net), .I1(n10109[3]), .I2(n564), .I3(n37075), 
            .O(n9317[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3118_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_2_lut (.I0(GND_net), .I1(n17_adj_3554), .I2(n86_adj_3555), 
            .I3(GND_net), .O(n1800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_10_lut (.I0(GND_net), .I1(n1797[7]), .I2(GND_net), 
            .I3(n37644), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_4_lut (.I0(GND_net), .I1(n16029[1]), .I2(n343), .I3(n37562), 
            .O(n15848[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_11_lut (.I0(GND_net), .I1(n8377[8]), .I2(GND_net), 
            .I3(n37462), .O(n8362[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_6_lut (.I0(GND_net), .I1(n8206[3]), .I2(n513), .I3(n37304), 
            .O(n8182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_11 (.CI(n37462), .I0(n8377[8]), .I1(GND_net), .CO(n37463));
    SB_CARRY add_3062_6 (.CI(n37304), .I0(n8206[3]), .I1(n513), .CO(n37305));
    SB_CARRY add_3416_4 (.CI(n37562), .I0(n16029[1]), .I1(n343), .CO(n37563));
    SB_LUT4 add_3071_10_lut (.I0(GND_net), .I1(n8377[7]), .I2(GND_net), 
            .I3(n37461), .O(n8362[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_5_lut (.I0(GND_net), .I1(n8206[2]), .I2(n416_adj_3557), 
            .I3(n37303), .O(n8182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_10 (.CI(n37461), .I0(n8377[7]), .I1(GND_net), .CO(n37462));
    SB_CARRY add_3062_5 (.CI(n37303), .I0(n8206[2]), .I1(n416_adj_3557), 
            .CO(n37304));
    SB_CARRY mult_14_add_1211_10 (.CI(n37644), .I0(n1797[7]), .I1(GND_net), 
            .CO(n37645));
    SB_LUT4 add_3416_3_lut (.I0(GND_net), .I1(n16029[0]), .I2(n246_adj_3558), 
            .I3(n37561), .O(n15848[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_2 (.CI(GND_net), .I0(n17_adj_3554), .I1(n86_adj_3555), 
            .CO(n37729));
    SB_CARRY add_3270_8 (.CI(n36309), .I0(n13592[5]), .I1(n707_adj_3552), 
            .CO(n36310));
    SB_CARRY mult_10_add_2137_12 (.CI(n36624), .I0(n6540[9]), .I1(GND_net), 
            .CO(n36625));
    SB_LUT4 add_3071_9_lut (.I0(GND_net), .I1(n8377[6]), .I2(GND_net), 
            .I3(n37460), .O(n8362[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_4_lut (.I0(GND_net), .I1(n8206[1]), .I2(n319), .I3(n37302), 
            .O(n8182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_24_lut (.I0(GND_net), .I1(n1800[21]), .I2(GND_net), 
            .I3(n37727), .O(n1799[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_11_lut (.I0(GND_net), .I1(n6540[8]), .I2(GND_net), 
            .I3(n36623), .O(n58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_9 (.CI(n37460), .I0(n8377[6]), .I1(GND_net), .CO(n37461));
    SB_CARRY add_3062_4 (.CI(n37302), .I0(n8206[1]), .I1(n319), .CO(n37303));
    SB_CARRY add_3079_18 (.CI(n37858), .I0(n9325[15]), .I1(GND_net), .CO(n37859));
    SB_LUT4 add_3270_7_lut (.I0(GND_net), .I1(n13592[4]), .I2(n610_adj_3559), 
            .I3(n36308), .O(n13107[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3416_3 (.CI(n37561), .I0(n16029[0]), .I1(n246_adj_3558), 
            .CO(n37562));
    SB_CARRY add_3270_7 (.CI(n36308), .I0(n13592[4]), .I1(n610_adj_3559), 
            .CO(n36309));
    SB_LUT4 add_3071_8_lut (.I0(GND_net), .I1(n8377[5]), .I2(n734), .I3(n37459), 
            .O(n8362[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_3_lut (.I0(GND_net), .I1(n8206[0]), .I2(n222_adj_3560), 
            .I3(n37301), .O(n8182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i11_1_lut (.I0(\PID_CONTROLLER.err[10] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[10]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3071_8 (.CI(n37459), .I0(n8377[5]), .I1(n734), .CO(n37460));
    SB_CARRY add_3118_6 (.CI(n37075), .I0(n10109[3]), .I1(n564), .CO(n37076));
    SB_LUT4 add_3079_17_lut (.I0(GND_net), .I1(n9325[14]), .I2(GND_net), 
            .I3(n37857), .O(n8470[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_3 (.CI(n37301), .I0(n8206[0]), .I1(n222_adj_3560), 
            .CO(n37302));
    SB_CARRY add_3079_17 (.CI(n37857), .I0(n9325[14]), .I1(GND_net), .CO(n37858));
    SB_CARRY mult_14_add_1214_24 (.CI(n37727), .I0(n1800[21]), .I1(GND_net), 
            .CO(n1695));
    SB_LUT4 mult_14_add_1211_9_lut (.I0(GND_net), .I1(n1797[6]), .I2(GND_net), 
            .I3(n37643), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3416_2_lut (.I0(GND_net), .I1(n56), .I2(n149), .I3(GND_net), 
            .O(n15848[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3416_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_7_lut (.I0(GND_net), .I1(n8377[4]), .I2(n637), .I3(n37458), 
            .O(n8362[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3062_2_lut (.I0(GND_net), .I1(n32_adj_3562), .I2(n125), 
            .I3(GND_net), .O(n8182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3062_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3118_5_lut (.I0(GND_net), .I1(n10844[2]), .I2(n464_adj_3563), 
            .I3(n37074), .O(n9317[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3118_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3062_2 (.CI(GND_net), .I0(n32_adj_3562), .I1(n125), .CO(n37301));
    SB_CARRY add_3118_5 (.CI(n37074), .I0(n10844[2]), .I1(n464_adj_3563), 
            .CO(n37075));
    SB_LUT4 add_3118_4_lut (.I0(GND_net), .I1(n10844[1]), .I2(n370_adj_3544), 
            .I3(n37073), .O(n9317[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3118_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_7 (.CI(n37458), .I0(n8377[4]), .I1(n637), .CO(n37459));
    SB_LUT4 add_3061_24_lut (.I0(GND_net), .I1(n8182[21]), .I2(GND_net), 
            .I3(n37300), .O(n8157[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3118_4 (.CI(n37073), .I0(n10844[1]), .I1(n370_adj_3544), 
            .CO(n37074));
    SB_LUT4 add_3118_3_lut (.I0(GND_net), .I1(n10109[0]), .I2(n276_adj_3564), 
            .I3(n37072), .O(n9317[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3118_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_23_lut (.I0(GND_net), .I1(n1800[20]), .I2(GND_net), 
            .I3(n37726), .O(n1799[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_16_lut (.I0(GND_net), .I1(n9325[13]), .I2(GND_net), 
            .I3(n37856), .O(n8470[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_11 (.CI(n36623), .I0(n6540[8]), .I1(GND_net), 
            .CO(n36624));
    SB_LUT4 add_3061_23_lut (.I0(GND_net), .I1(n8182[20]), .I2(GND_net), 
            .I3(n37299), .O(n8157[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3118_3 (.CI(n37072), .I0(n10109[0]), .I1(n276_adj_3564), 
            .CO(n37073));
    SB_LUT4 mult_10_add_2137_10_lut (.I0(GND_net), .I1(n6540[7]), .I2(GND_net), 
            .I3(n36622), .O(n58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_10 (.CI(n36622), .I0(n6540[7]), .I1(GND_net), 
            .CO(n36623));
    SB_LUT4 add_3118_2_lut (.I0(GND_net), .I1(n86), .I2(n182_adj_3565), 
            .I3(GND_net), .O(n9317[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3118_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3118_2 (.CI(GND_net), .I0(n86), .I1(n182_adj_3565), .CO(n37072));
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n546_adj_3514));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3416_2 (.CI(GND_net), .I0(n56), .I1(n149), .CO(n37561));
    SB_LUT4 add_3071_6_lut (.I0(GND_net), .I1(n8377[3]), .I2(n540), .I3(n37457), 
            .O(n8362[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_23 (.CI(n37299), .I0(n8182[20]), .I1(GND_net), .CO(n37300));
    SB_LUT4 add_3148_20_lut (.I0(GND_net), .I1(n10850[17]), .I2(GND_net), 
            .I3(n37071), .O(n10116[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_19_lut (.I0(GND_net), .I1(n10850[16]), .I2(GND_net), 
            .I3(n37070), .O(n10116[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_22_lut (.I0(GND_net), .I1(n8182[19]), .I2(GND_net), 
            .I3(n37298), .O(n8157[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_19 (.CI(n37070), .I0(n10850[16]), .I1(GND_net), 
            .CO(n37071));
    SB_LUT4 add_3148_18_lut (.I0(GND_net), .I1(n10850[15]), .I2(GND_net), 
            .I3(n37069), .O(n10116[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_6 (.CI(n37457), .I0(n8377[3]), .I1(n540), .CO(n37458));
    SB_CARRY add_3061_22 (.CI(n37298), .I0(n8182[19]), .I1(GND_net), .CO(n37299));
    SB_CARRY add_3148_18 (.CI(n37069), .I0(n10850[15]), .I1(GND_net), 
            .CO(n37070));
    SB_LUT4 add_3148_17_lut (.I0(GND_net), .I1(n10850[14]), .I2(GND_net), 
            .I3(n37068), .O(n10116[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_21_lut (.I0(GND_net), .I1(n8182[18]), .I2(GND_net), 
            .I3(n37297), .O(n8157[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_17 (.CI(n37068), .I0(n10850[14]), .I1(GND_net), 
            .CO(n37069));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[21]), .I3(n36008), .O(n43_adj_3566)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 sub_11_add_2_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[2] ), 
            .I2(n63[2]), .I3(n36106), .O(n69[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_4 (.CI(n36106), .I0(\PID_CONTROLLER.err_prev[2] ), 
            .I1(n63[2]), .CO(n36107));
    SB_LUT4 mult_10_add_2137_9_lut (.I0(GND_net), .I1(n6540[6]), .I2(GND_net), 
            .I3(n36621), .O(n58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_18_lut (.I0(GND_net), .I1(n282[16]), 
            .I2(n58[16]), .I3(n35902), .O(n57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_6_lut (.I0(GND_net), .I1(n13592[3]), .I2(n513_adj_3570), 
            .I3(n36307), .O(n13107[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_16_lut (.I0(GND_net), .I1(n10850[13]), .I2(GND_net), 
            .I3(n37067), .O(n10116[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3270_6 (.CI(n36307), .I0(n13592[3]), .I1(n513_adj_3570), 
            .CO(n36308));
    SB_CARRY mult_10_add_2137_9 (.CI(n36621), .I0(n6540[6]), .I1(GND_net), 
            .CO(n36622));
    SB_LUT4 sub_11_add_2_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[1] ), 
            .I2(n63[1]), .I3(n36105), .O(n69[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_9 (.CI(n37643), .I0(n1797[6]), .I1(GND_net), 
            .CO(n37644));
    SB_LUT4 add_3429_14_lut (.I0(GND_net), .I1(n16183[11]), .I2(GND_net), 
            .I3(n37560), .O(n16029[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_5_lut (.I0(GND_net), .I1(n8377[2]), .I2(n443_adj_3572), 
            .I3(n37456), .O(n8362[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_21 (.CI(n37297), .I0(n8182[18]), .I1(GND_net), .CO(n37298));
    SB_CARRY add_3148_16 (.CI(n37067), .I0(n10850[13]), .I1(GND_net), 
            .CO(n37068));
    SB_LUT4 add_3148_15_lut (.I0(GND_net), .I1(n10850[12]), .I2(GND_net), 
            .I3(n37066), .O(n10116[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_20_lut (.I0(GND_net), .I1(n8182[17]), .I2(GND_net), 
            .I3(n37296), .O(n8157[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_15 (.CI(n37066), .I0(n10850[12]), .I1(GND_net), 
            .CO(n37067));
    SB_LUT4 add_3148_14_lut (.I0(GND_net), .I1(n10850[11]), .I2(GND_net), 
            .I3(n37065), .O(n10116[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_5 (.CI(n37456), .I0(n8377[2]), .I1(n443_adj_3572), 
            .CO(n37457));
    SB_CARRY add_3061_20 (.CI(n37296), .I0(n8182[17]), .I1(GND_net), .CO(n37297));
    SB_LUT4 mult_10_add_2137_8_lut (.I0(GND_net), .I1(n6540[5]), .I2(n680_adj_3574), 
            .I3(n36620), .O(n58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_14 (.CI(n37065), .I0(n10850[11]), .I1(GND_net), 
            .CO(n37066));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n36008), .I0(GND_net), .I1(n75[21]), 
            .CO(n36009));
    SB_LUT4 add_3148_13_lut (.I0(GND_net), .I1(n10850[10]), .I2(GND_net), 
            .I3(n37064), .O(n10116[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_5_lut (.I0(GND_net), .I1(n13592[2]), .I2(n416_adj_3575), 
            .I3(n36306), .O(n13107[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_19_lut (.I0(GND_net), .I1(n8182[16]), .I2(GND_net), 
            .I3(n37295), .O(n8157[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[20]), .I3(n36007), .O(n41_adj_3576)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3270_5 (.CI(n36306), .I0(n13592[2]), .I1(n416_adj_3575), 
            .CO(n36307));
    SB_CARRY add_3148_13 (.CI(n37064), .I0(n10850[10]), .I1(GND_net), 
            .CO(n37065));
    SB_CARRY mult_10_add_2137_8 (.CI(n36620), .I0(n6540[5]), .I1(n680_adj_3574), 
            .CO(n36621));
    SB_LUT4 mult_10_add_2137_7_lut (.I0(GND_net), .I1(n6540[4]), .I2(n583_adj_3579), 
            .I3(n36619), .O(n58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_4_lut (.I0(GND_net), .I1(n13592[1]), .I2(n319_adj_3580), 
            .I3(n36305), .O(n13107[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_12_lut (.I0(GND_net), .I1(n10850[9]), .I2(GND_net), 
            .I3(n37063), .O(n10116[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_7 (.CI(n36619), .I0(n6540[4]), .I1(n583_adj_3579), 
            .CO(n36620));
    SB_CARRY add_3270_4 (.CI(n36305), .I0(n13592[1]), .I1(n319_adj_3580), 
            .CO(n36306));
    SB_LUT4 add_3429_13_lut (.I0(GND_net), .I1(n16183[10]), .I2(GND_net), 
            .I3(n37559), .O(n16029[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3071_4_lut (.I0(GND_net), .I1(n8377[1]), .I2(n346), .I3(n37455), 
            .O(n8362[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_19 (.CI(n37295), .I0(n8182[16]), .I1(GND_net), .CO(n37296));
    SB_CARRY add_3148_12 (.CI(n37063), .I0(n10850[9]), .I1(GND_net), .CO(n37064));
    SB_LUT4 add_3148_11_lut (.I0(GND_net), .I1(n10850[8]), .I2(GND_net), 
            .I3(n37062), .O(n10116[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_18_lut (.I0(GND_net), .I1(n8182[15]), .I2(GND_net), 
            .I3(n37294), .O(n8157[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_11 (.CI(n37062), .I0(n10850[8]), .I1(GND_net), .CO(n37063));
    SB_LUT4 add_3148_10_lut (.I0(GND_net), .I1(n10850[7]), .I2(GND_net), 
            .I3(n37061), .O(n10116[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3071_4 (.CI(n37455), .I0(n8377[1]), .I1(n346), .CO(n37456));
    SB_LUT4 mult_10_add_2137_6_lut (.I0(GND_net), .I1(n6540[3]), .I2(n486_adj_3581), 
            .I3(n36618), .O(n58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_18 (.CI(n37294), .I0(n8182[15]), .I1(GND_net), .CO(n37295));
    SB_CARRY add_3148_10 (.CI(n37061), .I0(n10850[7]), .I1(GND_net), .CO(n37062));
    SB_CARRY sub_11_add_2_3 (.CI(n36105), .I0(\PID_CONTROLLER.err_prev[1] ), 
            .I1(n63[1]), .CO(n36106));
    SB_LUT4 add_3148_9_lut (.I0(GND_net), .I1(n10850[6]), .I2(GND_net), 
            .I3(n37060), .O(n10116[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_17_lut (.I0(GND_net), .I1(n8182[14]), .I2(GND_net), 
            .I3(n37293), .O(n8157[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[0] ), 
            .I2(n63[0]), .I3(VCC_net), .O(n69[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_9 (.CI(n37060), .I0(n10850[6]), .I1(GND_net), .CO(n37061));
    SB_CARRY mult_10_add_2137_6 (.CI(n36618), .I0(n6540[3]), .I1(n486_adj_3581), 
            .CO(n36619));
    SB_LUT4 mult_10_i432_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n643_adj_3513));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i497_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_3511));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i12_1_lut (.I0(\PID_CONTROLLER.err[11] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[11]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n36007), .I0(GND_net), .I1(n75[20]), 
            .CO(n36008));
    SB_LUT4 add_3148_8_lut (.I0(GND_net), .I1(n10850[5]), .I2(n545), .I3(n37059), 
            .O(n10116[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_17 (.CI(n37293), .I0(n8182[14]), .I1(GND_net), .CO(n37294));
    SB_LUT4 mult_10_add_2137_5_lut (.I0(GND_net), .I1(n6540[2]), .I2(n389_adj_3583), 
            .I3(n36617), .O(n58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_23 (.CI(n37726), .I0(n1800[20]), .I1(GND_net), 
            .CO(n37727));
    SB_LUT4 mult_14_add_1211_8_lut (.I0(GND_net), .I1(n1797[5]), .I2(n512), 
            .I3(n37642), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3429_13 (.CI(n37559), .I0(n16183[10]), .I1(GND_net), 
            .CO(n37560));
    SB_LUT4 add_3071_3_lut (.I0(GND_net), .I1(n8377[0]), .I2(n249), .I3(n37454), 
            .O(n8362[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_16_lut (.I0(GND_net), .I1(n8182[13]), .I2(GND_net), 
            .I3(n37292), .O(n8157[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_8 (.CI(n37059), .I0(n10850[5]), .I1(n545), .CO(n37060));
    SB_CARRY add_3061_16 (.CI(n37292), .I0(n8182[13]), .I1(GND_net), .CO(n37293));
    SB_LUT4 add_3148_7_lut (.I0(GND_net), .I1(n10850[4]), .I2(n472), .I3(n37058), 
            .O(n10116[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_5 (.CI(n36617), .I0(n6540[2]), .I1(n389_adj_3583), 
            .CO(n36618));
    SB_LUT4 add_3270_3_lut (.I0(GND_net), .I1(n13592[0]), .I2(n222_adj_3585), 
            .I3(n36304), .O(n13107[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_7 (.CI(n37058), .I0(n10850[4]), .I1(n472), .CO(n37059));
    SB_LUT4 mult_10_add_2137_4_lut (.I0(GND_net), .I1(n6540[1]), .I2(n292_adj_3587), 
            .I3(n36616), .O(n58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3270_3 (.CI(n36304), .I0(n13592[0]), .I1(n222_adj_3585), 
            .CO(n36305));
    SB_LUT4 add_3148_6_lut (.I0(GND_net), .I1(n10850[3]), .I2(n399_c), 
            .I3(n37057), .O(n10116[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3270_2_lut (.I0(GND_net), .I1(n32_adj_3588), .I2(n125_adj_3589), 
            .I3(GND_net), .O(n13107[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3270_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_8 (.CI(n37642), .I0(n1797[5]), .I1(n512), 
            .CO(n37643));
    SB_CARRY mult_10_add_2137_4 (.CI(n36616), .I0(n6540[1]), .I1(n292_adj_3587), 
            .CO(n36617));
    SB_CARRY add_3270_2 (.CI(GND_net), .I0(n32_adj_3588), .I1(n125_adj_3589), 
            .CO(n36304));
    SB_CARRY add_3148_6 (.CI(n37057), .I0(n10850[3]), .I1(n399_c), .CO(n37058));
    SB_CARRY sub_11_add_2_2 (.CI(VCC_net), .I0(\PID_CONTROLLER.err_prev[0] ), 
            .I1(n63[0]), .CO(n36105));
    SB_LUT4 add_3292_22_lut (.I0(GND_net), .I1(n14033[19]), .I2(GND_net), 
            .I3(n36303), .O(n13592[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_21_lut (.I0(GND_net), .I1(n14033[18]), .I2(GND_net), 
            .I3(n36302), .O(n13592[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3429_12_lut (.I0(GND_net), .I1(n16183[9]), .I2(GND_net), 
            .I3(n37558), .O(n16029[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[19]), .I3(n36006), .O(n39_adj_3590)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3071_3 (.CI(n37454), .I0(n8377[0]), .I1(n249), .CO(n37455));
    SB_LUT4 mult_10_add_2137_3_lut (.I0(GND_net), .I1(n6540[0]), .I2(n195_adj_3593), 
            .I3(n36615), .O(n58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(GATES_5__N_3055), 
            .I3(n36104), .O(n853)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n36006), .I0(GND_net), .I1(n75[19]), 
            .CO(n36007));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[18]), .I3(n36005), .O(n37_adj_3594)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3061_15_lut (.I0(GND_net), .I1(n8182[12]), .I2(GND_net), 
            .I3(n37291), .O(n8157[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_15 (.CI(n37291), .I0(n8182[12]), .I1(GND_net), .CO(n37292));
    SB_LUT4 add_3148_5_lut (.I0(GND_net), .I1(n10850[2]), .I2(n326), .I3(n37056), 
            .O(n10116[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_3 (.CI(n36615), .I0(n6540[0]), .I1(n195_adj_3593), 
            .CO(n36616));
    SB_LUT4 mult_10_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3596), .I2(n98_adj_3597), 
            .I3(GND_net), .O(n58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_21 (.CI(n36302), .I0(n14033[18]), .I1(GND_net), 
            .CO(n36303));
    SB_CARRY mult_10_add_2137_2 (.CI(GND_net), .I0(n5_adj_3596), .I1(n98_adj_3597), 
            .CO(n36615));
    SB_LUT4 add_3292_20_lut (.I0(GND_net), .I1(n14033[17]), .I2(GND_net), 
            .I3(n36301), .O(n13592[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_5 (.CI(n37056), .I0(n10850[2]), .I1(n326), .CO(n37057));
    SB_CARRY add_3292_20 (.CI(n36301), .I0(n14033[17]), .I1(GND_net), 
            .CO(n36302));
    SB_LUT4 unary_minus_70_add_3_24_lut (.I0(n852[18]), .I1(GND_net), .I2(n76[22]), 
            .I3(n36103), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY unary_minus_70_add_3_24 (.CI(n36103), .I0(GND_net), .I1(n76[22]), 
            .CO(n36104));
    SB_LUT4 add_3292_19_lut (.I0(GND_net), .I1(n14033[16]), .I2(GND_net), 
            .I3(n36300), .O(n13592[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_19 (.CI(n36300), .I0(n14033[16]), .I1(GND_net), 
            .CO(n36301));
    SB_LUT4 add_3292_18_lut (.I0(GND_net), .I1(n14033[15]), .I2(GND_net), 
            .I3(n36299), .O(n13592[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n76[21]), 
            .I3(n36102), .O(n855)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n36005), .I0(GND_net), .I1(n75[18]), 
            .CO(n36006));
    SB_CARRY add_3292_18 (.CI(n36299), .I0(n14033[15]), .I1(GND_net), 
            .CO(n36300));
    SB_CARRY unary_minus_70_add_3_23 (.CI(n36102), .I0(GND_net), .I1(n76[21]), 
            .CO(n36103));
    SB_LUT4 add_3292_17_lut (.I0(GND_net), .I1(n14033[14]), .I2(GND_net), 
            .I3(n36298), .O(n13592[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3429_12 (.CI(n37558), .I0(n16183[9]), .I1(GND_net), .CO(n37559));
    SB_LUT4 add_3071_2_lut (.I0(GND_net), .I1(n59), .I2(n152_adj_3601), 
            .I3(GND_net), .O(n8362[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_16 (.CI(n37856), .I0(n9325[13]), .I1(GND_net), .CO(n37857));
    SB_LUT4 unary_minus_70_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n76[20]), 
            .I3(n36101), .O(n856)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_14_lut (.I0(GND_net), .I1(n8182[11]), .I2(GND_net), 
            .I3(n37290), .O(n8157[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_14 (.CI(n37290), .I0(n8182[11]), .I1(GND_net), .CO(n37291));
    SB_CARRY add_3292_17 (.CI(n36298), .I0(n14033[14]), .I1(GND_net), 
            .CO(n36299));
    SB_LUT4 add_3148_4_lut (.I0(GND_net), .I1(n10850[1]), .I2(n253), .I3(n37055), 
            .O(n10116[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_16_lut (.I0(GND_net), .I1(n14033[13]), .I2(GND_net), 
            .I3(n36297), .O(n13592[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_4 (.CI(n37055), .I0(n10850[1]), .I1(n253), .CO(n37056));
    SB_CARRY add_3292_16 (.CI(n36297), .I0(n14033[13]), .I1(GND_net), 
            .CO(n36298));
    SB_LUT4 add_3292_15_lut (.I0(GND_net), .I1(n14033[12]), .I2(GND_net), 
            .I3(n36296), .O(n13592[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_22 (.CI(n36101), .I0(GND_net), .I1(n76[20]), 
            .CO(n36102));
    SB_CARRY add_3292_15 (.CI(n36296), .I0(n14033[12]), .I1(GND_net), 
            .CO(n36297));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[17]), .I3(n36004), .O(n35_adj_3603)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3148_3_lut (.I0(GND_net), .I1(n10850[0]), .I2(n180), .I3(n37054), 
            .O(n10116[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_14_lut (.I0(GND_net), .I1(n14033[11]), .I2(GND_net), 
            .I3(n36295), .O(n13592[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n76[19]), 
            .I3(n36100), .O(n857)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_14 (.CI(n36295), .I0(n14033[11]), .I1(GND_net), 
            .CO(n36296));
    SB_LUT4 add_3292_13_lut (.I0(GND_net), .I1(n14033[10]), .I2(GND_net), 
            .I3(n36294), .O(n13592[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_21 (.CI(n36100), .I0(GND_net), .I1(n76[19]), 
            .CO(n36101));
    SB_CARRY add_3292_13 (.CI(n36294), .I0(n14033[10]), .I1(GND_net), 
            .CO(n36295));
    SB_CARRY add_3071_2 (.CI(GND_net), .I0(n59), .I1(n152_adj_3601), .CO(n37454));
    SB_LUT4 add_3061_13_lut (.I0(GND_net), .I1(n8182[10]), .I2(GND_net), 
            .I3(n37289), .O(n8157[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_3 (.CI(n37054), .I0(n10850[0]), .I1(n180), .CO(n37055));
    SB_CARRY add_3061_13 (.CI(n37289), .I0(n8182[10]), .I1(GND_net), .CO(n37290));
    SB_LUT4 add_3148_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n10116[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_12_lut (.I0(GND_net), .I1(n14033[9]), .I2(GND_net), 
            .I3(n36293), .O(n13592[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_12 (.CI(n36293), .I0(n14033[9]), .I1(GND_net), .CO(n36294));
    SB_LUT4 add_2980_31_lut (.I0(GND_net), .I1(n7758[28]), .I2(GND_net), 
            .I3(n36607), .O(n6540[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n76[18]), 
            .I3(n36099), .O(n852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_11_lut (.I0(GND_net), .I1(n14033[8]), .I2(GND_net), 
            .I3(n36292), .O(n13592[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_22_lut (.I0(GND_net), .I1(n1800[19]), .I2(GND_net), 
            .I3(n37725), .O(n1799[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_11 (.CI(n36292), .I0(n14033[8]), .I1(GND_net), .CO(n36293));
    SB_CARRY add_3148_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n37054));
    SB_CARRY unary_minus_5_add_3_19 (.CI(n36004), .I0(GND_net), .I1(n75[17]), 
            .CO(n36005));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[16]), .I3(n36003), .O(n33_adj_3607)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_2980_30_lut (.I0(GND_net), .I1(n7758[27]), .I2(GND_net), 
            .I3(n36606), .O(n6540[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_30 (.CI(n36606), .I0(n7758[27]), .I1(GND_net), .CO(n36607));
    SB_LUT4 add_3292_10_lut (.I0(GND_net), .I1(n14033[7]), .I2(GND_net), 
            .I3(n36291), .O(n13592[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_20 (.CI(n36099), .I0(GND_net), .I1(n76[18]), 
            .CO(n36100));
    SB_CARRY unary_minus_5_add_3_18 (.CI(n36003), .I0(GND_net), .I1(n75[16]), 
            .CO(n36004));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[15]), .I3(n36002), .O(n31_adj_3609)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_70_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n76[17]), 
            .I3(n36098), .O(n859)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_10 (.CI(n36291), .I0(n14033[7]), .I1(GND_net), .CO(n36292));
    SB_LUT4 add_2980_29_lut (.I0(GND_net), .I1(n7758[26]), .I2(GND_net), 
            .I3(n36605), .O(n6540[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_9_lut (.I0(GND_net), .I1(n14033[6]), .I2(GND_net), 
            .I3(n36290), .O(n13592[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_19 (.CI(n36098), .I0(GND_net), .I1(n76[17]), 
            .CO(n36099));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n36002), .I0(GND_net), .I1(n75[15]), 
            .CO(n36003));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[14]), .I3(n36001), .O(n29_adj_3612)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_70_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n76[16]), 
            .I3(n36097), .O(n860)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_9 (.CI(n36290), .I0(n14033[6]), .I1(GND_net), .CO(n36291));
    SB_LUT4 mult_14_add_1211_7_lut (.I0(GND_net), .I1(n1797[4]), .I2(n439), 
            .I3(n37641), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3429_11_lut (.I0(GND_net), .I1(n16183[8]), .I2(GND_net), 
            .I3(n37557), .O(n16029[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_7 (.CI(n37641), .I0(n1797[4]), .I1(n439), 
            .CO(n37642));
    SB_LUT4 add_3176_19_lut (.I0(GND_net), .I1(n11529[16]), .I2(GND_net), 
            .I3(n37053), .O(n10850[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_15_lut (.I0(GND_net), .I1(n8362[12]), .I2(GND_net), 
            .I3(n37453), .O(n8346[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_29 (.CI(n36605), .I0(n7758[26]), .I1(GND_net), .CO(n36606));
    SB_LUT4 add_3061_12_lut (.I0(GND_net), .I1(n8182[9]), .I2(GND_net), 
            .I3(n37288), .O(n8157[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_12 (.CI(n37288), .I0(n8182[9]), .I1(GND_net), .CO(n37289));
    SB_LUT4 add_3176_18_lut (.I0(GND_net), .I1(n11529[15]), .I2(GND_net), 
            .I3(n37052), .O(n10850[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_6_lut (.I0(GND_net), .I1(n1797[3]), .I2(n366), 
            .I3(n37640), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_11_lut (.I0(GND_net), .I1(n8182[8]), .I2(GND_net), 
            .I3(n37287), .O(n8157[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_28_lut (.I0(GND_net), .I1(n7758[25]), .I2(GND_net), 
            .I3(n36604), .O(n6540[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_8_lut (.I0(GND_net), .I1(n14033[5]), .I2(n710_adj_3616), 
            .I3(n36289), .O(n13592[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_28 (.CI(n36604), .I0(n7758[25]), .I1(GND_net), .CO(n36605));
    SB_CARRY add_3292_8 (.CI(n36289), .I0(n14033[5]), .I1(n710_adj_3616), 
            .CO(n36290));
    SB_CARRY add_3176_18 (.CI(n37052), .I0(n11529[15]), .I1(GND_net), 
            .CO(n37053));
    SB_LUT4 add_2980_27_lut (.I0(GND_net), .I1(n7758[24]), .I2(GND_net), 
            .I3(n36603), .O(n6540[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_7_lut (.I0(GND_net), .I1(n14033[4]), .I2(n613_adj_3617), 
            .I3(n36288), .O(n13592[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_18 (.CI(n36097), .I0(GND_net), .I1(n76[16]), 
            .CO(n36098));
    SB_CARRY add_3292_7 (.CI(n36288), .I0(n14033[4]), .I1(n613_adj_3617), 
            .CO(n36289));
    SB_CARRY add_2980_27 (.CI(n36603), .I0(n7758[24]), .I1(GND_net), .CO(n36604));
    SB_LUT4 add_3292_6_lut (.I0(GND_net), .I1(n14033[3]), .I2(n516_adj_3618), 
            .I3(n36287), .O(n13592[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n76[15]), 
            .I3(n36096), .O(n861)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_6 (.CI(n36287), .I0(n14033[3]), .I1(n516_adj_3618), 
            .CO(n36288));
    SB_LUT4 add_3070_14_lut (.I0(GND_net), .I1(n8362[11]), .I2(GND_net), 
            .I3(n37452), .O(n8346[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_11 (.CI(n37287), .I0(n8182[8]), .I1(GND_net), .CO(n37288));
    SB_LUT4 add_3176_17_lut (.I0(GND_net), .I1(n11529[14]), .I2(GND_net), 
            .I3(n37051), .O(n10850[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1014__i0 (.Q(pwm_count[0]), .C(clk32MHz), .D(n64[0]));   // verilog/motorControl.v(110[18:29])
    SB_LUT4 add_3061_10_lut (.I0(GND_net), .I1(n8182[7]), .I2(GND_net), 
            .I3(n37286), .O(n8157[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_17 (.CI(n37051), .I0(n11529[14]), .I1(GND_net), 
            .CO(n37052));
    SB_LUT4 add_2980_26_lut (.I0(GND_net), .I1(n7758[23]), .I2(GND_net), 
            .I3(n36602), .O(n6540[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_26 (.CI(n36602), .I0(n7758[23]), .I1(GND_net), .CO(n36603));
    SB_LUT4 add_3292_5_lut (.I0(GND_net), .I1(n14033[2]), .I2(n419_adj_3620), 
            .I3(n36286), .O(n13592[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_5 (.CI(n36286), .I0(n14033[2]), .I1(n419_adj_3620), 
            .CO(n36287));
    SB_LUT4 add_2980_25_lut (.I0(GND_net), .I1(n7758[22]), .I2(GND_net), 
            .I3(n36601), .O(n6540[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_4_lut (.I0(GND_net), .I1(n14033[1]), .I2(n322_adj_3621), 
            .I3(n36285), .O(n13592[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_16_lut (.I0(GND_net), .I1(n11529[13]), .I2(GND_net), 
            .I3(n37050), .O(n10850[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_25 (.CI(n36601), .I0(n7758[22]), .I1(GND_net), .CO(n36602));
    SB_CARRY add_3292_4 (.CI(n36285), .I0(n14033[1]), .I1(n322_adj_3621), 
            .CO(n36286));
    SB_CARRY unary_minus_70_add_3_17 (.CI(n36096), .I0(GND_net), .I1(n76[15]), 
            .CO(n36097));
    SB_CARRY unary_minus_5_add_3_16 (.CI(n36001), .I0(GND_net), .I1(n75[14]), 
            .CO(n36002));
    SB_LUT4 unary_minus_70_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n76[14]), 
            .I3(n36095), .O(n862)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3292_3_lut (.I0(GND_net), .I1(n14033[0]), .I2(n225_adj_3623), 
            .I3(n36284), .O(n13592[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_24_lut (.I0(GND_net), .I1(n7758[21]), .I2(GND_net), 
            .I3(n36600), .O(n6540[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_3 (.CI(n36284), .I0(n14033[0]), .I1(n225_adj_3623), 
            .CO(n36285));
    SB_LUT4 add_3292_2_lut (.I0(GND_net), .I1(n35_adj_3624), .I2(n128_adj_3625), 
            .I3(GND_net), .O(n13592[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3292_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_16 (.CI(n36095), .I0(GND_net), .I1(n76[14]), 
            .CO(n36096));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[13]), .I3(n36000), .O(n27_adj_3626)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_70_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n76[13]), 
            .I3(n36094), .O(n863)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3292_2 (.CI(GND_net), .I0(n35_adj_3624), .I1(n128_adj_3625), 
            .CO(n36284));
    SB_CARRY add_3429_11 (.CI(n37557), .I0(n16183[8]), .I1(GND_net), .CO(n37558));
    SB_CARRY add_3070_14 (.CI(n37452), .I0(n8362[11]), .I1(GND_net), .CO(n37453));
    SB_CARRY add_3061_10 (.CI(n37286), .I0(n8182[7]), .I1(GND_net), .CO(n37287));
    SB_LUT4 add_3061_9_lut (.I0(GND_net), .I1(n8182[6]), .I2(GND_net), 
            .I3(n37285), .O(n8157[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_16 (.CI(n37050), .I0(n11529[13]), .I1(GND_net), 
            .CO(n37051));
    SB_CARRY unary_minus_70_add_3_15 (.CI(n36094), .I0(GND_net), .I1(n76[13]), 
            .CO(n36095));
    SB_LUT4 add_3176_15_lut (.I0(GND_net), .I1(n11529[12]), .I2(GND_net), 
            .I3(n37049), .O(n10850[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_24 (.CI(n36600), .I0(n7758[21]), .I1(GND_net), .CO(n36601));
    SB_LUT4 add_2980_23_lut (.I0(GND_net), .I1(n7758[20]), .I2(GND_net), 
            .I3(n36599), .O(n6540[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_22 (.CI(n37725), .I0(n1800[19]), .I1(GND_net), 
            .CO(n37726));
    SB_LUT4 add_3462_11_lut (.I0(GND_net), .I1(n16503[8]), .I2(GND_net), 
            .I3(n36283), .O(n16418[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_23 (.CI(n36599), .I0(n7758[20]), .I1(GND_net), .CO(n36600));
    SB_LUT4 add_3462_10_lut (.I0(GND_net), .I1(n16503[7]), .I2(GND_net), 
            .I3(n36282), .O(n16418[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_15 (.CI(n37049), .I0(n11529[12]), .I1(GND_net), 
            .CO(n37050));
    SB_LUT4 add_2980_22_lut (.I0(GND_net), .I1(n7758[19]), .I2(GND_net), 
            .I3(n36598), .O(n6540[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_10 (.CI(n36282), .I0(n16503[7]), .I1(GND_net), .CO(n36283));
    SB_LUT4 mult_12_i304_2_lut (.I0(\Kd[4] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n452_c));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n76[12]), 
            .I3(n36093), .O(n864)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3462_9_lut (.I0(GND_net), .I1(n16503[6]), .I2(GND_net), 
            .I3(n36281), .O(n16418[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_22 (.CI(n36598), .I0(n7758[19]), .I1(GND_net), .CO(n36599));
    SB_CARRY unary_minus_70_add_3_14 (.CI(n36093), .I0(GND_net), .I1(n76[12]), 
            .CO(n36094));
    SB_LUT4 add_2980_21_lut (.I0(GND_net), .I1(n7758[18]), .I2(GND_net), 
            .I3(n36597), .O(n6540[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_9 (.CI(n36281), .I0(n16503[6]), .I1(GND_net), .CO(n36282));
    SB_LUT4 unary_minus_70_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n76[11]), 
            .I3(n36092), .O(n865)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3462_8_lut (.I0(GND_net), .I1(n16503[5]), .I2(n743_adj_3631), 
            .I3(n36280), .O(n16418[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_9 (.CI(n37285), .I0(n8182[6]), .I1(GND_net), .CO(n37286));
    SB_LUT4 mult_14_add_1214_21_lut (.I0(GND_net), .I1(n1800[18]), .I2(GND_net), 
            .I3(n37724), .O(n1799[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_21 (.CI(n36597), .I0(n7758[18]), .I1(GND_net), .CO(n36598));
    SB_LUT4 add_3070_13_lut (.I0(GND_net), .I1(n8362[10]), .I2(GND_net), 
            .I3(n37451), .O(n8346[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_8_lut (.I0(GND_net), .I1(n8182[5]), .I2(n704_adj_3632), 
            .I3(n37284), .O(n8157[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_8 (.CI(n37284), .I0(n8182[5]), .I1(n704_adj_3632), 
            .CO(n37285));
    SB_LUT4 add_3176_14_lut (.I0(GND_net), .I1(n11529[11]), .I2(GND_net), 
            .I3(n37048), .O(n10850[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_6 (.CI(n37640), .I0(n1797[3]), .I1(n366), 
            .CO(n37641));
    SB_LUT4 add_3079_15_lut (.I0(GND_net), .I1(n9325[12]), .I2(GND_net), 
            .I3(n37855), .O(n8470[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_20_lut (.I0(GND_net), .I1(n7758[17]), .I2(GND_net), 
            .I3(n36596), .O(n6540[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_8 (.CI(n36280), .I0(n16503[5]), .I1(n743_adj_3631), 
            .CO(n36281));
    SB_CARRY mult_14_add_1214_21 (.CI(n37724), .I0(n1800[18]), .I1(GND_net), 
            .CO(n37725));
    SB_CARRY add_2980_20 (.CI(n36596), .I0(n7758[17]), .I1(GND_net), .CO(n36597));
    SB_LUT4 add_3462_7_lut (.I0(GND_net), .I1(n16503[4]), .I2(n646_adj_3633), 
            .I3(n36279), .O(n16418[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_14 (.CI(n37048), .I0(n11529[11]), .I1(GND_net), 
            .CO(n37049));
    SB_LUT4 add_2980_19_lut (.I0(GND_net), .I1(n7758[16]), .I2(GND_net), 
            .I3(n36595), .O(n6540[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_7 (.CI(n36279), .I0(n16503[4]), .I1(n646_adj_3633), 
            .CO(n36280));
    SB_CARRY unary_minus_70_add_3_13 (.CI(n36092), .I0(GND_net), .I1(n76[11]), 
            .CO(n36093));
    SB_CARRY unary_minus_5_add_3_15 (.CI(n36000), .I0(GND_net), .I1(n75[13]), 
            .CO(n36001));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[12]), .I3(n35999), .O(n25_adj_3634)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_70_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n76[10]), 
            .I3(n36091), .O(n866)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3462_6_lut (.I0(GND_net), .I1(n16503[3]), .I2(n549_adj_3637), 
            .I3(n36278), .O(n16418[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_15 (.CI(n37855), .I0(n9325[12]), .I1(GND_net), .CO(n37856));
    SB_LUT4 add_3079_14_lut (.I0(GND_net), .I1(n9325[11]), .I2(GND_net), 
            .I3(n37854), .O(n8470[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_14 (.CI(n37854), .I0(n9325[11]), .I1(GND_net), .CO(n37855));
    SB_LUT4 add_3079_13_lut (.I0(GND_net), .I1(n9325[10]), .I2(GND_net), 
            .I3(n37853), .O(n8470[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_13 (.CI(n37853), .I0(n9325[10]), .I1(GND_net), .CO(n37854));
    SB_LUT4 mult_14_add_1214_20_lut (.I0(GND_net), .I1(n1800[17]), .I2(GND_net), 
            .I3(n37723), .O(n1799[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_12_lut (.I0(GND_net), .I1(n9325[9]), .I2(GND_net), 
            .I3(n37852), .O(n8470[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n35999), .I0(GND_net), .I1(n75[12]), 
            .CO(n36000));
    SB_CARRY add_3070_13 (.CI(n37451), .I0(n8362[10]), .I1(GND_net), .CO(n37452));
    SB_LUT4 add_3070_12_lut (.I0(GND_net), .I1(n8362[9]), .I2(GND_net), 
            .I3(n37450), .O(n8346[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3429_10_lut (.I0(GND_net), .I1(n16183[7]), .I2(GND_net), 
            .I3(n37556), .O(n16029[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_20 (.CI(n37723), .I0(n1800[17]), .I1(GND_net), 
            .CO(n37724));
    SB_CARRY add_2980_19 (.CI(n36595), .I0(n7758[16]), .I1(GND_net), .CO(n36596));
    SB_LUT4 sub_11_inv_0_i13_1_lut (.I0(\PID_CONTROLLER.err[12] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[12]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3079_12 (.CI(n37852), .I0(n9325[9]), .I1(GND_net), .CO(n37853));
    SB_LUT4 add_3079_11_lut (.I0(GND_net), .I1(n9325[8]), .I2(GND_net), 
            .I3(n37851), .O(n8470[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_19_lut (.I0(GND_net), .I1(n1800[16]), .I2(GND_net), 
            .I3(n37722), .O(n1799[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_7_lut (.I0(GND_net), .I1(n8182[4]), .I2(n607_adj_3638), 
            .I3(n37283), .O(n8157[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_19 (.CI(n37722), .I0(n1800[16]), .I1(GND_net), 
            .CO(n37723));
    SB_LUT4 mult_14_add_1211_5_lut (.I0(GND_net), .I1(n1797[2]), .I2(n293), 
            .I3(n37639), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3429_10 (.CI(n37556), .I0(n16183[7]), .I1(GND_net), .CO(n37557));
    SB_LUT4 add_2980_18_lut (.I0(GND_net), .I1(n7758[15]), .I2(GND_net), 
            .I3(n36594), .O(n6540[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_18 (.CI(n36594), .I0(n7758[15]), .I1(GND_net), .CO(n36595));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[11]), .I3(n35998), .O(n23_adj_3640)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3070_12 (.CI(n37450), .I0(n8362[9]), .I1(GND_net), .CO(n37451));
    SB_CARRY add_3061_7 (.CI(n37283), .I0(n8182[4]), .I1(n607_adj_3638), 
            .CO(n37284));
    SB_LUT4 add_3176_13_lut (.I0(GND_net), .I1(n11529[10]), .I2(GND_net), 
            .I3(n37047), .O(n10850[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_13 (.CI(n37047), .I0(n11529[10]), .I1(GND_net), 
            .CO(n37048));
    SB_LUT4 add_3061_6_lut (.I0(GND_net), .I1(n8182[3]), .I2(n510_adj_3642), 
            .I3(n37282), .O(n8157[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_12_lut (.I0(GND_net), .I1(n11529[9]), .I2(GND_net), 
            .I3(n37046), .O(n10850[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_6 (.CI(n37282), .I0(n8182[3]), .I1(n510_adj_3642), 
            .CO(n37283));
    SB_CARRY add_3176_12 (.CI(n37046), .I0(n11529[9]), .I1(GND_net), .CO(n37047));
    SB_LUT4 add_3176_11_lut (.I0(GND_net), .I1(n11529[8]), .I2(GND_net), 
            .I3(n37045), .O(n10850[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n35998), .I0(GND_net), .I1(n75[11]), 
            .CO(n35999));
    SB_CARRY add_3176_11 (.CI(n37045), .I0(n11529[8]), .I1(GND_net), .CO(n37046));
    SB_LUT4 add_3429_9_lut (.I0(GND_net), .I1(n16183[6]), .I2(GND_net), 
            .I3(n37555), .O(n16029[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_11_lut (.I0(GND_net), .I1(n8362[8]), .I2(GND_net), 
            .I3(n37449), .O(n8346[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3462_6 (.CI(n36278), .I0(n16503[3]), .I1(n549_adj_3637), 
            .CO(n36279));
    SB_LUT4 add_3061_5_lut (.I0(GND_net), .I1(n8182[2]), .I2(n413_adj_3643), 
            .I3(n37281), .O(n8157[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3462_5_lut (.I0(GND_net), .I1(n16503[2]), .I2(n452_adj_3644), 
            .I3(n36277), .O(n16418[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_10_lut (.I0(GND_net), .I1(n11529[7]), .I2(GND_net), 
            .I3(n37044), .O(n10850[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_17_lut (.I0(GND_net), .I1(n7758[14]), .I2(GND_net), 
            .I3(n36593), .O(n6540[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_10 (.CI(n37044), .I0(n11529[7]), .I1(GND_net), .CO(n37045));
    SB_CARRY mult_14_add_1211_5 (.CI(n37639), .I0(n1797[2]), .I1(n293), 
            .CO(n37640));
    SB_CARRY add_3061_5 (.CI(n37281), .I0(n8182[2]), .I1(n413_adj_3643), 
            .CO(n37282));
    SB_CARRY add_3429_9 (.CI(n37555), .I0(n16183[6]), .I1(GND_net), .CO(n37556));
    SB_CARRY add_3070_11 (.CI(n37449), .I0(n8362[8]), .I1(GND_net), .CO(n37450));
    SB_LUT4 add_3061_4_lut (.I0(GND_net), .I1(n8182[1]), .I2(n316_adj_3645), 
            .I3(n37280), .O(n8157[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_9_lut (.I0(GND_net), .I1(n11529[6]), .I2(GND_net), 
            .I3(n37043), .O(n10850[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_17 (.CI(n36593), .I0(n7758[14]), .I1(GND_net), .CO(n36594));
    SB_CARRY add_3462_5 (.CI(n36277), .I0(n16503[2]), .I1(n452_adj_3644), 
            .CO(n36278));
    SB_LUT4 add_3462_4_lut (.I0(GND_net), .I1(n16503[1]), .I2(n355_adj_3646), 
            .I3(n36276), .O(n16418[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_16_lut (.I0(GND_net), .I1(n7758[13]), .I2(GND_net), 
            .I3(n36592), .O(n6540[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_16 (.CI(n36592), .I0(n7758[13]), .I1(GND_net), .CO(n36593));
    SB_CARRY add_3462_4 (.CI(n36276), .I0(n16503[1]), .I1(n355_adj_3646), 
            .CO(n36277));
    SB_LUT4 add_3462_3_lut (.I0(GND_net), .I1(n16503[0]), .I2(n258_adj_3647), 
            .I3(n36275), .O(n16418[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_15_lut (.I0(GND_net), .I1(n7758[12]), .I2(GND_net), 
            .I3(n36591), .O(n6540[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_9 (.CI(n37043), .I0(n11529[6]), .I1(GND_net), .CO(n37044));
    SB_CARRY add_2980_15 (.CI(n36591), .I0(n7758[12]), .I1(GND_net), .CO(n36592));
    SB_CARRY add_3462_3 (.CI(n36275), .I0(n16503[0]), .I1(n258_adj_3647), 
            .CO(n36276));
    SB_LUT4 add_3462_2_lut (.I0(GND_net), .I1(n68_adj_3648), .I2(n161_adj_3649), 
            .I3(GND_net), .O(n16418[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3462_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_14_lut (.I0(GND_net), .I1(n7758[11]), .I2(GND_net), 
            .I3(n36590), .O(n6540[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_14 (.CI(n36590), .I0(n7758[11]), .I1(GND_net), .CO(n36591));
    SB_CARRY add_3462_2 (.CI(GND_net), .I0(n68_adj_3648), .I1(n161_adj_3649), 
            .CO(n36275));
    SB_LUT4 add_3313_21_lut (.I0(GND_net), .I1(n14432[18]), .I2(GND_net), 
            .I3(n36274), .O(n14033[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_13_lut (.I0(GND_net), .I1(n7758[10]), .I2(GND_net), 
            .I3(n36589), .O(n6540[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_4 (.CI(n37280), .I0(n8182[1]), .I1(n316_adj_3645), 
            .CO(n37281));
    SB_LUT4 add_3176_8_lut (.I0(GND_net), .I1(n11529[5]), .I2(n545), .I3(n37042), 
            .O(n10850[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_13 (.CI(n36589), .I0(n7758[10]), .I1(GND_net), .CO(n36590));
    SB_CARRY add_3176_8 (.CI(n37042), .I0(n11529[5]), .I1(n545), .CO(n37043));
    SB_LUT4 add_3313_20_lut (.I0(GND_net), .I1(n14432[17]), .I2(GND_net), 
            .I3(n36273), .O(n14033[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_7_lut (.I0(GND_net), .I1(n11529[4]), .I2(n472), .I3(n37041), 
            .O(n10850[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_4_lut (.I0(GND_net), .I1(n1797[1]), .I2(n220_adj_3651), 
            .I3(n37638), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3429_8_lut (.I0(GND_net), .I1(n16183[5]), .I2(n734_adj_3652), 
            .I3(n37554), .O(n16029[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_18 (.CI(n35902), .I0(n282[16]), .I1(n58[16]), 
            .CO(n35903));
    SB_CARRY unary_minus_70_add_3_12 (.CI(n36091), .I0(GND_net), .I1(n76[10]), 
            .CO(n36092));
    SB_LUT4 mult_14_add_1214_18_lut (.I0(GND_net), .I1(n1800[15]), .I2(GND_net), 
            .I3(n37721), .O(n1799[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_18 (.CI(n37721), .I0(n1800[15]), .I1(GND_net), 
            .CO(n37722));
    SB_CARRY add_3079_11 (.CI(n37851), .I0(n9325[8]), .I1(GND_net), .CO(n37852));
    SB_LUT4 mult_14_add_1214_17_lut (.I0(GND_net), .I1(n1800[14]), .I2(GND_net), 
            .I3(n37720), .O(n1799[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_10_lut (.I0(GND_net), .I1(n9325[7]), .I2(GND_net), 
            .I3(n37850), .O(n8470[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_4 (.CI(n37638), .I0(n1797[1]), .I1(n220_adj_3651), 
            .CO(n37639));
    SB_CARRY mult_14_add_1214_17 (.CI(n37720), .I0(n1800[14]), .I1(GND_net), 
            .CO(n37721));
    SB_CARRY add_3313_20 (.CI(n36273), .I0(n14432[17]), .I1(GND_net), 
            .CO(n36274));
    SB_LUT4 mult_14_add_1211_3_lut (.I0(GND_net), .I1(n1797[0]), .I2(n147_adj_3653), 
            .I3(n37637), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_16_lut (.I0(GND_net), .I1(n1800[13]), .I2(GND_net), 
            .I3(n37719), .O(n1799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[21]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[16]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[17]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2980_12_lut (.I0(GND_net), .I1(n7758[9]), .I2(GND_net), 
            .I3(n36588), .O(n6540[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_10 (.CI(n37850), .I0(n9325[7]), .I1(GND_net), .CO(n37851));
    SB_CARRY add_2980_12 (.CI(n36588), .I0(n7758[9]), .I1(GND_net), .CO(n36589));
    SB_LUT4 add_3313_19_lut (.I0(GND_net), .I1(n14432[16]), .I2(GND_net), 
            .I3(n36272), .O(n14033[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_3 (.CI(n37637), .I0(n1797[0]), .I1(n147_adj_3653), 
            .CO(n37638));
    SB_CARRY add_3313_19 (.CI(n36272), .I0(n14432[16]), .I1(GND_net), 
            .CO(n36273));
    SB_LUT4 add_2980_11_lut (.I0(GND_net), .I1(n7758[8]), .I2(GND_net), 
            .I3(n36587), .O(n6540[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_7 (.CI(n37041), .I0(n11529[4]), .I1(n472), .CO(n37042));
    SB_LUT4 add_3079_9_lut (.I0(GND_net), .I1(n9325[6]), .I2(GND_net), 
            .I3(n37849), .O(n8470[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_16 (.CI(n37719), .I0(n1800[13]), .I1(GND_net), 
            .CO(n37720));
    SB_LUT4 mult_14_add_1214_15_lut (.I0(GND_net), .I1(n1800[12]), .I2(GND_net), 
            .I3(n37718), .O(n1799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_11 (.CI(n36587), .I0(n7758[8]), .I1(GND_net), .CO(n36588));
    SB_LUT4 add_3313_18_lut (.I0(GND_net), .I1(n14432[15]), .I2(GND_net), 
            .I3(n36271), .O(n14033[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_18 (.CI(n36271), .I0(n14432[15]), .I1(GND_net), 
            .CO(n36272));
    SB_LUT4 add_2980_10_lut (.I0(GND_net), .I1(n7758[7]), .I2(GND_net), 
            .I3(n36586), .O(n6540[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_10 (.CI(n36586), .I0(n7758[7]), .I1(GND_net), .CO(n36587));
    SB_LUT4 add_3313_17_lut (.I0(GND_net), .I1(n14432[14]), .I2(GND_net), 
            .I3(n36270), .O(n14033[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_17 (.CI(n36270), .I0(n14432[14]), .I1(GND_net), 
            .CO(n36271));
    SB_LUT4 add_2980_9_lut (.I0(GND_net), .I1(n7758[6]), .I2(GND_net), 
            .I3(n36585), .O(n6540[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_15 (.CI(n37718), .I0(n1800[12]), .I1(GND_net), 
            .CO(n37719));
    SB_LUT4 add_3070_10_lut (.I0(GND_net), .I1(n8362[7]), .I2(GND_net), 
            .I3(n37448), .O(n8346[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3313_16_lut (.I0(GND_net), .I1(n14432[13]), .I2(GND_net), 
            .I3(n36269), .O(n14033[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_3_lut (.I0(GND_net), .I1(n8182[0]), .I2(n219_adj_3654), 
            .I3(n37279), .O(n8157[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_6_lut (.I0(GND_net), .I1(n11529[3]), .I2(n399_c), 
            .I3(n37040), .O(n10850[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_10 (.CI(n37448), .I0(n8362[7]), .I1(GND_net), .CO(n37449));
    SB_CARRY add_3061_3 (.CI(n37279), .I0(n8182[0]), .I1(n219_adj_3654), 
            .CO(n37280));
    SB_CARRY add_3176_6 (.CI(n37040), .I0(n11529[3]), .I1(n399_c), .CO(n37041));
    SB_LUT4 add_3176_5_lut (.I0(GND_net), .I1(n11529[2]), .I2(n326), .I3(n37039), 
            .O(n10850[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_9 (.CI(n36585), .I0(n7758[6]), .I1(GND_net), .CO(n36586));
    SB_CARRY add_3313_16 (.CI(n36269), .I0(n14432[13]), .I1(GND_net), 
            .CO(n36270));
    SB_LUT4 add_3313_15_lut (.I0(GND_net), .I1(n14432[12]), .I2(GND_net), 
            .I3(n36268), .O(n14033[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_8_lut (.I0(GND_net), .I1(n7758[5]), .I2(n683_adj_3655), 
            .I3(n36584), .O(n6540[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i369_2_lut (.I0(\Kd[5] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n549));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_14_lut (.I0(GND_net), .I1(n1800[11]), .I2(GND_net), 
            .I3(n37717), .O(n1799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i430_2_lut (.I0(\Kd[6] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n640));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i430_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3079_9 (.CI(n37849), .I0(n9325[6]), .I1(GND_net), .CO(n37850));
    SB_CARRY add_2980_8 (.CI(n36584), .I0(n7758[5]), .I1(n683_adj_3655), 
            .CO(n36585));
    SB_CARRY add_3313_15 (.CI(n36268), .I0(n14432[12]), .I1(GND_net), 
            .CO(n36269));
    SB_LUT4 add_3313_14_lut (.I0(GND_net), .I1(n14432[11]), .I2(GND_net), 
            .I3(n36267), .O(n14033[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_7_lut (.I0(GND_net), .I1(n7758[4]), .I2(n586_adj_3656), 
            .I3(n36583), .O(n6540[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_5 (.CI(n37039), .I0(n11529[2]), .I1(n326), .CO(n37040));
    SB_CARRY add_2980_7 (.CI(n36583), .I0(n7758[4]), .I1(n586_adj_3656), 
            .CO(n36584));
    SB_CARRY add_3313_14 (.CI(n36267), .I0(n14432[11]), .I1(GND_net), 
            .CO(n36268));
    SB_LUT4 add_3313_13_lut (.I0(GND_net), .I1(n14432[10]), .I2(GND_net), 
            .I3(n36266), .O(n14033[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_6_lut (.I0(GND_net), .I1(n7758[3]), .I2(n489_adj_3657), 
            .I3(n36582), .O(n6540[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_6 (.CI(n36582), .I0(n7758[3]), .I1(n489_adj_3657), 
            .CO(n36583));
    SB_LUT4 mult_10_i164_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n243));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i164_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3313_13 (.CI(n36266), .I0(n14432[10]), .I1(GND_net), 
            .CO(n36267));
    SB_LUT4 add_3313_12_lut (.I0(GND_net), .I1(n14432[9]), .I2(GND_net), 
            .I3(n36265), .O(n14033[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_5_lut (.I0(GND_net), .I1(n7758[2]), .I2(n392_adj_3658), 
            .I3(n36581), .O(n6540[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3061_2_lut (.I0(GND_net), .I1(n29_adj_3659), .I2(n122_adj_3660), 
            .I3(GND_net), .O(n8157[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3061_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3176_4_lut (.I0(GND_net), .I1(n11529[1]), .I2(n253), .I3(n37038), 
            .O(n10850[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3061_2 (.CI(GND_net), .I0(n29_adj_3659), .I1(n122_adj_3660), 
            .CO(n37279));
    SB_CARRY add_3176_4 (.CI(n37038), .I0(n11529[1]), .I1(n253), .CO(n37039));
    SB_CARRY add_2980_5 (.CI(n36581), .I0(n7758[2]), .I1(n392_adj_3658), 
            .CO(n36582));
    SB_CARRY add_3313_12 (.CI(n36265), .I0(n14432[9]), .I1(GND_net), .CO(n36266));
    SB_LUT4 add_3313_11_lut (.I0(GND_net), .I1(n14432[8]), .I2(GND_net), 
            .I3(n36264), .O(n14033[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_4_lut (.I0(GND_net), .I1(n7758[1]), .I2(n295_adj_3661), 
            .I3(n36580), .O(n6540[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_4 (.CI(n36580), .I0(n7758[1]), .I1(n295_adj_3661), 
            .CO(n36581));
    SB_CARRY add_3313_11 (.CI(n36264), .I0(n14432[8]), .I1(GND_net), .CO(n36265));
    SB_LUT4 add_3313_10_lut (.I0(GND_net), .I1(n14432[7]), .I2(GND_net), 
            .I3(n36263), .O(n14033[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_3_lut (.I0(GND_net), .I1(n7758[0]), .I2(n198_adj_3662), 
            .I3(n36579), .O(n6540[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[18]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3176_3_lut (.I0(GND_net), .I1(n11529[0]), .I2(n180), .I3(n37037), 
            .O(n10850[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_3 (.CI(n36579), .I0(n7758[0]), .I1(n198_adj_3662), 
            .CO(n36580));
    SB_CARRY add_3313_10 (.CI(n36263), .I0(n14432[7]), .I1(GND_net), .CO(n36264));
    SB_LUT4 add_3313_9_lut (.I0(GND_net), .I1(n14432[6]), .I2(GND_net), 
            .I3(n36262), .O(n14033[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2980_2_lut (.I0(GND_net), .I1(n8_adj_3663), .I2(n101_adj_3664), 
            .I3(GND_net), .O(n6540[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2980_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2980_2 (.CI(GND_net), .I0(n8_adj_3663), .I1(n101_adj_3664), 
            .CO(n36579));
    SB_LUT4 add_3047_30_lut (.I0(GND_net), .I1(n9123[27]), .I2(GND_net), 
            .I3(n36578), .O(n7758[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_9 (.CI(n36262), .I0(n14432[6]), .I1(GND_net), .CO(n36263));
    SB_LUT4 add_3313_8_lut (.I0(GND_net), .I1(n14432[5]), .I2(n713_adj_3665), 
            .I3(n36261), .O(n14033[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_29_lut (.I0(GND_net), .I1(n9123[26]), .I2(GND_net), 
            .I3(n36577), .O(n7758[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_8 (.CI(n36261), .I0(n14432[5]), .I1(n713_adj_3665), 
            .CO(n36262));
    SB_CARRY add_3429_8 (.CI(n37554), .I0(n16183[5]), .I1(n734_adj_3652), 
            .CO(n37555));
    SB_LUT4 add_3070_9_lut (.I0(GND_net), .I1(n8362[6]), .I2(GND_net), 
            .I3(n37447), .O(n8346[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_25_lut (.I0(GND_net), .I1(n8157[22]), .I2(GND_net), 
            .I3(n37278), .O(n8131[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3176_3 (.CI(n37037), .I0(n11529[0]), .I1(n180), .CO(n37038));
    SB_LUT4 unary_minus_70_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n76[9]), 
            .I3(n36090), .O(n867)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_29 (.CI(n36577), .I0(n9123[26]), .I1(GND_net), .CO(n36578));
    SB_LUT4 add_3176_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n10850[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3176_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3313_7_lut (.I0(GND_net), .I1(n14432[4]), .I2(n616_adj_3667), 
            .I3(n36260), .O(n14033[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_7 (.CI(n36260), .I0(n14432[4]), .I1(n616_adj_3667), 
            .CO(n36261));
    SB_LUT4 add_3313_6_lut (.I0(GND_net), .I1(n14432[3]), .I2(n519_adj_3668), 
            .I3(n36259), .O(n14033[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_28_lut (.I0(GND_net), .I1(n9123[25]), .I2(GND_net), 
            .I3(n36576), .O(n7758[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_28 (.CI(n36576), .I0(n9123[25]), .I1(GND_net), .CO(n36577));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[10]), .I3(n35997), .O(n21_adj_3669)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3313_6 (.CI(n36259), .I0(n14432[3]), .I1(n519_adj_3668), 
            .CO(n36260));
    SB_CARRY unary_minus_70_add_3_11 (.CI(n36090), .I0(GND_net), .I1(n76[9]), 
            .CO(n36091));
    SB_LUT4 unary_minus_21_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[22]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3047_27_lut (.I0(GND_net), .I1(n9123[24]), .I2(GND_net), 
            .I3(n36575), .O(n7758[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[19]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3176_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n37037));
    SB_LUT4 add_3429_7_lut (.I0(GND_net), .I1(n16183[4]), .I2(n637_adj_3671), 
            .I3(n37553), .O(n16029[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3203_18_lut (.I0(GND_net), .I1(n12155[15]), .I2(GND_net), 
            .I3(n37036), .O(n11529[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_9 (.CI(n37447), .I0(n8362[6]), .I1(GND_net), .CO(n37448));
    SB_LUT4 add_13_add_1_21902_add_1_17_lut (.I0(GND_net), .I1(n282[15]), 
            .I2(n58[15]), .I3(n35901), .O(n57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3429_7 (.CI(n37553), .I0(n16183[4]), .I1(n637_adj_3671), 
            .CO(n37554));
    SB_LUT4 add_13_add_1_21902_add_1_31_lut (.I0(GND_net), .I1(n7063[6]), 
            .I2(n58[29]), .I3(n35915), .O(n57[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_24_lut (.I0(GND_net), .I1(n8157[21]), .I2(GND_net), 
            .I3(n37277), .O(n8131[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i14_1_lut (.I0(\PID_CONTROLLER.err[13] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[13]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_14_add_1214_14 (.CI(n37717), .I0(n1800[11]), .I1(GND_net), 
            .CO(n37718));
    SB_LUT4 add_3079_8_lut (.I0(GND_net), .I1(n9325[5]), .I2(n545), .I3(n37848), 
            .O(n8470[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_32 (.CI(n35916), .I0(n7063[7]), .I1(n58[30]), 
            .CO(n35917));
    SB_CARRY add_13_add_1_21902_add_1_17 (.CI(n35901), .I0(n282[15]), .I1(n58[15]), 
            .CO(n35902));
    SB_LUT4 mult_14_add_1214_13_lut (.I0(GND_net), .I1(n1800[10]), .I2(GND_net), 
            .I3(n37716), .O(n1799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_8 (.CI(n37848), .I0(n9325[5]), .I1(n545), .CO(n37849));
    SB_CARRY mult_14_add_1214_13 (.CI(n37716), .I0(n1800[10]), .I1(GND_net), 
            .CO(n37717));
    SB_LUT4 add_3079_7_lut (.I0(GND_net), .I1(n9325[4]), .I2(n472), .I3(n37847), 
            .O(n8470[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3313_5_lut (.I0(GND_net), .I1(n14432[2]), .I2(n422_adj_3672), 
            .I3(n36258), .O(n14033[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_27 (.CI(n36575), .I0(n9123[24]), .I1(GND_net), .CO(n36576));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n35997), .I0(GND_net), .I1(n75[10]), 
            .CO(n35998));
    SB_LUT4 add_3047_26_lut (.I0(GND_net), .I1(n9123[23]), .I2(GND_net), 
            .I3(n36574), .O(n7758[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_7 (.CI(n37847), .I0(n9325[4]), .I1(n472), .CO(n37848));
    SB_CARRY add_3047_26 (.CI(n36574), .I0(n9123[23]), .I1(GND_net), .CO(n36575));
    SB_LUT4 mult_14_add_1211_2_lut (.I0(GND_net), .I1(n5_adj_3673), .I2(n74_adj_3674), 
            .I3(GND_net), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n76[8]), 
            .I3(n36089), .O(n868)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_12_lut (.I0(GND_net), .I1(n1800[9]), .I2(GND_net), 
            .I3(n37715), .O(n1799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_8_lut (.I0(GND_net), .I1(n8362[5]), .I2(n731_adj_3676), 
            .I3(n37446), .O(n8346[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3203_17_lut (.I0(GND_net), .I1(n12155[14]), .I2(GND_net), 
            .I3(n37035), .O(n11529[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_32_lut (.I0(GND_net), .I1(n7063[7]), 
            .I2(n58[30]), .I3(n35916), .O(n57[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_6_lut (.I0(GND_net), .I1(n9325[3]), .I2(n399_c), 
            .I3(n37846), .O(n8470[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_6 (.CI(n37846), .I0(n9325[3]), .I1(n399_c), .CO(n37847));
    SB_CARRY add_3060_24 (.CI(n37277), .I0(n8157[21]), .I1(GND_net), .CO(n37278));
    SB_LUT4 add_13_add_1_21902_add_1_16_lut (.I0(GND_net), .I1(n282[14]), 
            .I2(n58[14]), .I3(n35900), .O(n57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[20]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_14_add_1211_2 (.CI(GND_net), .I0(n5_adj_3673), .I1(n74_adj_3674), 
            .CO(n37637));
    SB_LUT4 add_3429_6_lut (.I0(GND_net), .I1(n16183[3]), .I2(n540_adj_3677), 
            .I3(n37552), .O(n16029[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_25_lut (.I0(GND_net), .I1(n9123[22]), .I2(GND_net), 
            .I3(n36573), .O(n7758[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_5 (.CI(n36258), .I0(n14432[2]), .I1(n422_adj_3672), 
            .CO(n36259));
    SB_LUT4 add_3313_4_lut (.I0(GND_net), .I1(n14432[1]), .I2(n325_adj_3678), 
            .I3(n36257), .O(n14033[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_25 (.CI(n36573), .I0(n9123[22]), .I1(GND_net), .CO(n36574));
    SB_LUT4 add_3047_24_lut (.I0(GND_net), .I1(n9123[21]), .I2(GND_net), 
            .I3(n36572), .O(n7758[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_4 (.CI(n36257), .I0(n14432[1]), .I1(n325_adj_3678), 
            .CO(n36258));
    SB_LUT4 add_3313_3_lut (.I0(GND_net), .I1(n14432[0]), .I2(n228_adj_3679), 
            .I3(n36256), .O(n14033[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_24 (.CI(n36572), .I0(n9123[21]), .I1(GND_net), .CO(n36573));
    SB_LUT4 add_3060_23_lut (.I0(GND_net), .I1(n8157[20]), .I2(GND_net), 
            .I3(n37276), .O(n8131[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_17 (.CI(n37035), .I0(n12155[14]), .I1(GND_net), 
            .CO(n37036));
    SB_LUT4 add_3047_23_lut (.I0(GND_net), .I1(n9123[20]), .I2(GND_net), 
            .I3(n36571), .O(n7758[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_3 (.CI(n36256), .I0(n14432[0]), .I1(n228_adj_3679), 
            .CO(n36257));
    SB_LUT4 add_3313_2_lut (.I0(GND_net), .I1(n38_adj_3680), .I2(n131_adj_3681), 
            .I3(GND_net), .O(n14033[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3313_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_23 (.CI(n36571), .I0(n9123[20]), .I1(GND_net), .CO(n36572));
    SB_CARRY mult_14_add_1214_12 (.CI(n37715), .I0(n1800[9]), .I1(GND_net), 
            .CO(n37716));
    SB_LUT4 add_3047_22_lut (.I0(GND_net), .I1(n9123[19]), .I2(GND_net), 
            .I3(n36570), .O(n7758[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3313_2 (.CI(GND_net), .I0(n38_adj_3680), .I1(n131_adj_3681), 
            .CO(n36256));
    SB_LUT4 add_3333_20_lut (.I0(GND_net), .I1(n14791[17]), .I2(GND_net), 
            .I3(n36255), .O(n14432[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_22 (.CI(n36570), .I0(n9123[19]), .I1(GND_net), .CO(n36571));
    SB_LUT4 add_3203_16_lut (.I0(GND_net), .I1(n12155[13]), .I2(GND_net), 
            .I3(n37034), .O(n11529[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_10 (.CI(n36089), .I0(GND_net), .I1(n76[8]), 
            .CO(n36090));
    SB_CARRY add_3070_8 (.CI(n37446), .I0(n8362[5]), .I1(n731_adj_3676), 
            .CO(n37447));
    SB_LUT4 add_13_add_1_21902_add_1_33_lut (.I0(GND_net), .I1(n7063[8]), 
            .I2(n5784[0]), .I3(n35917), .O(n57[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_16 (.CI(n35900), .I0(n282[14]), .I1(n58[14]), 
            .CO(n35901));
    SB_CARRY add_3060_23 (.CI(n37276), .I0(n8157[20]), .I1(GND_net), .CO(n37277));
    SB_LUT4 add_3060_22_lut (.I0(GND_net), .I1(n8157[19]), .I2(GND_net), 
            .I3(n37275), .O(n8131[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_15_lut (.I0(GND_net), .I1(n282[13]), 
            .I2(n58[13]), .I3(n35899), .O(n57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_16 (.CI(n37034), .I0(n12155[13]), .I1(GND_net), 
            .CO(n37035));
    SB_LUT4 add_3079_5_lut (.I0(GND_net), .I1(n9325[2]), .I2(n326), .I3(n37845), 
            .O(n8470[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3203_15_lut (.I0(GND_net), .I1(n12155[12]), .I2(GND_net), 
            .I3(n37033), .O(n11529[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_21_lut (.I0(GND_net), .I1(n9123[18]), .I2(GND_net), 
            .I3(n36569), .O(n7758[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_15 (.CI(n37033), .I0(n12155[12]), .I1(GND_net), 
            .CO(n37034));
    SB_CARRY add_3047_21 (.CI(n36569), .I0(n9123[18]), .I1(GND_net), .CO(n36570));
    SB_LUT4 add_3333_19_lut (.I0(GND_net), .I1(n14791[16]), .I2(GND_net), 
            .I3(n36254), .O(n14432[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_19 (.CI(n36254), .I0(n14791[16]), .I1(GND_net), 
            .CO(n36255));
    SB_LUT4 add_3047_20_lut (.I0(GND_net), .I1(n9123[17]), .I2(GND_net), 
            .I3(n36568), .O(n7758[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_20 (.CI(n36568), .I0(n9123[17]), .I1(GND_net), .CO(n36569));
    SB_LUT4 add_3333_18_lut (.I0(GND_net), .I1(n14791[15]), .I2(GND_net), 
            .I3(n36253), .O(n14432[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_18 (.CI(n36253), .I0(n14791[15]), .I1(GND_net), 
            .CO(n36254));
    SB_LUT4 add_3047_19_lut (.I0(GND_net), .I1(n9123[16]), .I2(GND_net), 
            .I3(n36567), .O(n7758[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_7_lut (.I0(GND_net), .I1(n8362[4]), .I2(n634_adj_3682), 
            .I3(n37445), .O(n8346[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_22 (.CI(n37275), .I0(n8157[19]), .I1(GND_net), .CO(n37276));
    SB_LUT4 add_3203_14_lut (.I0(GND_net), .I1(n12155[11]), .I2(GND_net), 
            .I3(n37032), .O(n11529[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_19 (.CI(n36567), .I0(n9123[16]), .I1(GND_net), .CO(n36568));
    SB_LUT4 add_3333_17_lut (.I0(GND_net), .I1(n14791[14]), .I2(GND_net), 
            .I3(n36252), .O(n14432[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_18_lut (.I0(GND_net), .I1(n9123[15]), .I2(GND_net), 
            .I3(n36566), .O(n7758[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_17 (.CI(n36252), .I0(n14791[14]), .I1(GND_net), 
            .CO(n36253));
    SB_CARRY add_3047_18 (.CI(n36566), .I0(n9123[15]), .I1(GND_net), .CO(n36567));
    SB_LUT4 add_3047_17_lut (.I0(GND_net), .I1(n9123[14]), .I2(GND_net), 
            .I3(n36565), .O(n7758[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_16_lut (.I0(GND_net), .I1(n14791[13]), .I2(GND_net), 
            .I3(n36251), .O(n14432[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_16 (.CI(n36251), .I0(n14791[13]), .I1(GND_net), 
            .CO(n36252));
    SB_CARRY add_3047_17 (.CI(n36565), .I0(n9123[14]), .I1(GND_net), .CO(n36566));
    SB_CARRY add_3203_14 (.CI(n37032), .I0(n12155[11]), .I1(GND_net), 
            .CO(n37033));
    SB_LUT4 add_3047_16_lut (.I0(GND_net), .I1(n9123[13]), .I2(GND_net), 
            .I3(n36564), .O(n7758[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3203_13_lut (.I0(GND_net), .I1(n12155[10]), .I2(GND_net), 
            .I3(n37031), .O(n11529[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i434_2_lut (.I0(\Kd[6] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n646));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n75[9]), .I3(n35996), .O(n19_adj_3683)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3079_5 (.CI(n37845), .I0(n9325[2]), .I1(n326), .CO(n37846));
    SB_LUT4 unary_minus_70_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n76[7]), 
            .I3(n36088), .O(n869)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_21_lut (.I0(GND_net), .I1(n8157[18]), .I2(GND_net), 
            .I3(n37274), .O(n8131[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_13 (.CI(n37031), .I0(n12155[10]), .I1(GND_net), 
            .CO(n37032));
    SB_LUT4 mult_14_add_1214_11_lut (.I0(GND_net), .I1(n1800[8]), .I2(GND_net), 
            .I3(n37714), .O(n1799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_18_lut (.I0(GND_net), .I1(n15397[15]), .I2(GND_net), 
            .I3(n37636), .O(n15112[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3429_6 (.CI(n37552), .I0(n16183[3]), .I1(n540_adj_3677), 
            .CO(n37553));
    SB_CARRY add_3070_7 (.CI(n37445), .I0(n8362[4]), .I1(n634_adj_3682), 
            .CO(n37446));
    SB_CARRY add_3060_21 (.CI(n37274), .I0(n8157[18]), .I1(GND_net), .CO(n37275));
    SB_LUT4 add_3060_20_lut (.I0(GND_net), .I1(n8157[17]), .I2(GND_net), 
            .I3(n37273), .O(n8131[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3429_5_lut (.I0(GND_net), .I1(n16183[2]), .I2(n443_adj_3686), 
            .I3(n37551), .O(n16029[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_6_lut (.I0(GND_net), .I1(n8362[3]), .I2(n537_adj_3687), 
            .I3(n37444), .O(n8346[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_20 (.CI(n37273), .I0(n8157[17]), .I1(GND_net), .CO(n37274));
    SB_LUT4 add_3060_19_lut (.I0(GND_net), .I1(n8157[16]), .I2(GND_net), 
            .I3(n37272), .O(n8131[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_17_lut (.I0(GND_net), .I1(n15397[14]), .I2(GND_net), 
            .I3(n37635), .O(n15112[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_15_lut (.I0(GND_net), .I1(n14791[12]), .I2(GND_net), 
            .I3(n36250), .O(n14432[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_15 (.CI(n36250), .I0(n14791[12]), .I1(GND_net), 
            .CO(n36251));
    SB_CARRY add_3047_16 (.CI(n36564), .I0(n9123[13]), .I1(GND_net), .CO(n36565));
    SB_LUT4 add_3047_15_lut (.I0(GND_net), .I1(n9123[12]), .I2(GND_net), 
            .I3(n36563), .O(n7758[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_14_lut (.I0(GND_net), .I1(n14791[11]), .I2(GND_net), 
            .I3(n36249), .O(n14432[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i229_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n340));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[21]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3333_14 (.CI(n36249), .I0(n14791[11]), .I1(GND_net), 
            .CO(n36250));
    SB_CARRY add_3047_15 (.CI(n36563), .I0(n9123[12]), .I1(GND_net), .CO(n36564));
    SB_CARRY add_3060_19 (.CI(n37272), .I0(n8157[16]), .I1(GND_net), .CO(n37273));
    SB_LUT4 unary_minus_21_inv_0_i32_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[31]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3203_12_lut (.I0(GND_net), .I1(n12155[9]), .I2(GND_net), 
            .I3(n37030), .O(n11529[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[22]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3047_14_lut (.I0(GND_net), .I1(n9123[11]), .I2(GND_net), 
            .I3(n36562), .O(n7758[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i499_2_lut (.I0(\Kd[7] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3079_4_lut (.I0(GND_net), .I1(n9325[1]), .I2(n253), .I3(n37844), 
            .O(n8470[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3429_5 (.CI(n37551), .I0(n16183[2]), .I1(n443_adj_3686), 
            .CO(n37552));
    SB_CARRY add_3070_6 (.CI(n37444), .I0(n8362[3]), .I1(n537_adj_3687), 
            .CO(n37445));
    SB_LUT4 add_3060_18_lut (.I0(GND_net), .I1(n8157[15]), .I2(GND_net), 
            .I3(n37271), .O(n8131[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_18 (.CI(n37271), .I0(n8157[15]), .I1(GND_net), .CO(n37272));
    SB_LUT4 add_3429_4_lut (.I0(GND_net), .I1(n16183[1]), .I2(n346_adj_3688), 
            .I3(n37550), .O(n16029[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_5_lut (.I0(GND_net), .I1(n8362[2]), .I2(n440_adj_3689), 
            .I3(n37443), .O(n8346[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_13_lut (.I0(GND_net), .I1(n14791[10]), .I2(GND_net), 
            .I3(n36248), .O(n14432[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_13 (.CI(n36248), .I0(n14791[10]), .I1(GND_net), 
            .CO(n36249));
    SB_CARRY add_3047_14 (.CI(n36562), .I0(n9123[11]), .I1(GND_net), .CO(n36563));
    SB_LUT4 add_3047_13_lut (.I0(GND_net), .I1(n9123[10]), .I2(GND_net), 
            .I3(n36561), .O(n7758[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_12_lut (.I0(GND_net), .I1(n14791[9]), .I2(GND_net), 
            .I3(n36247), .O(n14432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[23]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[0]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3410));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3333_12 (.CI(n36247), .I0(n14791[9]), .I1(GND_net), .CO(n36248));
    SB_CARRY add_3047_13 (.CI(n36561), .I0(n9123[10]), .I1(GND_net), .CO(n36562));
    SB_LUT4 mult_10_i144_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n213));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i144_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3203_12 (.CI(n37030), .I0(n12155[9]), .I1(GND_net), .CO(n37031));
    SB_LUT4 mult_12_i73_2_lut (.I0(\Kd[1] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_3409));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i10_2_lut (.I0(\Kd[0] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i209_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n310));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i91_2_lut (.I0(\Kd[1] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n134));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3047_12_lut (.I0(GND_net), .I1(n9123[9]), .I2(GND_net), 
            .I3(n36560), .O(n7758[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_11_lut (.I0(GND_net), .I1(n14791[8]), .I2(GND_net), 
            .I3(n36246), .O(n14432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i28_2_lut (.I0(\Kd[0] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_c));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i138_2_lut (.I0(\Kd[2] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i138_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3070_5 (.CI(n37443), .I0(n8362[2]), .I1(n440_adj_3689), 
            .CO(n37444));
    SB_LUT4 add_3060_17_lut (.I0(GND_net), .I1(n8157[14]), .I2(GND_net), 
            .I3(n37270), .O(n8131[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_17 (.CI(n37270), .I0(n8157[14]), .I1(GND_net), .CO(n37271));
    SB_CARRY add_3079_4 (.CI(n37844), .I0(n9325[1]), .I1(n253), .CO(n37845));
    SB_CARRY mult_14_add_1214_11 (.CI(n37714), .I0(n1800[8]), .I1(GND_net), 
            .CO(n37715));
    SB_CARRY add_3370_17 (.CI(n37635), .I0(n15397[14]), .I1(GND_net), 
            .CO(n37636));
    SB_CARRY add_3429_4 (.CI(n37550), .I0(n16183[1]), .I1(n346_adj_3688), 
            .CO(n37551));
    SB_LUT4 mult_12_i156_2_lut (.I0(\Kd[2] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n231));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3070_4_lut (.I0(GND_net), .I1(n8362[1]), .I2(n343_adj_3690), 
            .I3(n37442), .O(n8346[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_16_lut (.I0(GND_net), .I1(n8157[13]), .I2(GND_net), 
            .I3(n37269), .O(n8131[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n35996), .I0(GND_net), .I1(n75[9]), 
            .CO(n35997));
    SB_CARRY add_3060_16 (.CI(n37269), .I0(n8157[13]), .I1(GND_net), .CO(n37270));
    SB_CARRY add_3047_12 (.CI(n36560), .I0(n9123[9]), .I1(GND_net), .CO(n36561));
    SB_LUT4 mult_10_i294_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n437));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3203_11_lut (.I0(GND_net), .I1(n12155[8]), .I2(GND_net), 
            .I3(n37029), .O(n11529[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_11_lut (.I0(GND_net), .I1(n9123[8]), .I2(GND_net), 
            .I3(n36559), .O(n7758[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_15_lut (.I0(GND_net), .I1(n8157[12]), .I2(GND_net), 
            .I3(n37268), .O(n8131[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_11 (.CI(n37029), .I0(n12155[8]), .I1(GND_net), .CO(n37030));
    SB_LUT4 add_3203_10_lut (.I0(GND_net), .I1(n12155[7]), .I2(GND_net), 
            .I3(n37028), .O(n11529[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_10 (.CI(n37028), .I0(n12155[7]), .I1(GND_net), .CO(n37029));
    SB_CARRY add_3060_15 (.CI(n37268), .I0(n8157[12]), .I1(GND_net), .CO(n37269));
    SB_CARRY add_3070_4 (.CI(n37442), .I0(n8362[1]), .I1(n343_adj_3690), 
            .CO(n37443));
    SB_LUT4 mult_14_add_1214_10_lut (.I0(GND_net), .I1(n1800[7]), .I2(GND_net), 
            .I3(n37713), .O(n1799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_14_lut (.I0(GND_net), .I1(n8157[11]), .I2(GND_net), 
            .I3(n37267), .O(n8131[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_3_lut (.I0(GND_net), .I1(n8362[0]), .I2(n246_adj_3691), 
            .I3(n37441), .O(n8346[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3203_9_lut (.I0(GND_net), .I1(n12155[6]), .I2(GND_net), 
            .I3(n37027), .O(n11529[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_9 (.CI(n36088), .I0(GND_net), .I1(n76[7]), 
            .CO(n36089));
    SB_CARRY add_3333_11 (.CI(n36246), .I0(n14791[8]), .I1(GND_net), .CO(n36247));
    SB_CARRY add_3203_9 (.CI(n37027), .I0(n12155[6]), .I1(GND_net), .CO(n37028));
    SB_LUT4 add_3333_10_lut (.I0(GND_net), .I1(n14791[7]), .I2(GND_net), 
            .I3(n36245), .O(n14432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3429_3_lut (.I0(GND_net), .I1(n16183[0]), .I2(n249_adj_3692), 
            .I3(n37549), .O(n16029[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_14 (.CI(n37267), .I0(n8157[11]), .I1(GND_net), .CO(n37268));
    SB_CARRY add_3429_3 (.CI(n37549), .I0(n16183[0]), .I1(n249_adj_3692), 
            .CO(n37550));
    SB_LUT4 add_3203_8_lut (.I0(GND_net), .I1(n12155[5]), .I2(n545), .I3(n37026), 
            .O(n11529[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_16_lut (.I0(GND_net), .I1(n15397[13]), .I2(GND_net), 
            .I3(n37634), .O(n15112[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3203_8 (.CI(n37026), .I0(n12155[5]), .I1(n545), .CO(n37027));
    SB_LUT4 add_3429_2_lut (.I0(GND_net), .I1(n59_adj_3693), .I2(n152_adj_3694), 
            .I3(GND_net), .O(n16029[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3429_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3429_2 (.CI(GND_net), .I0(n59_adj_3693), .I1(n152_adj_3694), 
            .CO(n37549));
    SB_CARRY add_3047_11 (.CI(n36559), .I0(n9123[8]), .I1(GND_net), .CO(n36560));
    SB_CARRY add_13_add_1_21902_add_1_15 (.CI(n35899), .I0(n282[13]), .I1(n58[13]), 
            .CO(n35900));
    SB_LUT4 add_3441_13_lut (.I0(GND_net), .I1(n16312[10]), .I2(GND_net), 
            .I3(n37548), .O(n16183[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_3 (.CI(n37441), .I0(n8362[0]), .I1(n246_adj_3691), 
            .CO(n37442));
    SB_LUT4 add_13_add_1_21902_add_1_14_lut (.I0(GND_net), .I1(n282[12]), 
            .I2(n58[12]), .I3(n35898), .O(n57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_13_lut (.I0(GND_net), .I1(n8157[10]), .I2(GND_net), 
            .I3(n37266), .O(n8131[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3203_7_lut (.I0(GND_net), .I1(n12155[4]), .I2(n472), .I3(n37025), 
            .O(n11529[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_12_lut (.I0(GND_net), .I1(n16312[9]), .I2(GND_net), 
            .I3(n37547), .O(n16183[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_16 (.CI(n37634), .I0(n15397[13]), .I1(GND_net), 
            .CO(n37635));
    SB_CARRY add_3203_7 (.CI(n37025), .I0(n12155[4]), .I1(n472), .CO(n37026));
    SB_LUT4 mult_12_i203_2_lut (.I0(\Kd[3] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n301));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i268_2_lut (.I0(\Kd[4] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n398));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i268_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3060_13 (.CI(n37266), .I0(n8157[10]), .I1(GND_net), .CO(n37267));
    SB_CARRY mult_14_add_1214_10 (.CI(n37713), .I0(n1800[7]), .I1(GND_net), 
            .CO(n37714));
    SB_LUT4 add_3203_6_lut (.I0(GND_net), .I1(n12155[3]), .I2(n399_c), 
            .I3(n37024), .O(n11529[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n76[6]), 
            .I3(n36087), .O(n870)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_6 (.CI(n37024), .I0(n12155[3]), .I1(n399_c), .CO(n37025));
    SB_LUT4 add_3203_5_lut (.I0(GND_net), .I1(n12155[2]), .I2(n326), .I3(n37023), 
            .O(n11529[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3070_2_lut (.I0(GND_net), .I1(n56_adj_3696), .I2(n149_adj_3697), 
            .I3(GND_net), .O(n8346[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3070_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_12_lut (.I0(GND_net), .I1(n8157[9]), .I2(GND_net), 
            .I3(n37265), .O(n8131[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n75[8]), .I3(n35995), .O(n17_adj_3698)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3047_10_lut (.I0(GND_net), .I1(n9123[7]), .I2(GND_net), 
            .I3(n36558), .O(n7758[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3079_3_lut (.I0(GND_net), .I1(n9325[0]), .I2(n180), .I3(n37843), 
            .O(n8470[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_5 (.CI(n37023), .I0(n12155[2]), .I1(n326), .CO(n37024));
    SB_LUT4 add_3370_15_lut (.I0(GND_net), .I1(n15397[12]), .I2(GND_net), 
            .I3(n37633), .O(n15112[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_10 (.CI(n36245), .I0(n14791[7]), .I1(GND_net), .CO(n36246));
    SB_LUT4 add_3203_4_lut (.I0(GND_net), .I1(n12155[1]), .I2(n253), .I3(n37022), 
            .O(n11529[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_12 (.CI(n37265), .I0(n8157[9]), .I1(GND_net), .CO(n37266));
    SB_CARRY add_3203_4 (.CI(n37022), .I0(n12155[1]), .I1(n253), .CO(n37023));
    SB_CARRY add_13_add_1_21902_add_1_14 (.CI(n35898), .I0(n282[12]), .I1(n58[12]), 
            .CO(n35899));
    SB_LUT4 add_3203_3_lut (.I0(GND_net), .I1(n12155[0]), .I2(n180), .I3(n37021), 
            .O(n11529[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_12 (.CI(n37547), .I0(n16312[9]), .I1(GND_net), .CO(n37548));
    SB_CARRY add_3047_10 (.CI(n36558), .I0(n9123[7]), .I1(GND_net), .CO(n36559));
    SB_LUT4 add_3047_9_lut (.I0(GND_net), .I1(n9123[6]), .I2(GND_net), 
            .I3(n36557), .O(n7758[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_15 (.CI(n37633), .I0(n15397[12]), .I1(GND_net), 
            .CO(n37634));
    SB_LUT4 add_13_add_1_21902_add_1_13_lut (.I0(GND_net), .I1(n282[11]), 
            .I2(n58[11]), .I3(n35897), .O(n57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_11_lut (.I0(GND_net), .I1(n16312[8]), .I2(GND_net), 
            .I3(n37546), .O(n16183[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3070_2 (.CI(GND_net), .I0(n56_adj_3696), .I1(n149_adj_3697), 
            .CO(n37441));
    SB_CARRY add_3079_3 (.CI(n37843), .I0(n9325[0]), .I1(n180), .CO(n37844));
    SB_LUT4 add_3060_11_lut (.I0(GND_net), .I1(n8157[8]), .I2(GND_net), 
            .I3(n37264), .O(n8131[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_8 (.CI(n36087), .I0(GND_net), .I1(n76[6]), 
            .CO(n36088));
    SB_LUT4 add_3079_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n8470[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3079_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3079_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n37843));
    SB_LUT4 mult_12_i221_2_lut (.I0(\Kd[3] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n328));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_24_lut (.I0(GND_net), .I1(n8446[21]), .I2(GND_net), 
            .I3(n37842), .O(n1804[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_9_lut (.I0(GND_net), .I1(n1800[6]), .I2(GND_net), 
            .I3(n37712), .O(n1799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n35995), .I0(GND_net), .I1(n75[8]), 
            .CO(n35996));
    SB_CARRY add_13_add_1_21902_add_1_13 (.CI(n35897), .I0(n282[11]), .I1(n58[11]), 
            .CO(n35898));
    SB_CARRY add_13_add_1_21902_add_1_31 (.CI(n35915), .I0(n7063[6]), .I1(n58[29]), 
            .CO(n35916));
    SB_CARRY add_3203_3 (.CI(n37021), .I0(n12155[0]), .I1(n180), .CO(n37022));
    SB_CARRY add_3047_9 (.CI(n36557), .I0(n9123[6]), .I1(GND_net), .CO(n36558));
    SB_LUT4 add_3333_9_lut (.I0(GND_net), .I1(n14791[6]), .I2(GND_net), 
            .I3(n36244), .O(n14432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n76[5]), 
            .I3(n36086), .O(n871)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n75[7]), .I3(n35994), .O(n15_adj_3702)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_70_add_3_7 (.CI(n36086), .I0(GND_net), .I1(n76[5]), 
            .CO(n36087));
    SB_LUT4 add_3069_16_lut (.I0(GND_net), .I1(n8346[13]), .I2(GND_net), 
            .I3(n37440), .O(n8329[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_8_lut (.I0(GND_net), .I1(n9123[5]), .I2(n686_adj_3704), 
            .I3(n36556), .O(n7758[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_8 (.CI(n36556), .I0(n9123[5]), .I1(n686_adj_3704), 
            .CO(n36557));
    SB_LUT4 mult_14_add_1219_23_lut (.I0(GND_net), .I1(n8446[20]), .I2(GND_net), 
            .I3(n37841), .O(n1804[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_14_lut (.I0(GND_net), .I1(n15397[11]), .I2(GND_net), 
            .I3(n37632), .O(n15112[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_14 (.CI(n37632), .I0(n15397[11]), .I1(GND_net), 
            .CO(n37633));
    SB_LUT4 unary_minus_70_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n76[4]), 
            .I3(n36085), .O(n872)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i333_2_lut (.I0(\Kd[5] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n495));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_21902_add_1_12_lut (.I0(GND_net), .I1(n282[10]), 
            .I2(n58[10]), .I3(n35896), .O(n57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_12 (.CI(n35896), .I0(n282[10]), .I1(n58[10]), 
            .CO(n35897));
    SB_LUT4 add_13_add_1_21902_add_1_11_lut (.I0(GND_net), .I1(n282[9]), 
            .I2(n58[9]), .I3(n35895), .O(n57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_11 (.CI(n35895), .I0(n282[9]), .I1(n58[9]), 
            .CO(n35896));
    SB_CARRY add_3060_11 (.CI(n37264), .I0(n8157[8]), .I1(GND_net), .CO(n37265));
    SB_LUT4 add_13_add_1_21902_add_1_10_lut (.I0(GND_net), .I1(n282[8]), 
            .I2(n58[8]), .I3(n35894), .O(n57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_7_lut (.I0(GND_net), .I1(n9123[4]), .I2(n589_adj_3706), 
            .I3(n36555), .O(n7758[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_7 (.CI(n36555), .I0(n9123[4]), .I1(n589_adj_3706), 
            .CO(n36556));
    SB_LUT4 add_3203_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n11529[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3203_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_10 (.CI(n35894), .I0(n282[8]), .I1(n58[8]), 
            .CO(n35895));
    SB_CARRY unary_minus_70_add_3_6 (.CI(n36085), .I0(GND_net), .I1(n76[4]), 
            .CO(n36086));
    SB_LUT4 add_3047_6_lut (.I0(GND_net), .I1(n9123[3]), .I2(n492_adj_3707), 
            .I3(n36554), .O(n7758[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n76[3]), 
            .I3(n36084), .O(n873)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_10_lut (.I0(GND_net), .I1(n8157[7]), .I2(GND_net), 
            .I3(n37263), .O(n8131[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3203_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n37021));
    SB_CARRY add_3060_10 (.CI(n37263), .I0(n8157[7]), .I1(GND_net), .CO(n37264));
    SB_LUT4 add_3069_15_lut (.I0(GND_net), .I1(n8346[12]), .I2(GND_net), 
            .I3(n37439), .O(n8329[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_23 (.CI(n37841), .I0(n8446[20]), .I1(GND_net), 
            .CO(n37842));
    SB_LUT4 add_13_add_1_21902_add_1_9_lut (.I0(GND_net), .I1(n282[7]), 
            .I2(n58[7]), .I3(n35893), .O(n57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_15 (.CI(n37439), .I0(n8346[12]), .I1(GND_net), .CO(n37440));
    SB_CARRY mult_14_add_1214_9 (.CI(n37712), .I0(n1800[6]), .I1(GND_net), 
            .CO(n37713));
    SB_CARRY add_3441_11 (.CI(n37546), .I0(n16312[8]), .I1(GND_net), .CO(n37547));
    SB_LUT4 add_3229_17_lut (.I0(GND_net), .I1(n12730[14]), .I2(GND_net), 
            .I3(n37020), .O(n12155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_9_lut (.I0(GND_net), .I1(n8157[6]), .I2(GND_net), 
            .I3(n37262), .O(n8131[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_9 (.CI(n37262), .I0(n8157[6]), .I1(GND_net), .CO(n37263));
    SB_LUT4 add_3370_13_lut (.I0(GND_net), .I1(n15397[10]), .I2(GND_net), 
            .I3(n37631), .O(n15112[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_8_lut (.I0(GND_net), .I1(n8157[5]), .I2(n701_adj_3709), 
            .I3(n37261), .O(n8131[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_14_lut (.I0(GND_net), .I1(n8346[11]), .I2(GND_net), 
            .I3(n37438), .O(n8329[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_10_lut (.I0(GND_net), .I1(n16312[7]), .I2(GND_net), 
            .I3(n37545), .O(n16183[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3229_16_lut (.I0(GND_net), .I1(n12730[13]), .I2(GND_net), 
            .I3(n37019), .O(n12155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_13 (.CI(n37631), .I0(n15397[10]), .I1(GND_net), 
            .CO(n37632));
    SB_LUT4 mult_14_add_1214_8_lut (.I0(GND_net), .I1(n1800[5]), .I2(n521), 
            .I3(n37711), .O(n1799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_12_lut (.I0(GND_net), .I1(n15397[9]), .I2(GND_net), 
            .I3(n37630), .O(n15112[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_22_lut (.I0(GND_net), .I1(n8446[19]), .I2(GND_net), 
            .I3(n37840), .O(n1804[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_8 (.CI(n37711), .I0(n1800[5]), .I1(n521), 
            .CO(n37712));
    SB_CARRY add_13_add_1_21902_add_1_9 (.CI(n35893), .I0(n282[7]), .I1(n58[7]), 
            .CO(n35894));
    SB_CARRY add_3229_16 (.CI(n37019), .I0(n12730[13]), .I1(GND_net), 
            .CO(n37020));
    SB_LUT4 add_13_add_1_21902_add_1_8_lut (.I0(GND_net), .I1(n282[6]), 
            .I2(n58[6]), .I3(n35892), .O(n57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_10 (.CI(n37545), .I0(n16312[7]), .I1(GND_net), .CO(n37546));
    SB_LUT4 add_3441_9_lut (.I0(GND_net), .I1(n16312[6]), .I2(GND_net), 
            .I3(n37544), .O(n16183[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_12 (.CI(n37630), .I0(n15397[9]), .I1(GND_net), .CO(n37631));
    SB_CARRY add_3333_9 (.CI(n36244), .I0(n14791[6]), .I1(GND_net), .CO(n36245));
    SB_CARRY mult_14_add_1219_22 (.CI(n37840), .I0(n8446[19]), .I1(GND_net), 
            .CO(n37841));
    SB_LUT4 add_3370_11_lut (.I0(GND_net), .I1(n15397[8]), .I2(GND_net), 
            .I3(n37629), .O(n15112[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_8 (.CI(n35892), .I0(n282[6]), .I1(n58[6]), 
            .CO(n35893));
    SB_LUT4 mult_14_add_1219_21_lut (.I0(GND_net), .I1(n8446[18]), .I2(GND_net), 
            .I3(n37839), .O(n1804[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_7_lut (.I0(GND_net), .I1(n1800[4]), .I2(n448_c), 
            .I3(n37710), .O(n1799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_21 (.CI(n37839), .I0(n8446[18]), .I1(GND_net), 
            .CO(n37840));
    SB_LUT4 mult_14_add_1219_20_lut (.I0(GND_net), .I1(n8446[17]), .I2(GND_net), 
            .I3(n37838), .O(n1804[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i495_2_lut (.I0(\Kd[7] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i495_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1219_20 (.CI(n37838), .I0(n8446[17]), .I1(GND_net), 
            .CO(n37839));
    SB_CARRY mult_14_add_1214_7 (.CI(n37710), .I0(n1800[4]), .I1(n448_c), 
            .CO(n37711));
    SB_CARRY add_3069_14 (.CI(n37438), .I0(n8346[11]), .I1(GND_net), .CO(n37439));
    SB_CARRY add_3441_9 (.CI(n37544), .I0(n16312[6]), .I1(GND_net), .CO(n37545));
    SB_LUT4 add_3229_15_lut (.I0(GND_net), .I1(n12730[12]), .I2(GND_net), 
            .I3(n37018), .O(n12155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3047_6 (.CI(n36554), .I0(n9123[3]), .I1(n492_adj_3707), 
            .CO(n36555));
    SB_CARRY add_3229_15 (.CI(n37018), .I0(n12730[12]), .I1(GND_net), 
            .CO(n37019));
    SB_CARRY unary_minus_70_add_3_5 (.CI(n36084), .I0(GND_net), .I1(n76[3]), 
            .CO(n36085));
    SB_LUT4 mult_12_i398_2_lut (.I0(\Kd[6] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n592_adj_3404));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3229_14_lut (.I0(GND_net), .I1(n12730[11]), .I2(GND_net), 
            .I3(n37017), .O(n12155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_8 (.CI(n37261), .I0(n8157[5]), .I1(n701_adj_3709), 
            .CO(n37262));
    SB_CARRY add_3229_14 (.CI(n37017), .I0(n12730[11]), .I1(GND_net), 
            .CO(n37018));
    SB_LUT4 add_3229_13_lut (.I0(GND_net), .I1(n12730[10]), .I2(GND_net), 
            .I3(n37016), .O(n12155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_13_lut (.I0(GND_net), .I1(n8346[10]), .I2(GND_net), 
            .I3(n37437), .O(n8329[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_7_lut (.I0(GND_net), .I1(n8157[4]), .I2(n604_adj_3712), 
            .I3(n37260), .O(n8131[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_13 (.CI(n37016), .I0(n12730[10]), .I1(GND_net), 
            .CO(n37017));
    SB_LUT4 add_3229_12_lut (.I0(GND_net), .I1(n12730[9]), .I2(GND_net), 
            .I3(n37015), .O(n12155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_7 (.CI(n37260), .I0(n8157[4]), .I1(n604_adj_3712), 
            .CO(n37261));
    SB_CARRY add_3229_12 (.CI(n37015), .I0(n12730[9]), .I1(GND_net), .CO(n37016));
    SB_LUT4 add_3229_11_lut (.I0(GND_net), .I1(n12730[8]), .I2(GND_net), 
            .I3(n37014), .O(n12155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_8_lut (.I0(GND_net), .I1(n16312[5]), .I2(n737_adj_3713), 
            .I3(n37543), .O(n16183[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_13 (.CI(n37437), .I0(n8346[10]), .I1(GND_net), .CO(n37438));
    SB_LUT4 add_3060_6_lut (.I0(GND_net), .I1(n8157[3]), .I2(n507_adj_3714), 
            .I3(n37259), .O(n8131[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_11 (.CI(n37014), .I0(n12730[8]), .I1(GND_net), .CO(n37015));
    SB_LUT4 add_3229_10_lut (.I0(GND_net), .I1(n12730[7]), .I2(GND_net), 
            .I3(n37013), .O(n12155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_6 (.CI(n37259), .I0(n8157[3]), .I1(n507_adj_3714), 
            .CO(n37260));
    SB_CARRY add_3229_10 (.CI(n37013), .I0(n12730[7]), .I1(GND_net), .CO(n37014));
    SB_LUT4 add_3229_9_lut (.I0(GND_net), .I1(n12730[6]), .I2(GND_net), 
            .I3(n37012), .O(n12155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_12_lut (.I0(GND_net), .I1(n8346[9]), .I2(GND_net), 
            .I3(n37436), .O(n8329[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_5_lut (.I0(GND_net), .I1(n8157[2]), .I2(n410_adj_3715), 
            .I3(n37258), .O(n8131[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_9 (.CI(n37012), .I0(n12730[6]), .I1(GND_net), .CO(n37013));
    SB_LUT4 add_3229_8_lut (.I0(GND_net), .I1(n12730[5]), .I2(n545), .I3(n37011), 
            .O(n12155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_5 (.CI(n37258), .I0(n8157[2]), .I1(n410_adj_3715), 
            .CO(n37259));
    SB_CARRY add_3229_8 (.CI(n37011), .I0(n12730[5]), .I1(n545), .CO(n37012));
    SB_LUT4 add_3229_7_lut (.I0(GND_net), .I1(n12730[4]), .I2(n472), .I3(n37010), 
            .O(n12155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_6_lut (.I0(GND_net), .I1(n1800[3]), .I2(n375), 
            .I3(n37709), .O(n1799[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_11 (.CI(n37629), .I0(n15397[8]), .I1(GND_net), .CO(n37630));
    SB_CARRY add_3441_8 (.CI(n37543), .I0(n16312[5]), .I1(n737_adj_3713), 
            .CO(n37544));
    SB_CARRY add_3069_12 (.CI(n37436), .I0(n8346[9]), .I1(GND_net), .CO(n37437));
    SB_LUT4 add_3060_4_lut (.I0(GND_net), .I1(n8157[1]), .I2(n313_adj_3716), 
            .I3(n37257), .O(n8131[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_7 (.CI(n37010), .I0(n12730[4]), .I1(n472), .CO(n37011));
    SB_CARRY add_3060_4 (.CI(n37257), .I0(n8157[1]), .I1(n313_adj_3716), 
            .CO(n37258));
    SB_LUT4 add_3069_11_lut (.I0(GND_net), .I1(n8346[8]), .I2(GND_net), 
            .I3(n37435), .O(n8329[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3060_3_lut (.I0(GND_net), .I1(n8157[0]), .I2(n216_adj_3717), 
            .I3(n37256), .O(n8131[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3229_6_lut (.I0(GND_net), .I1(n12730[3]), .I2(n399_c), 
            .I3(n37009), .O(n12155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_5_lut (.I0(GND_net), .I1(n9123[2]), .I2(n395_adj_3718), 
            .I3(n36553), .O(n7758[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_8_lut (.I0(GND_net), .I1(n14791[5]), .I2(n716_adj_3719), 
            .I3(n36243), .O(n14432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_6 (.CI(n37009), .I0(n12730[3]), .I1(n399_c), .CO(n37010));
    SB_CARRY add_3047_5 (.CI(n36553), .I0(n9123[2]), .I1(n395_adj_3718), 
            .CO(n36554));
    SB_CARRY add_3333_8 (.CI(n36243), .I0(n14791[5]), .I1(n716_adj_3719), 
            .CO(n36244));
    SB_LUT4 add_3333_7_lut (.I0(GND_net), .I1(n14791[4]), .I2(n619_adj_3720), 
            .I3(n36242), .O(n14432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3047_4_lut (.I0(GND_net), .I1(n9123[1]), .I2(n298_adj_3721), 
            .I3(n36552), .O(n7758[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_7 (.CI(n36242), .I0(n14791[4]), .I1(n619_adj_3720), 
            .CO(n36243));
    SB_CARRY add_3047_4 (.CI(n36552), .I0(n9123[1]), .I1(n298_adj_3721), 
            .CO(n36553));
    SB_LUT4 add_3047_3_lut (.I0(GND_net), .I1(n9123[0]), .I2(n201_adj_3722), 
            .I3(n36551), .O(n7758[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_7_lut (.I0(GND_net), .I1(n282[5]), 
            .I2(n58[5]), .I3(n35891), .O(n57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_19_lut (.I0(GND_net), .I1(n8446[16]), .I2(GND_net), 
            .I3(n37837), .O(n1804[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_7_lut (.I0(GND_net), .I1(n16312[4]), .I2(n640_adj_3723), 
            .I3(n37542), .O(n16183[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n76[2]), 
            .I3(n36083), .O(n874)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_19 (.CI(n37837), .I0(n8446[16]), .I1(GND_net), 
            .CO(n37838));
    SB_CARRY add_3441_7 (.CI(n37542), .I0(n16312[4]), .I1(n640_adj_3723), 
            .CO(n37543));
    SB_LUT4 add_3370_10_lut (.I0(GND_net), .I1(n15397[7]), .I2(GND_net), 
            .I3(n37628), .O(n15112[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_4 (.CI(n36083), .I0(GND_net), .I1(n76[2]), 
            .CO(n36084));
    SB_LUT4 add_3441_6_lut (.I0(GND_net), .I1(n16312[3]), .I2(n543_adj_3725), 
            .I3(n37541), .O(n16183[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_11 (.CI(n37435), .I0(n8346[8]), .I1(GND_net), .CO(n37436));
    SB_DFFE \PID_CONTROLLER.integral_1015__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[0]));   // verilog/motorControl.v(41[21:33])
    SB_LUT4 unary_minus_70_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n76[1]), 
            .I3(n36082), .O(n875)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_6_lut (.I0(GND_net), .I1(n14791[3]), .I2(n522_adj_3728), 
            .I3(n36241), .O(n14432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_3 (.CI(n37256), .I0(n8157[0]), .I1(n216_adj_3717), 
            .CO(n37257));
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i286_2_lut (.I0(\Kd[4] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n425));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i292_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n434));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3505));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3229_5_lut (.I0(GND_net), .I1(n12730[2]), .I2(n326), .I3(n37008), 
            .O(n12155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_5 (.CI(n37008), .I0(n12730[2]), .I1(n326), .CO(n37009));
    SB_CARRY add_3047_3 (.CI(n36551), .I0(n9123[0]), .I1(n201_adj_3722), 
            .CO(n36552));
    SB_CARRY unary_minus_70_add_3_3 (.CI(n36082), .I0(GND_net), .I1(n76[1]), 
            .CO(n36083));
    SB_CARRY add_3333_6 (.CI(n36241), .I0(n14791[3]), .I1(n522_adj_3728), 
            .CO(n36242));
    SB_LUT4 add_3047_2_lut (.I0(GND_net), .I1(n11_adj_3729), .I2(n104_adj_3730), 
            .I3(GND_net), .O(n7758[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3047_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_2_lut (.I0(n28817), .I1(GND_net), .I2(n76[0]), 
            .I3(VCC_net), .O(n46619)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_13_add_1_21902_add_1_7 (.CI(n35891), .I0(n282[5]), .I1(n58[5]), 
            .CO(n35892));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n35994), .I0(GND_net), .I1(n75[7]), 
            .CO(n35995));
    SB_LUT4 add_13_add_1_21902_add_1_6_lut (.I0(GND_net), .I1(n282[4]), 
            .I2(n58[4]), .I3(n35890), .O(n57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3229_4_lut (.I0(GND_net), .I1(n12730[1]), .I2(n253), .I3(n37007), 
            .O(n12155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_5_lut (.I0(GND_net), .I1(n14791[2]), .I2(n425_adj_3732), 
            .I3(n36240), .O(n14432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i463_2_lut (.I0(\Kd[7] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n689));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_13_add_1_21902_add_1_6 (.CI(n35890), .I0(n282[4]), .I1(n58[4]), 
            .CO(n35891));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n75[6]), .I3(n35993), .O(n13_adj_3733)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3047_2 (.CI(GND_net), .I0(n11_adj_3729), .I1(n104_adj_3730), 
            .CO(n36551));
    SB_LUT4 mult_14_add_1219_18_lut (.I0(GND_net), .I1(n8446[15]), .I2(GND_net), 
            .I3(n37836), .O(n1804[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_18 (.CI(n37836), .I0(n8446[15]), .I1(GND_net), 
            .CO(n37837));
    SB_CARRY mult_14_add_1214_6 (.CI(n37709), .I0(n1800[3]), .I1(n375), 
            .CO(n37710));
    SB_LUT4 mult_14_add_1219_17_lut (.I0(GND_net), .I1(n8446[14]), .I2(GND_net), 
            .I3(n37835), .O(n1804[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_17 (.CI(n37835), .I0(n8446[14]), .I1(GND_net), 
            .CO(n37836));
    SB_CARRY unary_minus_5_add_3_8 (.CI(n35993), .I0(GND_net), .I1(n75[6]), 
            .CO(n35994));
    SB_CARRY add_3333_5 (.CI(n36240), .I0(n14791[2]), .I1(n425_adj_3732), 
            .CO(n36241));
    SB_LUT4 add_3333_4_lut (.I0(GND_net), .I1(n14791[1]), .I2(n328_adj_3735), 
            .I3(n36239), .O(n14432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_5_lut (.I0(GND_net), .I1(n1800[2]), .I2(n302_adj_3737), 
            .I3(n37708), .O(n1799[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3277_15_lut (.I0(GND_net), .I1(n13732[12]), .I2(GND_net), 
            .I3(n36550), .O(n13254[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n75[5]), .I3(n35992), .O(n11_adj_3738)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3060_2_lut (.I0(GND_net), .I1(n26_adj_3740), .I2(n119_adj_3741), 
            .I3(GND_net), .O(n8131[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3060_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_16_lut (.I0(GND_net), .I1(n8446[13]), .I2(GND_net), 
            .I3(n37834), .O(n1804[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3277_14_lut (.I0(GND_net), .I1(n13732[11]), .I2(GND_net), 
            .I3(n36549), .O(n13254[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_4 (.CI(n36239), .I0(n14791[1]), .I1(n328_adj_3735), 
            .CO(n36240));
    SB_CARRY add_3277_14 (.CI(n36549), .I0(n13732[11]), .I1(GND_net), 
            .CO(n36550));
    SB_CARRY mult_14_add_1219_16 (.CI(n37834), .I0(n8446[13]), .I1(GND_net), 
            .CO(n37835));
    SB_CARRY mult_14_add_1214_5 (.CI(n37708), .I0(n1800[2]), .I1(n302_adj_3737), 
            .CO(n37709));
    SB_LUT4 mult_14_add_1219_15_lut (.I0(GND_net), .I1(n8446[12]), .I2(GND_net), 
            .I3(n37833), .O(n1804[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_15 (.CI(n37833), .I0(n8446[12]), .I1(GND_net), 
            .CO(n37834));
    SB_LUT4 add_3277_13_lut (.I0(GND_net), .I1(n13732[10]), .I2(GND_net), 
            .I3(n36548), .O(n13254[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3333_3_lut (.I0(GND_net), .I1(n14791[0]), .I2(n231_adj_3742), 
            .I3(n36238), .O(n14432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n76[0]), 
            .CO(n36082));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n35992), .I0(GND_net), .I1(n75[5]), 
            .CO(n35993));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n75[4]), .I3(n35991), .O(n9_adj_3743)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_13_add_1_21902_add_1_5_lut (.I0(GND_net), .I1(n282[3]), 
            .I2(n58[3]), .I3(n35889), .O(n57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n35991), .I0(GND_net), .I1(n75[4]), 
            .CO(n35992));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n75[3]), .I3(n35990), .O(n7_adj_3745)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3333_3 (.CI(n36238), .I0(n14791[0]), .I1(n231_adj_3742), 
            .CO(n36239));
    SB_CARRY add_3277_13 (.CI(n36548), .I0(n13732[10]), .I1(GND_net), 
            .CO(n36549));
    SB_LUT4 add_3277_12_lut (.I0(GND_net), .I1(n13732[9]), .I2(GND_net), 
            .I3(n36547), .O(n13254[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3277_12 (.CI(n36547), .I0(n13732[9]), .I1(GND_net), .CO(n36548));
    SB_CARRY add_3229_4 (.CI(n37007), .I0(n12730[1]), .I1(n253), .CO(n37008));
    SB_LUT4 mult_12_i351_2_lut (.I0(\Kd[5] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n522));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3229_3_lut (.I0(GND_net), .I1(n12730[0]), .I2(n180), .I3(n37006), 
            .O(n12155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3060_2 (.CI(GND_net), .I0(n26_adj_3740), .I1(n119_adj_3741), 
            .CO(n37256));
    SB_LUT4 mult_12_i111_2_lut (.I0(\Kd[1] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n164));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3333_2_lut (.I0(GND_net), .I1(n41_adj_3747), .I2(n134_adj_3748), 
            .I3(GND_net), .O(n14432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3333_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i48_2_lut (.I0(\Kd[0] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n71));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i416_2_lut (.I0(\Kd[6] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n619));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n534));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3069_10_lut (.I0(GND_net), .I1(n8346[7]), .I2(GND_net), 
            .I3(n37434), .O(n8329[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3277_11_lut (.I0(GND_net), .I1(n13732[8]), .I2(GND_net), 
            .I3(n36546), .O(n13254[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3333_2 (.CI(GND_net), .I0(n41_adj_3747), .I1(n134_adj_3748), 
            .CO(n36238));
    SB_LUT4 mult_14_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3059_26_lut (.I0(GND_net), .I1(n8131[23]), .I2(GND_net), 
            .I3(n37255), .O(n8104[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_3 (.CI(n37006), .I0(n12730[0]), .I1(n180), .CO(n37007));
    SB_LUT4 mult_12_i481_2_lut (.I0(\Kd[7] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n716));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3059_25_lut (.I0(GND_net), .I1(n8131[22]), .I2(GND_net), 
            .I3(n37254), .O(n8104[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3229_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n12155[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3229_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3277_11 (.CI(n36546), .I0(n13732[8]), .I1(GND_net), .CO(n36547));
    SB_LUT4 mult_14_add_1214_4_lut (.I0(GND_net), .I1(n1800[1]), .I2(n229_adj_3750), 
            .I3(n37707), .O(n1799[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_10_lut (.I0(GND_net), .I1(n16569[7]), .I2(GND_net), 
            .I3(n36237), .O(n16503[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_6 (.CI(n37541), .I0(n16312[3]), .I1(n543_adj_3725), 
            .CO(n37542));
    SB_LUT4 add_3277_10_lut (.I0(GND_net), .I1(n13732[7]), .I2(GND_net), 
            .I3(n36545), .O(n13254[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_10 (.CI(n37628), .I0(n15397[7]), .I1(GND_net), .CO(n37629));
    SB_LUT4 mult_14_add_1219_14_lut (.I0(GND_net), .I1(n8446[11]), .I2(GND_net), 
            .I3(n37832), .O(n1804[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i176_2_lut (.I0(\Kd[2] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n261));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i176_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1219_14 (.CI(n37832), .I0(n8446[11]), .I1(GND_net), 
            .CO(n37833));
    SB_CARRY add_13_add_1_21902_add_1_5 (.CI(n35889), .I0(n282[3]), .I1(n58[3]), 
            .CO(n35890));
    SB_LUT4 add_3370_9_lut (.I0(GND_net), .I1(n15397[6]), .I2(GND_net), 
            .I3(n37627), .O(n15112[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_13_lut (.I0(GND_net), .I1(n8446[10]), .I2(GND_net), 
            .I3(n37831), .O(n1804[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_25 (.CI(n37254), .I0(n8131[22]), .I1(GND_net), .CO(n37255));
    SB_CARRY add_3277_10 (.CI(n36545), .I0(n13732[7]), .I1(GND_net), .CO(n36546));
    SB_LUT4 add_3277_9_lut (.I0(GND_net), .I1(n13732[6]), .I2(GND_net), 
            .I3(n36544), .O(n13254[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_10 (.CI(n37434), .I0(n8346[7]), .I1(GND_net), .CO(n37435));
    SB_LUT4 add_3441_5_lut (.I0(GND_net), .I1(n16312[2]), .I2(n446_adj_3751), 
            .I3(n37540), .O(n16183[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_9_lut (.I0(GND_net), .I1(n16569[6]), .I2(GND_net), 
            .I3(n36236), .O(n16503[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_24_lut (.I0(GND_net), .I1(n8131[21]), .I2(GND_net), 
            .I3(n37253), .O(n8104[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_4 (.CI(n37707), .I0(n1800[1]), .I1(n229_adj_3750), 
            .CO(n37708));
    SB_CARRY add_3441_5 (.CI(n37540), .I0(n16312[2]), .I1(n446_adj_3751), 
            .CO(n37541));
    SB_CARRY mult_14_add_1219_13 (.CI(n37831), .I0(n8446[10]), .I1(GND_net), 
            .CO(n37832));
    SB_CARRY add_3059_24 (.CI(n37253), .I0(n8131[21]), .I1(GND_net), .CO(n37254));
    SB_CARRY add_3370_9 (.CI(n37627), .I0(n15397[6]), .I1(GND_net), .CO(n37628));
    SB_LUT4 add_3059_23_lut (.I0(GND_net), .I1(n8131[20]), .I2(GND_net), 
            .I3(n37252), .O(n8104[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n35990), .I0(GND_net), .I1(n75[3]), 
            .CO(n35991));
    SB_LUT4 add_3069_9_lut (.I0(GND_net), .I1(n8346[6]), .I2(GND_net), 
            .I3(n37433), .O(n8329[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3441_4_lut (.I0(GND_net), .I1(n16312[1]), .I2(n349_adj_3752), 
            .I3(n37539), .O(n16183[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_9 (.CI(n36236), .I0(n16569[6]), .I1(GND_net), .CO(n36237));
    SB_CARRY add_3277_9 (.CI(n36544), .I0(n13732[6]), .I1(GND_net), .CO(n36545));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n75[2]), .I3(n35989), .O(n5_adj_3753)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3471_8_lut (.I0(GND_net), .I1(n16569[5]), .I2(n746_adj_3755), 
            .I3(n36235), .O(n16503[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3277_8_lut (.I0(GND_net), .I1(n13732[5]), .I2(n545), .I3(n36543), 
            .O(n13254[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3229_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n37006));
    SB_LUT4 add_3370_8_lut (.I0(GND_net), .I1(n15397[5]), .I2(n722_adj_3756), 
            .I3(n37626), .O(n15112[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_9 (.CI(n37433), .I0(n8346[6]), .I1(GND_net), .CO(n37434));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n35989), .I0(GND_net), .I1(n75[2]), 
            .CO(n35990));
    SB_CARRY add_3277_8 (.CI(n36543), .I0(n13732[5]), .I1(n545), .CO(n36544));
    SB_LUT4 add_3277_7_lut (.I0(GND_net), .I1(n13732[4]), .I2(n472), .I3(n36542), 
            .O(n13254[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_8 (.CI(n36235), .I0(n16569[5]), .I1(n746_adj_3755), 
            .CO(n36236));
    SB_LUT4 add_3471_7_lut (.I0(GND_net), .I1(n16569[4]), .I2(n649_adj_3757), 
            .I3(n36234), .O(n16503[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n75[1]), .I3(n35988), .O(n3_adj_3758)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3441_4 (.CI(n37539), .I0(n16312[1]), .I1(n349_adj_3752), 
            .CO(n37540));
    SB_LUT4 add_3069_8_lut (.I0(GND_net), .I1(n8346[5]), .I2(n728_adj_3760), 
            .I3(n37432), .O(n8329[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_23 (.CI(n37252), .I0(n8131[20]), .I1(GND_net), .CO(n37253));
    SB_CARRY add_3370_8 (.CI(n37626), .I0(n15397[5]), .I1(n722_adj_3756), 
            .CO(n37627));
    SB_CARRY unary_minus_5_add_3_3 (.CI(n35988), .I0(GND_net), .I1(n75[1]), 
            .CO(n35989));
    SB_CARRY add_3069_8 (.CI(n37432), .I0(n8346[5]), .I1(n728_adj_3760), 
            .CO(n37433));
    SB_LUT4 add_3059_22_lut (.I0(GND_net), .I1(n8131[19]), .I2(GND_net), 
            .I3(n37251), .O(n8104[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_22 (.CI(n37251), .I0(n8131[19]), .I1(GND_net), .CO(n37252));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n75[0]), 
            .I3(VCC_net), .O(n73[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_7 (.CI(n36234), .I0(n16569[4]), .I1(n649_adj_3757), 
            .CO(n36235));
    SB_CARRY add_3277_7 (.CI(n36542), .I0(n13732[4]), .I1(n472), .CO(n36543));
    SB_LUT4 add_3441_3_lut (.I0(GND_net), .I1(n16312[0]), .I2(n252_adj_3763), 
            .I3(n37538), .O(n16183[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_7_lut (.I0(GND_net), .I1(n8346[4]), .I2(n631_adj_3764), 
            .I3(n37431), .O(n8329[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_3 (.CI(n37538), .I0(n16312[0]), .I1(n252_adj_3763), 
            .CO(n37539));
    SB_LUT4 add_3059_21_lut (.I0(GND_net), .I1(n8131[18]), .I2(GND_net), 
            .I3(n37250), .O(n8104[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_7_lut (.I0(GND_net), .I1(n15397[4]), .I2(n625_adj_3765), 
            .I3(n37625), .O(n15112[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i241_2_lut (.I0(\Kd[3] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n358));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3441_2_lut (.I0(GND_net), .I1(n62_adj_3766), .I2(n155_adj_3767), 
            .I3(GND_net), .O(n16183[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3441_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_7 (.CI(n37431), .I0(n8346[4]), .I1(n631_adj_3764), 
            .CO(n37432));
    SB_CARRY add_3059_21 (.CI(n37250), .I0(n8131[18]), .I1(GND_net), .CO(n37251));
    SB_LUT4 add_3277_6_lut (.I0(GND_net), .I1(n13732[3]), .I2(n399_c), 
            .I3(n36541), .O(n13254[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_6_lut (.I0(GND_net), .I1(n16569[3]), .I2(n552_adj_3768), 
            .I3(n36233), .O(n16503[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_3_lut (.I0(GND_net), .I1(n1800[0]), .I2(n156_adj_3769), 
            .I3(n37706), .O(n1799[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3277_6 (.CI(n36541), .I0(n13732[3]), .I1(n399_c), .CO(n36542));
    SB_LUT4 add_3277_5_lut (.I0(GND_net), .I1(n13732[2]), .I2(n326), .I3(n36540), 
            .O(n13254[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n631));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3471_6 (.CI(n36233), .I0(n16569[3]), .I1(n552_adj_3768), 
            .CO(n36234));
    SB_CARRY add_3277_5 (.CI(n36540), .I0(n13732[2]), .I1(n326), .CO(n36541));
    SB_LUT4 add_3471_5_lut (.I0(GND_net), .I1(n16569[2]), .I2(n455_adj_3770), 
            .I3(n36232), .O(n16503[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3277_4_lut (.I0(GND_net), .I1(n13732[1]), .I2(n253), .I3(n36539), 
            .O(n13254[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3069_6_lut (.I0(GND_net), .I1(n8346[3]), .I2(n534_adj_3771), 
            .I3(n37430), .O(n8329[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_6 (.CI(n37430), .I0(n8346[3]), .I1(n534_adj_3771), 
            .CO(n37431));
    SB_CARRY add_3277_4 (.CI(n36539), .I0(n13732[1]), .I1(n253), .CO(n36540));
    SB_LUT4 mult_12_i306_2_lut (.I0(\Kd[4] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n455_c));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3471_5 (.CI(n36232), .I0(n16569[2]), .I1(n455_adj_3770), 
            .CO(n36233));
    SB_LUT4 add_13_add_1_21902_add_1_4_lut (.I0(GND_net), .I1(n282[2]), 
            .I2(n58[2]), .I3(n35888), .O(n57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3441_2 (.CI(GND_net), .I0(n62_adj_3766), .I1(n155_adj_3767), 
            .CO(n37538));
    SB_LUT4 mult_10_i489_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n728));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3069_5_lut (.I0(GND_net), .I1(n8346[2]), .I2(n437_adj_3772), 
            .I3(n37429), .O(n8329[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_4_lut (.I0(GND_net), .I1(n16569[1]), .I2(n358_adj_3773), 
            .I3(n36231), .O(n16503[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_5 (.CI(n37429), .I0(n8346[2]), .I1(n437_adj_3772), 
            .CO(n37430));
    SB_LUT4 add_3277_3_lut (.I0(GND_net), .I1(n13732[0]), .I2(n180), .I3(n36538), 
            .O(n13254[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_23_lut (.I0(GND_net), .I1(n8470[20]), .I2(GND_net), 
            .I3(n37537), .O(n8446[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i249_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3471_4 (.CI(n36231), .I0(n16569[1]), .I1(n358_adj_3773), 
            .CO(n36232));
    SB_LUT4 mult_12_i371_2_lut (.I0(\Kd[5] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n552));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3277_3 (.CI(n36538), .I0(n13732[0]), .I1(n180), .CO(n36539));
    SB_LUT4 add_3471_3_lut (.I0(GND_net), .I1(n16569[0]), .I2(n261_adj_3774), 
            .I3(n36230), .O(n16503[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3277_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n13254[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3277_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_3 (.CI(n36230), .I0(n16569[0]), .I1(n261_adj_3774), 
            .CO(n36231));
    SB_LUT4 mult_12_i436_2_lut (.I0(\Kd[6] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n649));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i436_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1214_3 (.CI(n37706), .I0(n1800[0]), .I1(n156_adj_3769), 
            .CO(n37707));
    SB_CARRY add_13_add_1_21902_add_1_4 (.CI(n35888), .I0(n282[2]), .I1(n58[2]), 
            .CO(n35889));
    SB_LUT4 add_3059_20_lut (.I0(GND_net), .I1(n8131[17]), .I2(GND_net), 
            .I3(n37249), .O(n8104[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3277_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n36538));
    SB_LUT4 mult_12_i501_2_lut (.I0(\Kd[7] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_12_lut (.I0(GND_net), .I1(n8446[9]), .I2(GND_net), 
            .I3(n37830), .O(n1804[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_29_lut (.I0(GND_net), .I1(n9927[26]), .I2(GND_net), 
            .I3(n36537), .O(n9123[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_21902_add_1_3_lut (.I0(GND_net), .I1(n282[1]), 
            .I2(n58[1]), .I3(n35887), .O(n57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_2_lut (.I0(GND_net), .I1(n71_adj_3775), .I2(n164_adj_3776), 
            .I3(GND_net), .O(n16503[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_2 (.CI(GND_net), .I0(n71_adj_3775), .I1(n164_adj_3776), 
            .CO(n36230));
    SB_LUT4 add_3101_28_lut (.I0(GND_net), .I1(n9927[25]), .I2(GND_net), 
            .I3(n36536), .O(n9123[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_28 (.CI(n36536), .I0(n9927[25]), .I1(GND_net), .CO(n36537));
    SB_LUT4 add_3101_27_lut (.I0(GND_net), .I1(n9927[24]), .I2(GND_net), 
            .I3(n36535), .O(n9123[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_12 (.CI(n37830), .I0(n8446[9]), .I1(GND_net), 
            .CO(n37831));
    SB_CARRY add_3101_27 (.CI(n36535), .I0(n9927[24]), .I1(GND_net), .CO(n36536));
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n75[0]), 
            .CO(n35988));
    SB_LUT4 mult_14_add_1219_11_lut (.I0(GND_net), .I1(n8446[8]), .I2(GND_net), 
            .I3(n37829), .O(n1804[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_26_lut (.I0(GND_net), .I1(GND_net), .I2(n79[31]), 
            .I3(n35987), .O(pwm_23__N_2960[24])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n79[31]), 
            .I3(n35986), .O(pwm_23__N_2960[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_26_lut (.I0(GND_net), .I1(n9927[23]), .I2(GND_net), 
            .I3(n36534), .O(n9123[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_26 (.CI(n36534), .I0(n9927[23]), .I1(GND_net), .CO(n36535));
    SB_LUT4 mult_14_add_1214_2_lut (.I0(GND_net), .I1(n14_adj_3778), .I2(n83), 
            .I3(GND_net), .O(n1799[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_2 (.CI(GND_net), .I0(n14_adj_3778), .I1(n83), 
            .CO(n37706));
    SB_CARRY add_3370_7 (.CI(n37625), .I0(n15397[4]), .I1(n625_adj_3765), 
            .CO(n37626));
    SB_LUT4 unary_minus_21_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[1]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1213_24_lut (.I0(GND_net), .I1(n1799[21]), .I2(GND_net), 
            .I3(n37704), .O(n1798[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_22_lut (.I0(GND_net), .I1(n8470[19]), .I2(GND_net), 
            .I3(n37536), .O(n8446[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_21902_add_1_3 (.CI(n35887), .I0(n282[1]), .I1(n58[1]), 
            .CO(n35888));
    SB_LUT4 add_3101_25_lut (.I0(GND_net), .I1(n9927[22]), .I2(GND_net), 
            .I3(n36533), .O(n9123[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i274_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n407_c));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3069_4_lut (.I0(GND_net), .I1(n8346[1]), .I2(n340_adj_3779), 
            .I3(n37428), .O(n8329[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i339_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n504));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i93_2_lut (.I0(\Kd[1] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n137));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i93_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_17_add_3_25 (.CI(n35986), .I0(GND_net), .I1(n79[31]), 
            .CO(n35987));
    SB_LUT4 add_13_add_1_21902_add_1_2_lut (.I0(GND_net), .I1(n282[0]), 
            .I2(n58[0]), .I3(GND_net), .O(n57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_21902_add_1_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n79[22]), 
            .I3(n35985), .O(pwm_23__N_2960[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_4 (.CI(n37428), .I0(n8346[1]), .I1(n340_adj_3779), 
            .CO(n37429));
    SB_LUT4 add_3370_6_lut (.I0(GND_net), .I1(n15397[3]), .I2(n528_adj_3783), 
            .I3(n37624), .O(n15112[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_22 (.CI(n37536), .I0(n8470[19]), .I1(GND_net), .CO(n37537));
    SB_LUT4 mult_12_i30_2_lut (.I0(\Kd[0] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_3398));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3069_3_lut (.I0(GND_net), .I1(n8346[0]), .I2(n243_adj_3784), 
            .I3(n37427), .O(n8329[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_20 (.CI(n37249), .I0(n8131[17]), .I1(GND_net), .CO(n37250));
    SB_LUT4 add_3059_19_lut (.I0(GND_net), .I1(n8131[16]), .I2(GND_net), 
            .I3(n37248), .O(n8104[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3069_3 (.CI(n37427), .I0(n8346[0]), .I1(n243_adj_3784), 
            .CO(n37428));
    SB_CARRY add_13_add_1_21902_add_1_2 (.CI(GND_net), .I0(n282[0]), .I1(n58[0]), 
            .CO(n35887));
    SB_LUT4 add_3069_2_lut (.I0(GND_net), .I1(n53_adj_3785), .I2(n146_adj_3786), 
            .I3(GND_net), .O(n8329[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3069_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_11 (.CI(n37829), .I0(n8446[8]), .I1(GND_net), 
            .CO(n37830));
    SB_LUT4 mult_14_add_1219_10_lut (.I0(GND_net), .I1(n8446[7]), .I2(GND_net), 
            .I3(n37828), .O(n1804[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_10 (.CI(n37828), .I0(n8446[7]), .I1(GND_net), 
            .CO(n37829));
    SB_LUT4 mult_14_add_1219_9_lut (.I0(GND_net), .I1(n8446[6]), .I2(GND_net), 
            .I3(n37827), .O(n1804[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_6 (.CI(n37624), .I0(n15397[3]), .I1(n528_adj_3783), 
            .CO(n37625));
    SB_CARRY mult_14_add_1219_9 (.CI(n37827), .I0(n8446[6]), .I1(GND_net), 
            .CO(n37828));
    SB_LUT4 add_3370_5_lut (.I0(GND_net), .I1(n15397[2]), .I2(n431_adj_3789), 
            .I3(n37623), .O(n15112[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_8_lut (.I0(GND_net), .I1(n8446[5]), .I2(n536), 
            .I3(n37826), .O(n1804[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_25 (.CI(n36533), .I0(n9927[22]), .I1(GND_net), .CO(n36534));
    SB_CARRY mult_14_add_1219_8 (.CI(n37826), .I0(n8446[5]), .I1(n536), 
            .CO(n37827));
    SB_LUT4 add_3078_21_lut (.I0(GND_net), .I1(n8470[18]), .I2(GND_net), 
            .I3(n37535), .O(n8446[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_7_lut (.I0(GND_net), .I1(n8446[4]), .I2(n463_adj_3792), 
            .I3(n37825), .O(n1804[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n601));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3069_2 (.CI(GND_net), .I0(n53_adj_3785), .I1(n146_adj_3786), 
            .CO(n37427));
    SB_CARRY mult_14_add_1219_7 (.CI(n37825), .I0(n8446[4]), .I1(n463_adj_3792), 
            .CO(n37826));
    SB_CARRY add_3078_21 (.CI(n37535), .I0(n8470[18]), .I1(GND_net), .CO(n37536));
    SB_CARRY add_3370_5 (.CI(n37623), .I0(n15397[2]), .I1(n431_adj_3789), 
            .CO(n37624));
    SB_LUT4 add_3101_24_lut (.I0(GND_net), .I1(n9927[21]), .I2(GND_net), 
            .I3(n36532), .O(n9123[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_24 (.CI(n36532), .I0(n9927[21]), .I1(GND_net), .CO(n36533));
    SB_CARRY mult_14_add_1213_24 (.CI(n37704), .I0(n1799[21]), .I1(GND_net), 
            .CO(n1691));
    SB_LUT4 mult_14_add_1213_23_lut (.I0(GND_net), .I1(n1799[20]), .I2(GND_net), 
            .I3(n37703), .O(n1798[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_17_lut (.I0(GND_net), .I1(n8329[14]), .I2(GND_net), 
            .I3(n37426), .O(n8311[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_23 (.CI(n37703), .I0(n1799[20]), .I1(GND_net), 
            .CO(n37704));
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n698));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i158_2_lut (.I0(\Kd[2] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n234));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i158_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3059_19 (.CI(n37248), .I0(n8131[16]), .I1(GND_net), .CO(n37249));
    SB_LUT4 add_3370_4_lut (.I0(GND_net), .I1(n15397[1]), .I2(n334_adj_3793), 
            .I3(n37622), .O(n15112[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_23_lut (.I0(GND_net), .I1(n9927[20]), .I2(GND_net), 
            .I3(n36531), .O(n9123[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i148_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n219_adj_3502));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3078_20_lut (.I0(GND_net), .I1(n8470[17]), .I2(GND_net), 
            .I3(n37534), .O(n8446[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i15_1_lut (.I0(\PID_CONTROLLER.err[14] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[14]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_17_add_3_24 (.CI(n35985), .I0(GND_net), .I1(n79[22]), 
            .CO(n35986));
    SB_LUT4 add_3059_18_lut (.I0(GND_net), .I1(n8131[15]), .I2(GND_net), 
            .I3(n37247), .O(n8104[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_23 (.CI(n36531), .I0(n9927[20]), .I1(GND_net), .CO(n36532));
    SB_CARRY add_3059_18 (.CI(n37247), .I0(n8131[15]), .I1(GND_net), .CO(n37248));
    SB_LUT4 add_3101_22_lut (.I0(GND_net), .I1(n9927[19]), .I2(GND_net), 
            .I3(n36530), .O(n9123[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_22 (.CI(n36530), .I0(n9927[19]), .I1(GND_net), .CO(n36531));
    SB_LUT4 add_3101_21_lut (.I0(GND_net), .I1(n9927[18]), .I2(GND_net), 
            .I3(n36529), .O(n9123[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_21 (.CI(n36529), .I0(n9927[18]), .I1(GND_net), .CO(n36530));
    SB_LUT4 add_3101_20_lut (.I0(GND_net), .I1(n9927[17]), .I2(GND_net), 
            .I3(n36528), .O(n9123[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_20 (.CI(n36528), .I0(n9927[17]), .I1(GND_net), .CO(n36529));
    SB_LUT4 add_3101_19_lut (.I0(GND_net), .I1(n9927[16]), .I2(GND_net), 
            .I3(n36527), .O(n9123[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_4 (.CI(n37622), .I0(n15397[1]), .I1(n334_adj_3793), 
            .CO(n37623));
    SB_CARRY add_3101_19 (.CI(n36527), .I0(n9927[16]), .I1(GND_net), .CO(n36528));
    SB_LUT4 add_3068_16_lut (.I0(GND_net), .I1(n8329[13]), .I2(GND_net), 
            .I3(n37425), .O(n8311[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_17_lut (.I0(GND_net), .I1(n8131[14]), .I2(GND_net), 
            .I3(n37246), .O(n8104[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_18_lut (.I0(GND_net), .I1(n9927[15]), .I2(GND_net), 
            .I3(n36526), .O(n9123[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_33_lut (.I0(GND_net), .I1(n57[31]), .I2(n7059[0]), 
            .I3(n36224), .O(\PID_CONTROLLER.result_31__N_3003 [31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_18 (.CI(n36526), .I0(n9927[15]), .I1(GND_net), .CO(n36527));
    SB_LUT4 add_21902_32_lut (.I0(GND_net), .I1(n57[30]), .I2(n191[30]), 
            .I3(n36223), .O(\PID_CONTROLLER.result_31__N_3003 [30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_17_lut (.I0(GND_net), .I1(n9927[14]), .I2(GND_net), 
            .I3(n36525), .O(n9123[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n79[21]), 
            .I3(n35984), .O(pwm_23__N_2960[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[2]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3101_17 (.CI(n36525), .I0(n9927[14]), .I1(GND_net), .CO(n36526));
    SB_CARRY add_21902_32 (.CI(n36223), .I0(n57[30]), .I1(n191[30]), .CO(n36224));
    SB_LUT4 add_3101_16_lut (.I0(GND_net), .I1(n9927[13]), .I2(GND_net), 
            .I3(n36524), .O(n9123[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_16 (.CI(n36524), .I0(n9927[13]), .I1(GND_net), .CO(n36525));
    SB_CARRY add_3059_17 (.CI(n37246), .I0(n8131[14]), .I1(GND_net), .CO(n37247));
    SB_LUT4 add_21902_31_lut (.I0(GND_net), .I1(n57[29]), .I2(n191[29]), 
            .I3(n36222), .O(\PID_CONTROLLER.result_31__N_3003 [29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_15_lut (.I0(GND_net), .I1(n9927[12]), .I2(GND_net), 
            .I3(n36523), .O(n9123[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_31 (.CI(n36222), .I0(n57[29]), .I1(n191[29]), .CO(n36223));
    SB_LUT4 add_21902_30_lut (.I0(GND_net), .I1(n57[28]), .I2(n191[28]), 
            .I3(n36221), .O(\PID_CONTROLLER.result_31__N_3003 [28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_23 (.CI(n35984), .I0(GND_net), .I1(n79[21]), 
            .CO(n35985));
    SB_CARRY add_21902_30 (.CI(n36221), .I0(n57[28]), .I1(n191[28]), .CO(n36222));
    SB_LUT4 unary_minus_17_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n79[20]), 
            .I3(n35983), .O(\pwm_23__N_2960[20] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i75_2_lut (.I0(\Kd[1] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i213_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n316));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i213_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3101_15 (.CI(n36523), .I0(n9927[12]), .I1(GND_net), .CO(n36524));
    SB_LUT4 add_21902_29_lut (.I0(GND_net), .I1(n57[27]), .I2(n191[27]), 
            .I3(n36220), .O(\PID_CONTROLLER.result_31__N_3003 [27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_14_lut (.I0(GND_net), .I1(n9927[11]), .I2(GND_net), 
            .I3(n36522), .O(n9123[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_22 (.CI(n35983), .I0(GND_net), .I1(n79[20]), 
            .CO(n35984));
    SB_CARRY add_3101_14 (.CI(n36522), .I0(n9927[11]), .I1(GND_net), .CO(n36523));
    SB_LUT4 unary_minus_17_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n79[19]), 
            .I3(n35982), .O(pwm_23__N_2960[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_13_lut (.I0(GND_net), .I1(n9927[10]), .I2(GND_net), 
            .I3(n36521), .O(n9123[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_21 (.CI(n35982), .I0(GND_net), .I1(n79[19]), 
            .CO(n35983));
    SB_CARRY add_3101_13 (.CI(n36521), .I0(n9927[10]), .I1(GND_net), .CO(n36522));
    SB_CARRY add_21902_29 (.CI(n36220), .I0(n57[27]), .I1(n191[27]), .CO(n36221));
    SB_LUT4 add_3101_12_lut (.I0(GND_net), .I1(n9927[9]), .I2(GND_net), 
            .I3(n36520), .O(n9123[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_12 (.CI(n36520), .I0(n9927[9]), .I1(GND_net), .CO(n36521));
    SB_LUT4 add_3101_11_lut (.I0(GND_net), .I1(n9927[8]), .I2(GND_net), 
            .I3(n36519), .O(n9123[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i12_2_lut (.I0(\Kd[0] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i223_2_lut (.I0(\Kd[3] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n331));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_6_lut (.I0(GND_net), .I1(n8446[3]), .I2(n390), 
            .I3(n37824), .O(n1804[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_28_lut (.I0(GND_net), .I1(n57[26]), .I2(n191[26]), 
            .I3(n36219), .O(\PID_CONTROLLER.result_31__N_3003 [26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_11 (.CI(n36519), .I0(n9927[8]), .I1(GND_net), .CO(n36520));
    SB_LUT4 add_3101_10_lut (.I0(GND_net), .I1(n9927[7]), .I2(GND_net), 
            .I3(n36518), .O(n9123[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_28 (.CI(n36219), .I0(n57[26]), .I1(n191[26]), .CO(n36220));
    SB_CARRY add_3101_10 (.CI(n36518), .I0(n9927[7]), .I1(GND_net), .CO(n36519));
    SB_LUT4 add_3101_9_lut (.I0(GND_net), .I1(n9927[6]), .I2(GND_net), 
            .I3(n36517), .O(n9123[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_27_lut (.I0(GND_net), .I1(n57[25]), .I2(n191[25]), 
            .I3(n36218), .O(\PID_CONTROLLER.result_31__N_3003 [25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_9 (.CI(n36517), .I0(n9927[6]), .I1(GND_net), .CO(n36518));
    SB_LUT4 add_3059_16_lut (.I0(GND_net), .I1(n8131[13]), .I2(GND_net), 
            .I3(n37245), .O(n8104[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_8_lut (.I0(GND_net), .I1(n9927[5]), .I2(n689_adj_3797), 
            .I3(n36516), .O(n9123[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i140_2_lut (.I0(\Kd[2] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n207));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i288_2_lut (.I0(\Kd[4] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n428));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i288_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_21902_27 (.CI(n36218), .I0(n57[25]), .I1(n191[25]), .CO(n36219));
    SB_CARRY add_3101_8 (.CI(n36516), .I0(n9927[5]), .I1(n689_adj_3797), 
            .CO(n36517));
    SB_LUT4 add_3101_7_lut (.I0(GND_net), .I1(n9927[4]), .I2(n592_adj_3798), 
            .I3(n36515), .O(n9123[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_26_lut (.I0(GND_net), .I1(n57[24]), .I2(n191[24]), 
            .I3(n36217), .O(\PID_CONTROLLER.result_31__N_3003 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_7 (.CI(n36515), .I0(n9927[4]), .I1(n592_adj_3798), 
            .CO(n36516));
    SB_LUT4 mult_14_add_1213_22_lut (.I0(GND_net), .I1(n1799[19]), .I2(GND_net), 
            .I3(n37702), .O(n1798[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_3_lut (.I0(GND_net), .I1(n15397[0]), .I2(n237_adj_3799), 
            .I3(n37621), .O(n15112[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i278_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n413_adj_3500));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i278_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1219_6 (.CI(n37824), .I0(n8446[3]), .I1(n390), 
            .CO(n37825));
    SB_LUT4 unary_minus_17_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n79[18]), 
            .I3(n35981), .O(pwm_23__N_2960[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_20 (.CI(n35981), .I0(GND_net), .I1(n79[18]), 
            .CO(n35982));
    SB_LUT4 add_3101_6_lut (.I0(GND_net), .I1(n9927[3]), .I2(n495_adj_3801), 
            .I3(n36514), .O(n9123[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i113_2_lut (.I0(\Kd[1] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n167));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i50_2_lut (.I0(\Kd[0] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i347_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3101_6 (.CI(n36514), .I0(n9927[3]), .I1(n495_adj_3801), 
            .CO(n36515));
    SB_CARRY add_21902_26 (.CI(n36217), .I0(n57[24]), .I1(n191[24]), .CO(n36218));
    SB_LUT4 add_3101_5_lut (.I0(GND_net), .I1(n9927[2]), .I2(n398_adj_3802), 
            .I3(n36513), .O(n9123[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_5 (.CI(n36513), .I0(n9927[2]), .I1(n398_adj_3802), 
            .CO(n36514));
    SB_LUT4 add_21902_25_lut (.I0(GND_net), .I1(n57[23]), .I2(n191[23]), 
            .I3(n36216), .O(\PID_CONTROLLER.result_31__N_3003 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_4_lut (.I0(GND_net), .I1(n9927[1]), .I2(n301_adj_3803), 
            .I3(n36512), .O(n9123[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_20 (.CI(n37534), .I0(n8470[17]), .I1(GND_net), .CO(n37535));
    SB_LUT4 sub_11_inv_0_i16_1_lut (.I0(\PID_CONTROLLER.err[15] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[15]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[3]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i343_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n510_adj_3498));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i343_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3101_4 (.CI(n36512), .I0(n9927[1]), .I1(n301_adj_3803), 
            .CO(n36513));
    SB_CARRY add_21902_25 (.CI(n36216), .I0(n57[23]), .I1(n191[23]), .CO(n36217));
    SB_LUT4 unary_minus_17_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n79[17]), 
            .I3(n35980), .O(pwm_23__N_2960[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_16 (.CI(n37425), .I0(n8329[13]), .I1(GND_net), .CO(n37426));
    SB_CARRY add_3059_16 (.CI(n37245), .I0(n8131[13]), .I1(GND_net), .CO(n37246));
    SB_LUT4 add_3101_3_lut (.I0(GND_net), .I1(n9927[0]), .I2(n204_adj_3805), 
            .I3(n36511), .O(n9123[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_24_lut (.I0(GND_net), .I1(n57[22]), .I2(n191[22]), 
            .I3(n36215), .O(\PID_CONTROLLER.result_31__N_3003 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_3 (.CI(n36511), .I0(n9927[0]), .I1(n204_adj_3805), 
            .CO(n36512));
    SB_CARRY add_21902_24 (.CI(n36215), .I0(n57[22]), .I1(n191[22]), .CO(n36216));
    SB_CARRY unary_minus_17_add_3_19 (.CI(n35980), .I0(GND_net), .I1(n79[17]), 
            .CO(n35981));
    SB_LUT4 add_3101_2_lut (.I0(GND_net), .I1(n14_adj_3806), .I2(n107_adj_3807), 
            .I3(GND_net), .O(n9123[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n79[16]), 
            .I3(n35979), .O(pwm_23__N_2960[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_2 (.CI(GND_net), .I0(n14_adj_3806), .I1(n107_adj_3807), 
            .CO(n36511));
    SB_LUT4 add_21902_23_lut (.I0(GND_net), .I1(n57[21]), .I2(n191[21]), 
            .I3(n36214), .O(\PID_CONTROLLER.result_31__N_3003 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3299_14_lut (.I0(GND_net), .I1(n14166[11]), .I2(GND_net), 
            .I3(n36510), .O(n13732[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_18 (.CI(n35979), .I0(GND_net), .I1(n79[16]), 
            .CO(n35980));
    SB_LUT4 unary_minus_17_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n79[15]), 
            .I3(n35978), .O(pwm_23__N_2960[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[4]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i205_2_lut (.I0(\Kd[3] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n304));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i353_2_lut (.I0(\Kd[5] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n525));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3299_13_lut (.I0(GND_net), .I1(n14166[10]), .I2(GND_net), 
            .I3(n36509), .O(n13732[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_23 (.CI(n36214), .I0(n57[21]), .I1(n191[21]), .CO(n36215));
    SB_CARRY add_3299_13 (.CI(n36509), .I0(n14166[10]), .I1(GND_net), 
            .CO(n36510));
    SB_LUT4 add_21902_22_lut (.I0(GND_net), .I1(n57[20]), .I2(n191[20]), 
            .I3(n36213), .O(\PID_CONTROLLER.result_31__N_3003 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3299_12_lut (.I0(GND_net), .I1(n14166[9]), .I2(GND_net), 
            .I3(n36508), .O(n13732[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3299_12 (.CI(n36508), .I0(n14166[9]), .I1(GND_net), .CO(n36509));
    SB_LUT4 add_3059_15_lut (.I0(GND_net), .I1(n8131[12]), .I2(GND_net), 
            .I3(n37244), .O(n8104[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_15 (.CI(n37244), .I0(n8131[12]), .I1(GND_net), .CO(n37245));
    SB_LUT4 add_3299_11_lut (.I0(GND_net), .I1(n14166[8]), .I2(GND_net), 
            .I3(n36507), .O(n13732[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i270_2_lut (.I0(\Kd[4] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n401));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1219_5_lut (.I0(GND_net), .I1(n8446[2]), .I2(n317), 
            .I3(n37823), .O(n1804[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3299_11 (.CI(n36507), .I0(n14166[8]), .I1(GND_net), .CO(n36508));
    SB_CARRY mult_14_add_1213_22 (.CI(n37702), .I0(n1799[19]), .I1(GND_net), 
            .CO(n37703));
    SB_CARRY add_21902_22 (.CI(n36213), .I0(n57[20]), .I1(n191[20]), .CO(n36214));
    SB_LUT4 mult_14_add_1213_21_lut (.I0(GND_net), .I1(n1799[18]), .I2(GND_net), 
            .I3(n37701), .O(n1798[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3299_10_lut (.I0(GND_net), .I1(n14166[7]), .I2(GND_net), 
            .I3(n36506), .O(n13732[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_21 (.CI(n37701), .I0(n1799[18]), .I1(GND_net), 
            .CO(n37702));
    SB_CARRY add_3299_10 (.CI(n36506), .I0(n14166[7]), .I1(GND_net), .CO(n36507));
    SB_LUT4 add_3068_15_lut (.I0(GND_net), .I1(n8329[12]), .I2(GND_net), 
            .I3(n37424), .O(n8311[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_21_lut (.I0(GND_net), .I1(n57[19]), .I2(n191[19]), 
            .I3(n36212), .O(\PID_CONTROLLER.result_31__N_3003 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3299_9_lut (.I0(GND_net), .I1(n14166[6]), .I2(GND_net), 
            .I3(n36505), .O(n13732[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_5 (.CI(n37823), .I0(n8446[2]), .I1(n317), 
            .CO(n37824));
    SB_LUT4 add_3059_14_lut (.I0(GND_net), .I1(n8131[11]), .I2(GND_net), 
            .I3(n37243), .O(n8104[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_21 (.CI(n36212), .I0(n57[19]), .I1(n191[19]), .CO(n36213));
    SB_LUT4 mult_14_add_1219_4_lut (.I0(GND_net), .I1(n8446[1]), .I2(n244_adj_3811), 
            .I3(n37822), .O(n1804[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_15 (.CI(n37424), .I0(n8329[12]), .I1(GND_net), .CO(n37425));
    SB_LUT4 add_21902_20_lut (.I0(GND_net), .I1(n57[18]), .I2(n191[18]), 
            .I3(n36211), .O(\PID_CONTROLLER.result_31__N_3003 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_14 (.CI(n37243), .I0(n8131[11]), .I1(GND_net), .CO(n37244));
    SB_LUT4 add_3059_13_lut (.I0(GND_net), .I1(n8131[10]), .I2(GND_net), 
            .I3(n37242), .O(n8104[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_13 (.CI(n37242), .I0(n8131[10]), .I1(GND_net), .CO(n37243));
    SB_CARRY add_3299_9 (.CI(n36505), .I0(n14166[6]), .I1(GND_net), .CO(n36506));
    SB_CARRY add_21902_20 (.CI(n36211), .I0(n57[18]), .I1(n191[18]), .CO(n36212));
    SB_LUT4 mult_14_add_1213_20_lut (.I0(GND_net), .I1(n1799[17]), .I2(GND_net), 
            .I3(n37700), .O(n1798[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_3 (.CI(n37621), .I0(n15397[0]), .I1(n237_adj_3799), 
            .CO(n37622));
    SB_LUT4 mult_12_i418_2_lut (.I0(\Kd[6] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n622));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i178_2_lut (.I0(\Kd[2] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n264));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3078_19_lut (.I0(GND_net), .I1(n8470[16]), .I2(GND_net), 
            .I3(n37533), .O(n8446[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3299_8_lut (.I0(GND_net), .I1(n14166[5]), .I2(n545), .I3(n36504), 
            .O(n13732[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_19_lut (.I0(GND_net), .I1(n57[17]), .I2(n191[17]), 
            .I3(n36210), .O(\PID_CONTROLLER.result_31__N_3003 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3299_8 (.CI(n36504), .I0(n14166[5]), .I1(n545), .CO(n36505));
    SB_LUT4 add_3299_7_lut (.I0(GND_net), .I1(n14166[4]), .I2(n472), .I3(n36503), 
            .O(n13732[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_19 (.CI(n36210), .I0(n57[17]), .I1(n191[17]), .CO(n36211));
    SB_CARRY add_3299_7 (.CI(n36503), .I0(n14166[4]), .I1(n472), .CO(n36504));
    SB_LUT4 mult_12_i335_2_lut (.I0(\Kd[5] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n498));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[5]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i483_2_lut (.I0(\Kd[7] ), .I1(n69[13]), .I2(GND_net), 
            .I3(GND_net), .O(n719));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3299_6_lut (.I0(GND_net), .I1(n14166[3]), .I2(n399_c), 
            .I3(n36502), .O(n13732[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_18_lut (.I0(GND_net), .I1(n57[16]), .I2(n191[16]), 
            .I3(n36209), .O(\PID_CONTROLLER.result_31__N_3003 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3299_6 (.CI(n36502), .I0(n14166[3]), .I1(n399_c), .CO(n36503));
    SB_LUT4 mult_12_i400_2_lut (.I0(\Kd[6] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n595));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i243_2_lut (.I0(\Kd[3] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n361));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i465_2_lut (.I0(\Kd[7] ), .I1(n69[4]), .I2(GND_net), 
            .I3(GND_net), .O(n692));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i308_2_lut (.I0(\Kd[4] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n458));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3299_5_lut (.I0(GND_net), .I1(n14166[2]), .I2(n326), .I3(n36501), 
            .O(n13732[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_18 (.CI(n36209), .I0(n57[16]), .I1(n191[16]), .CO(n36210));
    SB_LUT4 add_3059_12_lut (.I0(GND_net), .I1(n8131[9]), .I2(GND_net), 
            .I3(n37241), .O(n8104[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3299_5 (.CI(n36501), .I0(n14166[2]), .I1(n326), .CO(n36502));
    SB_LUT4 add_21902_17_lut (.I0(GND_net), .I1(n57[15]), .I2(n191[15]), 
            .I3(n36208), .O(\PID_CONTROLLER.result_31__N_3003 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3299_4_lut (.I0(GND_net), .I1(n14166[1]), .I2(n253), .I3(n36500), 
            .O(n13732[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_17 (.CI(n36208), .I0(n57[15]), .I1(n191[15]), .CO(n36209));
    SB_CARRY add_3299_4 (.CI(n36500), .I0(n14166[1]), .I1(n253), .CO(n36501));
    SB_CARRY unary_minus_17_add_3_17 (.CI(n35978), .I0(GND_net), .I1(n79[15]), 
            .CO(n35979));
    SB_LUT4 add_3068_14_lut (.I0(GND_net), .I1(n8329[11]), .I2(GND_net), 
            .I3(n37423), .O(n8311[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_16_lut (.I0(GND_net), .I1(n57[14]), .I2(n191[14]), 
            .I3(n36207), .O(\PID_CONTROLLER.result_31__N_3003 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3299_3_lut (.I0(GND_net), .I1(n14166[0]), .I2(n180), .I3(n36499), 
            .O(n13732[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i17_1_lut (.I0(\PID_CONTROLLER.err[16] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[16]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i373_2_lut (.I0(\Kd[5] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n555));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i438_2_lut (.I0(\Kd[6] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n652));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n79[14]), 
            .I3(n35977), .O(\pwm_23__N_2960[14] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3299_3 (.CI(n36499), .I0(n14166[0]), .I1(n180), .CO(n36500));
    SB_LUT4 add_3299_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n13732[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3299_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_20 (.CI(n37700), .I0(n1799[17]), .I1(GND_net), 
            .CO(n37701));
    SB_CARRY add_3078_19 (.CI(n37533), .I0(n8470[16]), .I1(GND_net), .CO(n37534));
    SB_CARRY add_3299_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n36499));
    SB_CARRY add_21902_16 (.CI(n36207), .I0(n57[14]), .I1(n191[14]), .CO(n36208));
    SB_LUT4 mult_14_add_1213_19_lut (.I0(GND_net), .I1(n1799[16]), .I2(GND_net), 
            .I3(n37699), .O(n1798[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_28_lut (.I0(GND_net), .I1(n10669[25]), .I2(GND_net), 
            .I3(n36498), .O(n9927[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_2_lut (.I0(GND_net), .I1(n47_adj_3813), .I2(n140_adj_3814), 
            .I3(GND_net), .O(n15112[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_16 (.CI(n35977), .I0(GND_net), .I1(n79[14]), 
            .CO(n35978));
    SB_LUT4 mult_12_i503_2_lut (.I0(\Kd[7] ), .I1(n69[23]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i115_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n182));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n79[13]), 
            .I3(n35976), .O(\pwm_23__N_2960[13] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_15 (.CI(n35976), .I0(GND_net), .I1(n79[13]), 
            .CO(n35977));
    SB_LUT4 add_3140_27_lut (.I0(GND_net), .I1(n10669[24]), .I2(GND_net), 
            .I3(n36497), .O(n9927[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_27 (.CI(n36497), .I0(n10669[24]), .I1(GND_net), 
            .CO(n36498));
    SB_CARRY add_3068_14 (.CI(n37423), .I0(n8329[11]), .I1(GND_net), .CO(n37424));
    SB_LUT4 add_3140_26_lut (.I0(GND_net), .I1(n10669[23]), .I2(GND_net), 
            .I3(n36496), .O(n9927[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i115_2_lut (.I0(\Kd[1] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n170));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i52_2_lut (.I0(\Kd[0] ), .I1(n69[25]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i52_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i180_2_lut (.I0(\Kd[2] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n267));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i95_2_lut (.I0(\Kd[1] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n140));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i95_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3059_12 (.CI(n37241), .I0(n8131[9]), .I1(GND_net), .CO(n37242));
    SB_LUT4 add_3078_18_lut (.I0(GND_net), .I1(n8470[15]), .I2(GND_net), 
            .I3(n37532), .O(n8446[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_15_lut (.I0(GND_net), .I1(n57[13]), .I2(n191[13]), 
            .I3(n36206), .O(\PID_CONTROLLER.result_31__N_3003 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i32_2_lut (.I0(\Kd[0] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_3388));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1219_4 (.CI(n37822), .I0(n8446[1]), .I1(n244_adj_3811), 
            .CO(n37823));
    SB_CARRY add_21902_15 (.CI(n36206), .I0(n57[13]), .I1(n191[13]), .CO(n36207));
    SB_CARRY add_3140_26 (.CI(n36496), .I0(n10669[23]), .I1(GND_net), 
            .CO(n36497));
    SB_LUT4 mult_12_i245_2_lut (.I0(\Kd[3] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n364));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i160_2_lut (.I0(\Kd[2] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n237));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i310_2_lut (.I0(\Kd[4] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n461_adj_3387));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i225_2_lut (.I0(\Kd[3] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n334));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i375_2_lut (.I0(\Kd[5] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n558_adj_3386));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n79[12]), 
            .I3(n35975), .O(pwm_23__N_2960[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_25_lut (.I0(GND_net), .I1(n10669[22]), .I2(GND_net), 
            .I3(n36495), .O(n9927[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_14_lut (.I0(GND_net), .I1(n57[12]), .I2(n191[12]), 
            .I3(n36205), .O(\PID_CONTROLLER.result_31__N_3003 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i67_2_lut (.I0(\Kd[1] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i290_2_lut (.I0(\Kd[4] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n431));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i440_2_lut (.I0(\Kd[6] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n655));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i440_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i505_2_lut (.I0(\Kd[7] ), .I1(n69[24]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i355_2_lut (.I0(\Kd[5] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n528));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i95_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i46_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i77_2_lut (.I0(\Kd[1] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i77_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_17_add_3_14 (.CI(n35975), .I0(GND_net), .I1(n79[12]), 
            .CO(n35976));
    SB_LUT4 unary_minus_17_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n79[11]), 
            .I3(n35974), .O(pwm_23__N_2960[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i14_2_lut (.I0(\Kd[0] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_3384));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i420_2_lut (.I0(\Kd[6] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n625));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i142_2_lut (.I0(\Kd[2] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n210));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i207_2_lut (.I0(\Kd[3] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n307));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i485_2_lut (.I0(\Kd[7] ), .I1(n69[14]), .I2(GND_net), 
            .I3(GND_net), .O(n722));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i50_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3389));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i180_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n276));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i245_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n370));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22112_3_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n35561), .I2(n37873), 
            .I3(GND_net), .O(n16635[1]));   // verilog/motorControl.v(43[17:23])
    defparam i22112_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n464));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n558));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i442_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i4_2_lut (.I0(\Kd[0] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_3496));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i4_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3370_2 (.CI(GND_net), .I0(n47_adj_3813), .I1(n140_adj_3814), 
            .CO(n37621));
    SB_CARRY add_3078_18 (.CI(n37532), .I0(n8470[15]), .I1(GND_net), .CO(n37533));
    SB_LUT4 add_3479_9_lut (.I0(GND_net), .I1(n16618[6]), .I2(GND_net), 
            .I3(n37620), .O(n16569[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_13_lut (.I0(GND_net), .I1(n8329[10]), .I2(GND_net), 
            .I3(n37422), .O(n8311[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_11_lut (.I0(GND_net), .I1(n8131[8]), .I2(GND_net), 
            .I3(n37240), .O(n8104[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_3_lut (.I0(GND_net), .I1(n8446[0]), .I2(n171_adj_3819), 
            .I3(n37821), .O(n1804[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_14 (.CI(n36205), .I0(n57[12]), .I1(n191[12]), .CO(n36206));
    SB_CARRY unary_minus_17_add_3_13 (.CI(n35974), .I0(GND_net), .I1(n79[11]), 
            .CO(n35975));
    SB_CARRY mult_14_add_1219_3 (.CI(n37821), .I0(n8446[0]), .I1(n171_adj_3819), 
            .CO(n37822));
    SB_LUT4 add_21902_13_lut (.I0(GND_net), .I1(n57[11]), .I2(n191[11]), 
            .I3(n36204), .O(\PID_CONTROLLER.result_31__N_3003 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_17_lut (.I0(GND_net), .I1(n8470[14]), .I2(GND_net), 
            .I3(n37531), .O(n8446[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_13 (.CI(n37422), .I0(n8329[10]), .I1(GND_net), .CO(n37423));
    SB_CARRY add_3059_11 (.CI(n37240), .I0(n8131[8]), .I1(GND_net), .CO(n37241));
    SB_LUT4 add_3059_10_lut (.I0(GND_net), .I1(n8131[7]), .I2(GND_net), 
            .I3(n37239), .O(n8104[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_12_lut (.I0(GND_net), .I1(n8329[9]), .I2(GND_net), 
            .I3(n37421), .O(n8311[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_10 (.CI(n37239), .I0(n8131[7]), .I1(GND_net), .CO(n37240));
    SB_CARRY add_3078_17 (.CI(n37531), .I0(n8470[14]), .I1(GND_net), .CO(n37532));
    SB_CARRY add_3140_25 (.CI(n36495), .I0(n10669[22]), .I1(GND_net), 
            .CO(n36496));
    SB_CARRY add_21902_13 (.CI(n36204), .I0(n57[11]), .I1(n191[11]), .CO(n36205));
    SB_LUT4 mult_14_add_1219_2_lut (.I0(GND_net), .I1(n35), .I2(n98_adj_3820), 
            .I3(GND_net), .O(n1804[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_24_lut (.I0(GND_net), .I1(n10669[21]), .I2(GND_net), 
            .I3(n36494), .O(n9927[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_12_lut (.I0(GND_net), .I1(n57[10]), .I2(n191[10]), 
            .I3(n36203), .O(\PID_CONTROLLER.result_31__N_3003 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_24 (.CI(n36494), .I0(n10669[21]), .I1(GND_net), 
            .CO(n36495));
    SB_CARRY add_21902_12 (.CI(n36203), .I0(n57[10]), .I1(n191[10]), .CO(n36204));
    SB_LUT4 add_21902_11_lut (.I0(GND_net), .I1(n57[9]), .I2(n191[9]), 
            .I3(n36202), .O(\PID_CONTROLLER.result_31__N_3003 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_23_lut (.I0(GND_net), .I1(n10669[20]), .I2(GND_net), 
            .I3(n36493), .O(n9927[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_11 (.CI(n36202), .I0(n57[9]), .I1(n191[9]), .CO(n36203));
    SB_LUT4 unary_minus_17_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n79[10]), 
            .I3(n35973), .O(pwm_23__N_2960[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut (.I0(n35561), .I1(n7_adj_3822), .I2(n8_adj_3823), 
            .I3(n8_adj_3824), .O(n43968));   // verilog/motorControl.v(43[17:23])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3140_23 (.CI(n36493), .I0(n10669[20]), .I1(GND_net), 
            .CO(n36494));
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n607));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1219_2 (.CI(GND_net), .I0(n35), .I1(n98_adj_3820), 
            .CO(n37821));
    SB_LUT4 mult_14_add_1218_24_lut (.I0(GND_net), .I1(n1804[21]), .I2(GND_net), 
            .I3(n37819), .O(n1803[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_24 (.CI(n37819), .I0(n1804[21]), .I1(GND_net), 
            .CO(n1711));
    SB_CARRY mult_14_add_1213_19 (.CI(n37699), .I0(n1799[16]), .I1(GND_net), 
            .CO(n37700));
    SB_LUT4 add_3479_8_lut (.I0(GND_net), .I1(n16618[5]), .I2(n749_adj_3825), 
            .I3(n37619), .O(n16569[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_23_lut (.I0(GND_net), .I1(n1804[20]), .I2(GND_net), 
            .I3(n37818), .O(n1803[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_23 (.CI(n37818), .I0(n1804[20]), .I1(GND_net), 
            .CO(n37819));
    SB_LUT4 add_3078_16_lut (.I0(GND_net), .I1(n8470[13]), .I2(GND_net), 
            .I3(n37530), .O(n8446[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_10_lut (.I0(GND_net), .I1(n57[8]), .I2(n191[8]), 
            .I3(n36201), .O(\PID_CONTROLLER.result_31__N_3003 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_22_lut (.I0(GND_net), .I1(n10669[19]), .I2(GND_net), 
            .I3(n36492), .O(n9927[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_10 (.CI(n36201), .I0(n57[8]), .I1(n191[8]), .CO(n36202));
    SB_LUT4 add_3059_9_lut (.I0(GND_net), .I1(n8131[6]), .I2(GND_net), 
            .I3(n37238), .O(n8104[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i473_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n704));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i473_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3068_12 (.CI(n37421), .I0(n8329[9]), .I1(GND_net), .CO(n37422));
    SB_LUT4 sub_11_inv_0_i18_1_lut (.I0(\PID_CONTROLLER.err[17] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[17]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3479_8 (.CI(n37619), .I0(n16618[5]), .I1(n749_adj_3825), 
            .CO(n37620));
    SB_LUT4 mult_14_add_1213_18_lut (.I0(GND_net), .I1(n1799[15]), .I2(GND_net), 
            .I3(n37698), .O(n1798[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_18 (.CI(n37698), .I0(n1799[15]), .I1(GND_net), 
            .CO(n37699));
    SB_LUT4 unary_minus_21_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[6]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1218_22_lut (.I0(GND_net), .I1(n1804[19]), .I2(GND_net), 
            .I3(n37817), .O(n1803[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_22 (.CI(n37817), .I0(n1804[19]), .I1(GND_net), 
            .CO(n37818));
    SB_LUT4 mult_14_add_1218_21_lut (.I0(GND_net), .I1(n1804[18]), .I2(GND_net), 
            .I3(n37816), .O(n1803[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_21 (.CI(n37816), .I0(n1804[18]), .I1(GND_net), 
            .CO(n37817));
    SB_LUT4 mult_14_add_1218_20_lut (.I0(GND_net), .I1(n1804[17]), .I2(GND_net), 
            .I3(n37815), .O(n1803[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_20 (.CI(n37815), .I0(n1804[17]), .I1(GND_net), 
            .CO(n37816));
    SB_LUT4 mult_14_add_1218_19_lut (.I0(GND_net), .I1(n1804[16]), .I2(GND_net), 
            .I3(n37814), .O(n1803[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_19 (.CI(n37814), .I0(n1804[16]), .I1(GND_net), 
            .CO(n37815));
    SB_LUT4 add_3479_7_lut (.I0(GND_net), .I1(n16618[4]), .I2(n652_adj_3826), 
            .I3(n37618), .O(n16569[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i132_2_lut (.I0(\Kd[2] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1213_17_lut (.I0(GND_net), .I1(n1799[14]), .I2(GND_net), 
            .I3(n37697), .O(n1798[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3479_7 (.CI(n37618), .I0(n16618[4]), .I1(n652_adj_3826), 
            .CO(n37619));
    SB_LUT4 mult_14_add_1218_18_lut (.I0(GND_net), .I1(n1804[15]), .I2(GND_net), 
            .I3(n37813), .O(n1803[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_17 (.CI(n37697), .I0(n1799[14]), .I1(GND_net), 
            .CO(n37698));
    SB_CARRY mult_14_add_1218_18 (.CI(n37813), .I0(n1804[15]), .I1(GND_net), 
            .CO(n37814));
    SB_LUT4 mult_14_add_1218_17_lut (.I0(GND_net), .I1(n1804[14]), .I2(GND_net), 
            .I3(n37812), .O(n1803[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_9 (.CI(n37238), .I0(n8131[6]), .I1(GND_net), .CO(n37239));
    SB_LUT4 mult_14_add_1213_16_lut (.I0(GND_net), .I1(n1799[13]), .I2(GND_net), 
            .I3(n37696), .O(n1798[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_11_lut (.I0(GND_net), .I1(n8329[8]), .I2(GND_net), 
            .I3(n37420), .O(n8311[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_8_lut (.I0(GND_net), .I1(n8131[5]), .I2(n698_adj_3827), 
            .I3(n37237), .O(n8104[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3479_6_lut (.I0(GND_net), .I1(n16618[3]), .I2(n555_adj_3828), 
            .I3(n37617), .O(n16569[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_16 (.CI(n37530), .I0(n8470[13]), .I1(GND_net), .CO(n37531));
    SB_CARRY add_3068_11 (.CI(n37420), .I0(n8329[8]), .I1(GND_net), .CO(n37421));
    SB_CARRY mult_14_add_1213_16 (.CI(n37696), .I0(n1799[13]), .I1(GND_net), 
            .CO(n37697));
    SB_CARRY add_3059_8 (.CI(n37237), .I0(n8131[5]), .I1(n698_adj_3827), 
            .CO(n37238));
    SB_CARRY unary_minus_17_add_3_12 (.CI(n35973), .I0(GND_net), .I1(n79[10]), 
            .CO(n35974));
    SB_LUT4 add_3068_10_lut (.I0(GND_net), .I1(n8329[7]), .I2(GND_net), 
            .I3(n37419), .O(n8311[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_9_lut (.I0(GND_net), .I1(n57[7]), .I2(n191[7]), 
            .I3(n36200), .O(\PID_CONTROLLER.result_31__N_3003 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_7_lut (.I0(GND_net), .I1(n8131[4]), .I2(n601_adj_3829), 
            .I3(n37236), .O(n8104[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3479_6 (.CI(n37617), .I0(n16618[3]), .I1(n555_adj_3828), 
            .CO(n37618));
    SB_CARRY add_3140_22 (.CI(n36492), .I0(n10669[19]), .I1(GND_net), 
            .CO(n36493));
    SB_LUT4 unary_minus_17_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n79[9]), 
            .I3(n35972), .O(pwm_23__N_2960[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_21_lut (.I0(GND_net), .I1(n10669[18]), .I2(GND_net), 
            .I3(n36491), .O(n9927[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_11 (.CI(n35972), .I0(GND_net), .I1(n79[9]), 
            .CO(n35973));
    SB_CARRY add_3140_21 (.CI(n36491), .I0(n10669[18]), .I1(GND_net), 
            .CO(n36492));
    SB_CARRY mult_14_add_1218_17 (.CI(n37812), .I0(n1804[14]), .I1(GND_net), 
            .CO(n37813));
    SB_LUT4 add_3140_20_lut (.I0(GND_net), .I1(n10669[17]), .I2(GND_net), 
            .I3(n36490), .O(n9927[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_9 (.CI(n36200), .I0(n57[7]), .I1(n191[7]), .CO(n36201));
    SB_LUT4 add_3479_5_lut (.I0(GND_net), .I1(n16618[2]), .I2(n458_adj_3831), 
            .I3(n37616), .O(n16569[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3479_5 (.CI(n37616), .I0(n16618[2]), .I1(n458_adj_3831), 
            .CO(n37617));
    SB_CARRY add_3140_20 (.CI(n36490), .I0(n10669[17]), .I1(GND_net), 
            .CO(n36491));
    SB_LUT4 unary_minus_17_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n79[8]), 
            .I3(n35971), .O(pwm_23__N_2960[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3479_4_lut (.I0(GND_net), .I1(n16618[1]), .I2(n361_adj_3833), 
            .I3(n37615), .O(n16569[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_10 (.CI(n35971), .I0(GND_net), .I1(n79[8]), 
            .CO(n35972));
    SB_LUT4 sub_11_inv_0_i19_1_lut (.I0(\PID_CONTROLLER.err[18] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[18]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1213_15_lut (.I0(GND_net), .I1(n1799[12]), .I2(GND_net), 
            .I3(n37695), .O(n1798[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_19_lut (.I0(GND_net), .I1(n10669[16]), .I2(GND_net), 
            .I3(n36489), .O(n9927[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i20_1_lut (.I0(\PID_CONTROLLER.err[19] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[19]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3140_19 (.CI(n36489), .I0(n10669[16]), .I1(GND_net), 
            .CO(n36490));
    SB_LUT4 mult_12_i197_2_lut (.I0(\Kd[3] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n292));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_21902_8_lut (.I0(GND_net), .I1(n57[6]), .I2(n191[6]), 
            .I3(n36199), .O(\PID_CONTROLLER.result_31__N_3003 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[7]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i21_1_lut (.I0(\PID_CONTROLLER.err[20] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[20]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21902_8 (.CI(n36199), .I0(n57[6]), .I1(n191[6]), .CO(n36200));
    SB_CARRY mult_14_add_1213_15 (.CI(n37695), .I0(n1799[12]), .I1(GND_net), 
            .CO(n37696));
    SB_LUT4 mult_14_i144_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3140_18_lut (.I0(GND_net), .I1(n10669[15]), .I2(GND_net), 
            .I3(n36488), .O(n9927[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3479_4 (.CI(n37615), .I0(n16618[1]), .I1(n361_adj_3833), 
            .CO(n37616));
    SB_CARRY add_3140_18 (.CI(n36488), .I0(n10669[15]), .I1(GND_net), 
            .CO(n36489));
    SB_LUT4 mult_14_add_1213_14_lut (.I0(GND_net), .I1(n1799[11]), .I2(GND_net), 
            .I3(n37694), .O(n1798[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_7 (.CI(n37236), .I0(n8131[4]), .I1(n601_adj_3829), 
            .CO(n37237));
    SB_LUT4 add_3078_15_lut (.I0(GND_net), .I1(n8470[12]), .I2(GND_net), 
            .I3(n37529), .O(n8446[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_17_lut (.I0(GND_net), .I1(n10669[14]), .I2(GND_net), 
            .I3(n36487), .O(n9927[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3078_15 (.CI(n37529), .I0(n8470[12]), .I1(GND_net), .CO(n37530));
    SB_LUT4 add_21902_7_lut (.I0(GND_net), .I1(n57[5]), .I2(n191[5]), 
            .I3(n36198), .O(\PID_CONTROLLER.result_31__N_3003 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_16_lut (.I0(GND_net), .I1(n1804[13]), .I2(GND_net), 
            .I3(n37811), .O(n1803[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_17 (.CI(n36487), .I0(n10669[14]), .I1(GND_net), 
            .CO(n36488));
    SB_CARRY add_21902_7 (.CI(n36198), .I0(n57[5]), .I1(n191[5]), .CO(n36199));
    SB_CARRY add_3068_10 (.CI(n37419), .I0(n8329[7]), .I1(GND_net), .CO(n37420));
    SB_LUT4 unary_minus_17_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n79[7]), 
            .I3(n35970), .O(pwm_23__N_2960[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_9 (.CI(n35970), .I0(GND_net), .I1(n79[7]), 
            .CO(n35971));
    SB_LUT4 add_3140_16_lut (.I0(GND_net), .I1(n10669[13]), .I2(GND_net), 
            .I3(n36486), .O(n9927[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_16 (.CI(n36486), .I0(n10669[13]), .I1(GND_net), 
            .CO(n36487));
    SB_LUT4 add_3140_15_lut (.I0(GND_net), .I1(n10669[12]), .I2(GND_net), 
            .I3(n36485), .O(n9927[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_14 (.CI(n37694), .I0(n1799[11]), .I1(GND_net), 
            .CO(n37695));
    SB_LUT4 unary_minus_21_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[8]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i262_2_lut (.I0(\Kd[4] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n389));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i262_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1218_16 (.CI(n37811), .I0(n1804[13]), .I1(GND_net), 
            .CO(n37812));
    SB_LUT4 mult_12_i272_2_lut (.I0(\Kd[4] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n404));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3059_6_lut (.I0(GND_net), .I1(n8131[3]), .I2(n504_adj_3835), 
            .I3(n37235), .O(n8104[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_6 (.CI(n37235), .I0(n8131[3]), .I1(n504_adj_3835), 
            .CO(n37236));
    SB_LUT4 add_3059_5_lut (.I0(GND_net), .I1(n8131[2]), .I2(n407_adj_3836), 
            .I3(n37234), .O(n8104[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_15 (.CI(n36485), .I0(n10669[12]), .I1(GND_net), 
            .CO(n36486));
    SB_LUT4 add_3140_14_lut (.I0(GND_net), .I1(n10669[11]), .I2(GND_net), 
            .I3(n36484), .O(n9927[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_6_lut (.I0(GND_net), .I1(n57[4]), .I2(n191[4]), 
            .I3(n36197), .O(\PID_CONTROLLER.result_31__N_3003 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3479_3_lut (.I0(GND_net), .I1(n16618[0]), .I2(n264_adj_3837), 
            .I3(n37614), .O(n16569[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_9_lut (.I0(GND_net), .I1(n8329[6]), .I2(GND_net), 
            .I3(n37418), .O(n8311[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_14 (.CI(n36484), .I0(n10669[11]), .I1(GND_net), 
            .CO(n36485));
    SB_CARRY add_3059_5 (.CI(n37234), .I0(n8131[2]), .I1(n407_adj_3836), 
            .CO(n37235));
    SB_LUT4 add_3140_13_lut (.I0(GND_net), .I1(n10669[10]), .I2(GND_net), 
            .I3(n36483), .O(n9927[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_13_lut (.I0(GND_net), .I1(n1799[10]), .I2(GND_net), 
            .I3(n37693), .O(n1798[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_13 (.CI(n37693), .I0(n1799[10]), .I1(GND_net), 
            .CO(n37694));
    SB_CARRY add_3479_3 (.CI(n37614), .I0(n16618[0]), .I1(n264_adj_3837), 
            .CO(n37615));
    SB_LUT4 sub_11_inv_0_i22_1_lut (.I0(\PID_CONTROLLER.err[21] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[21]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21902_6 (.CI(n36197), .I0(n57[4]), .I1(n191[4]), .CO(n36198));
    SB_LUT4 mult_14_add_1213_12_lut (.I0(GND_net), .I1(n1799[9]), .I2(GND_net), 
            .I3(n37692), .O(n1798[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[9]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n79[6]), 
            .I3(n35969), .O(pwm_23__N_2960[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_13 (.CI(n36483), .I0(n10669[10]), .I1(GND_net), 
            .CO(n36484));
    SB_LUT4 sub_11_inv_0_i23_1_lut (.I0(\PID_CONTROLLER.err[22] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[22]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_14_add_1213_12 (.CI(n37692), .I0(n1799[9]), .I1(GND_net), 
            .CO(n37693));
    SB_CARRY unary_minus_17_add_3_8 (.CI(n35969), .I0(GND_net), .I1(n79[6]), 
            .CO(n35970));
    SB_LUT4 mult_14_add_1213_11_lut (.I0(GND_net), .I1(n1799[8]), .I2(GND_net), 
            .I3(n37691), .O(n1798[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_15_lut (.I0(GND_net), .I1(n1804[12]), .I2(GND_net), 
            .I3(n37810), .O(n1803[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_15 (.CI(n37810), .I0(n1804[12]), .I1(GND_net), 
            .CO(n37811));
    SB_LUT4 add_21902_5_lut (.I0(GND_net), .I1(n57[3]), .I2(n191[3]), 
            .I3(n36196), .O(\PID_CONTROLLER.result_31__N_3003 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_14_lut (.I0(GND_net), .I1(n1804[11]), .I2(GND_net), 
            .I3(n37809), .O(n1803[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3479_2_lut (.I0(GND_net), .I1(n86_adj_3389), .I2(n167_adj_3839), 
            .I3(GND_net), .O(n16569[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3479_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3479_2 (.CI(GND_net), .I0(n86_adj_3389), .I1(n167_adj_3839), 
            .CO(n37614));
    SB_LUT4 add_3140_12_lut (.I0(GND_net), .I1(n10669[9]), .I2(GND_net), 
            .I3(n36482), .O(n9927[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_11 (.CI(n37691), .I0(n1799[8]), .I1(GND_net), 
            .CO(n37692));
    SB_CARRY mult_14_add_1218_14 (.CI(n37809), .I0(n1804[11]), .I1(GND_net), 
            .CO(n37810));
    SB_LUT4 mult_14_add_1218_13_lut (.I0(GND_net), .I1(n1804[10]), .I2(GND_net), 
            .I3(n37808), .O(n1803[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_13 (.CI(n37808), .I0(n1804[10]), .I1(GND_net), 
            .CO(n37809));
    SB_LUT4 mult_14_add_1218_12_lut (.I0(GND_net), .I1(n1804[9]), .I2(GND_net), 
            .I3(n37807), .O(n1803[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_12 (.CI(n37807), .I0(n1804[9]), .I1(GND_net), 
            .CO(n37808));
    SB_LUT4 unary_minus_17_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n79[5]), 
            .I3(n35968), .O(pwm_23__N_2960[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_11_lut (.I0(GND_net), .I1(n1804[8]), .I2(GND_net), 
            .I3(n37806), .O(n1803[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_11 (.CI(n37806), .I0(n1804[8]), .I1(GND_net), 
            .CO(n37807));
    SB_LUT4 mult_14_add_1218_10_lut (.I0(GND_net), .I1(n1804[7]), .I2(GND_net), 
            .I3(n37805), .O(n1803[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_7 (.CI(n35968), .I0(GND_net), .I1(n79[5]), 
            .CO(n35969));
    SB_LUT4 add_3387_17_lut (.I0(GND_net), .I1(n15638[14]), .I2(GND_net), 
            .I3(n37613), .O(n15397[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i327_2_lut (.I0(\Kd[5] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n486));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i327_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3140_12 (.CI(n36482), .I0(n10669[9]), .I1(GND_net), .CO(n36483));
    SB_LUT4 mult_12_i87_2_lut (.I0(\Kd[1] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n128));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i24_2_lut (.I0(\Kd[0] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3487));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i24_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1218_10 (.CI(n37805), .I0(n1804[7]), .I1(GND_net), 
            .CO(n37806));
    SB_LUT4 add_3387_16_lut (.I0(GND_net), .I1(n15638[13]), .I2(GND_net), 
            .I3(n37612), .O(n15397[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_16 (.CI(n37612), .I0(n15638[13]), .I1(GND_net), 
            .CO(n37613));
    SB_LUT4 add_3387_15_lut (.I0(GND_net), .I1(n15638[12]), .I2(GND_net), 
            .I3(n37611), .O(n15397[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_11_lut (.I0(GND_net), .I1(n10669[8]), .I2(GND_net), 
            .I3(n36481), .O(n9927[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_9 (.CI(n37418), .I0(n8329[6]), .I1(GND_net), .CO(n37419));
    SB_LUT4 mult_12_i392_2_lut (.I0(\Kd[6] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n583_adj_3486));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1218_9_lut (.I0(GND_net), .I1(n1804[6]), .I2(GND_net), 
            .I3(n37804), .O(n1803[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_9 (.CI(n37804), .I0(n1804[6]), .I1(GND_net), 
            .CO(n37805));
    SB_LUT4 mult_12_i152_2_lut (.I0(\Kd[2] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n225_adj_3485));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i457_2_lut (.I0(\Kd[7] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n680));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1218_8_lut (.I0(GND_net), .I1(n1804[5]), .I2(n533), 
            .I3(n37803), .O(n1803[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i337_2_lut (.I0(\Kd[5] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n501));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i337_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1218_8 (.CI(n37803), .I0(n1804[5]), .I1(n533), 
            .CO(n37804));
    SB_LUT4 unary_minus_21_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[10]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_add_1218_7_lut (.I0(GND_net), .I1(n1804[4]), .I2(n460_adj_3845), 
            .I3(n37802), .O(n1803[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_5 (.CI(n36196), .I0(n57[3]), .I1(n191[3]), .CO(n36197));
    SB_CARRY add_3387_15 (.CI(n37611), .I0(n15638[12]), .I1(GND_net), 
            .CO(n37612));
    SB_LUT4 add_21902_4_lut (.I0(GND_net), .I1(n57[2]), .I2(n191[2]), 
            .I3(n36195), .O(\PID_CONTROLLER.result_31__N_3003 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_11 (.CI(n36481), .I0(n10669[8]), .I1(GND_net), .CO(n36482));
    SB_CARRY mult_14_add_1218_7 (.CI(n37802), .I0(n1804[4]), .I1(n460_adj_3845), 
            .CO(n37803));
    SB_LUT4 mult_14_add_1213_10_lut (.I0(GND_net), .I1(n1799[7]), .I2(GND_net), 
            .I3(n37690), .O(n1798[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_4_lut (.I0(GND_net), .I1(n8131[1]), .I2(n310_adj_3846), 
            .I3(n37233), .O(n8104[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_25_lut (.I0(\PID_CONTROLLER.result [23]), 
            .I1(n49815), .I2(n60[31]), .I3(n36057), .O(n448)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3140_10_lut (.I0(GND_net), .I1(n10669[7]), .I2(GND_net), 
            .I3(n36480), .O(n9927[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3387_14_lut (.I0(GND_net), .I1(n15638[11]), .I2(GND_net), 
            .I3(n37610), .O(n15397[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_24_lut (.I0(\PID_CONTROLLER.result [22]), 
            .I1(n49815), .I2(n60[22]), .I3(n36056), .O(n449)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mult_12_i217_2_lut (.I0(\Kd[3] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n322));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n79[4]), 
            .I3(n35967), .O(pwm_23__N_2960[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_10 (.CI(n36480), .I0(n10669[7]), .I1(GND_net), .CO(n36481));
    SB_CARRY unary_minus_23_add_3_24 (.CI(n36056), .I0(n49815), .I1(n60[22]), 
            .CO(n36057));
    SB_LUT4 add_3140_9_lut (.I0(GND_net), .I1(n10669[6]), .I2(GND_net), 
            .I3(n36479), .O(n9927[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_6 (.CI(n35967), .I0(GND_net), .I1(n79[4]), 
            .CO(n35968));
    SB_CARRY mult_14_add_1213_10 (.CI(n37690), .I0(n1799[7]), .I1(GND_net), 
            .CO(n37691));
    SB_LUT4 unary_minus_23_add_3_23_lut (.I0(\PID_CONTROLLER.result[21] ), 
            .I1(n49815), .I2(n60[21]), .I3(n36055), .O(n28362)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3078_14_lut (.I0(GND_net), .I1(n8470[11]), .I2(GND_net), 
            .I3(n37528), .O(n8446[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21902_4 (.CI(n36195), .I0(n57[2]), .I1(n191[2]), .CO(n36196));
    SB_LUT4 mult_14_add_1213_9_lut (.I0(GND_net), .I1(n1799[6]), .I2(GND_net), 
            .I3(n37689), .O(n1798[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_9 (.CI(n36479), .I0(n10669[6]), .I1(GND_net), .CO(n36480));
    SB_LUT4 add_3140_8_lut (.I0(GND_net), .I1(n10669[5]), .I2(n692_adj_3850), 
            .I3(n36478), .O(n9927[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_9 (.CI(n37689), .I0(n1799[6]), .I1(GND_net), 
            .CO(n37690));
    SB_LUT4 mult_14_add_1218_6_lut (.I0(GND_net), .I1(n1804[3]), .I2(n387_c), 
            .I3(n37801), .O(n1803[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_8_lut (.I0(GND_net), .I1(n1799[5]), .I2(n518), 
            .I3(n37688), .O(n1798[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_8 (.CI(n37688), .I0(n1799[5]), .I1(n518), 
            .CO(n37689));
    SB_CARRY mult_14_add_1218_6 (.CI(n37801), .I0(n1804[3]), .I1(n387_c), 
            .CO(n37802));
    SB_CARRY add_3078_14 (.CI(n37528), .I0(n8470[11]), .I1(GND_net), .CO(n37529));
    SB_LUT4 mult_14_add_1218_5_lut (.I0(GND_net), .I1(n1804[2]), .I2(n314_adj_3852), 
            .I3(n37800), .O(n1803[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_5 (.CI(n37800), .I0(n1804[2]), .I1(n314_adj_3852), 
            .CO(n37801));
    SB_LUT4 mult_14_add_1218_4_lut (.I0(GND_net), .I1(n1804[1]), .I2(n241_adj_3854), 
            .I3(n37799), .O(n1803[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_4 (.CI(n37799), .I0(n1804[1]), .I1(n241_adj_3854), 
            .CO(n37800));
    SB_LUT4 mult_14_add_1218_3_lut (.I0(GND_net), .I1(n1804[0]), .I2(n168_adj_3856), 
            .I3(n37798), .O(n1803[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_14 (.CI(n37610), .I0(n15638[11]), .I1(GND_net), 
            .CO(n37611));
    SB_CARRY add_3140_8 (.CI(n36478), .I0(n10669[5]), .I1(n692_adj_3850), 
            .CO(n36479));
    SB_CARRY mult_14_add_1218_3 (.CI(n37798), .I0(n1804[0]), .I1(n168_adj_3856), 
            .CO(n37799));
    SB_LUT4 mult_14_add_1213_7_lut (.I0(GND_net), .I1(n1799[4]), .I2(n445), 
            .I3(n37687), .O(n1798[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_7 (.CI(n37687), .I0(n1799[4]), .I1(n445), 
            .CO(n37688));
    SB_LUT4 mult_14_add_1218_2_lut (.I0(GND_net), .I1(n26_adj_3857), .I2(n95), 
            .I3(GND_net), .O(n1803[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_2 (.CI(GND_net), .I0(n26_adj_3857), .I1(n95), 
            .CO(n37798));
    SB_LUT4 mult_14_i193_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i193_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i402_2_lut (.I0(\Kd[6] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n598));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_23_add_3_23 (.CI(n36055), .I0(n49815), .I1(n60[21]), 
            .CO(n36056));
    SB_LUT4 mult_12_i467_2_lut (.I0(\Kd[7] ), .I1(n69[5]), .I2(GND_net), 
            .I3(GND_net), .O(n695));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i242_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i242_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3387_13_lut (.I0(GND_net), .I1(n15638[10]), .I2(GND_net), 
            .I3(n37609), .O(n15397[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i97_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n143_adj_3380));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3379));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n79[3]), 
            .I3(n35966), .O(pwm_23__N_2960[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_inv_0_i24_1_lut (.I0(\PID_CONTROLLER.err[23] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[23]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3078_13_lut (.I0(GND_net), .I1(n8470[10]), .I2(GND_net), 
            .I3(n37527), .O(n8446[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_24_lut (.I0(GND_net), .I1(n1803[21]), .I2(GND_net), 
            .I3(n37796), .O(n1802[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_7_lut (.I0(GND_net), .I1(n10669[4]), .I2(n595_adj_3859), 
            .I3(n36477), .O(n9927[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21902_3_lut (.I0(GND_net), .I1(n57[1]), .I2(n191[1]), 
            .I3(n36194), .O(\PID_CONTROLLER.result_31__N_3003 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_7 (.CI(n36477), .I0(n10669[4]), .I1(n595_adj_3859), 
            .CO(n36478));
    SB_CARRY unary_minus_17_add_3_5 (.CI(n35966), .I0(GND_net), .I1(n79[3]), 
            .CO(n35967));
    SB_LUT4 add_3140_6_lut (.I0(GND_net), .I1(n10669[3]), .I2(n498_adj_3860), 
            .I3(n36476), .O(n9927[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_6 (.CI(n36476), .I0(n10669[3]), .I1(n498_adj_3860), 
            .CO(n36477));
    SB_CARRY add_21902_3 (.CI(n36194), .I0(n57[1]), .I1(n191[1]), .CO(n36195));
    SB_LUT4 add_3068_8_lut (.I0(GND_net), .I1(n8329[5]), .I2(n725), .I3(n37417), 
            .O(n8311[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_5_lut (.I0(GND_net), .I1(n10669[2]), .I2(n401_adj_3861), 
            .I3(n36475), .O(n9927[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3059_4 (.CI(n37233), .I0(n8131[1]), .I1(n310_adj_3846), 
            .CO(n37234));
    SB_CARRY add_3387_13 (.CI(n37609), .I0(n15638[10]), .I1(GND_net), 
            .CO(n37610));
    SB_CARRY add_3078_13 (.CI(n37527), .I0(n8470[10]), .I1(GND_net), .CO(n37528));
    SB_CARRY add_3140_5 (.CI(n36475), .I0(n10669[2]), .I1(n401_adj_3861), 
            .CO(n36476));
    SB_CARRY mult_14_add_1217_24 (.CI(n37796), .I0(n1803[21]), .I1(GND_net), 
            .CO(n1707));
    SB_LUT4 mult_14_add_1213_6_lut (.I0(GND_net), .I1(n1799[3]), .I2(n372), 
            .I3(n37686), .O(n1798[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3068_8 (.CI(n37417), .I0(n8329[5]), .I1(n725), .CO(n37418));
    SB_LUT4 mult_14_add_1217_23_lut (.I0(GND_net), .I1(n1803[20]), .I2(GND_net), 
            .I3(n37795), .O(n1802[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_23 (.CI(n37795), .I0(n1803[20]), .I1(GND_net), 
            .CO(n37796));
    SB_LUT4 mult_14_add_1217_22_lut (.I0(GND_net), .I1(n1803[19]), .I2(GND_net), 
            .I3(n37794), .O(n1802[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_6 (.CI(n37686), .I0(n1799[3]), .I1(n372), 
            .CO(n37687));
    SB_LUT4 add_3059_3_lut (.I0(GND_net), .I1(n8131[0]), .I2(n213_adj_3862), 
            .I3(n37232), .O(n8104[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_4_lut (.I0(GND_net), .I1(n10669[1]), .I2(n304_adj_3863), 
            .I3(n36474), .O(n9927[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3078_12_lut (.I0(GND_net), .I1(n8470[9]), .I2(GND_net), 
            .I3(n37526), .O(n8446[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_4 (.CI(n36474), .I0(n10669[1]), .I1(n304_adj_3863), 
            .CO(n36475));
    SB_LUT4 add_21902_2_lut (.I0(GND_net), .I1(n57[0]), .I2(n191[0]), 
            .I3(GND_net), .O(\PID_CONTROLLER.result_31__N_3003 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21902_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3140_3_lut (.I0(GND_net), .I1(n10669[0]), .I2(n207_adj_3864), 
            .I3(n36473), .O(n9927[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_3 (.CI(n36473), .I0(n10669[0]), .I1(n207_adj_3864), 
            .CO(n36474));
    SB_CARRY add_21902_2 (.CI(GND_net), .I0(n57[0]), .I1(n191[0]), .CO(n36194));
    SB_LUT4 add_3140_2_lut (.I0(GND_net), .I1(n17_adj_3865), .I2(n110_adj_3866), 
            .I3(GND_net), .O(n9927[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3140_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3140_2 (.CI(GND_net), .I0(n17_adj_3865), .I1(n110_adj_3866), 
            .CO(n36473));
    SB_LUT4 add_3352_19_lut (.I0(GND_net), .I1(n15112[16]), .I2(GND_net), 
            .I3(n36193), .O(n14791[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3320_13_lut (.I0(GND_net), .I1(n14558[10]), .I2(GND_net), 
            .I3(n36472), .O(n14166[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3320_12_lut (.I0(GND_net), .I1(n14558[9]), .I2(GND_net), 
            .I3(n36471), .O(n14166[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i2  (.Q(\PID_CONTROLLER.err_prev[1] ), 
           .C(clk32MHz), .D(n23732));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i3  (.Q(\PID_CONTROLLER.err_prev[2] ), 
           .C(clk32MHz), .D(n23731));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY mult_14_add_1217_22 (.CI(n37794), .I0(n1803[19]), .I1(GND_net), 
            .CO(n37795));
    SB_DFF \PID_CONTROLLER.err_prev__i4  (.Q(\PID_CONTROLLER.err_prev[3] ), 
           .C(clk32MHz), .D(n23730));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i5  (.Q(\PID_CONTROLLER.err_prev[4] ), 
           .C(clk32MHz), .D(n23729));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i6  (.Q(\PID_CONTROLLER.err_prev[5] ), 
           .C(clk32MHz), .D(n23728));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i7  (.Q(\PID_CONTROLLER.err_prev[6] ), 
           .C(clk32MHz), .D(n23727));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i8  (.Q(\PID_CONTROLLER.err_prev[7] ), 
           .C(clk32MHz), .D(n23726));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3352_18_lut (.I0(GND_net), .I1(n15112[15]), .I2(GND_net), 
            .I3(n36192), .O(n14791[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i9  (.Q(\PID_CONTROLLER.err_prev[8] ), 
           .C(clk32MHz), .D(n23725));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_3320_12 (.CI(n36471), .I0(n14558[9]), .I1(GND_net), .CO(n36472));
    SB_DFF \PID_CONTROLLER.err_prev__i10  (.Q(\PID_CONTROLLER.err_prev[9] ), 
           .C(clk32MHz), .D(n23724));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_3059_3 (.CI(n37232), .I0(n8131[0]), .I1(n213_adj_3862), 
            .CO(n37233));
    SB_DFF \PID_CONTROLLER.err_prev__i11  (.Q(\PID_CONTROLLER.err_prev[10] ), 
           .C(clk32MHz), .D(n23723));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i12  (.Q(\PID_CONTROLLER.err_prev[11] ), 
           .C(clk32MHz), .D(n23722));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i13  (.Q(\PID_CONTROLLER.err_prev[12] ), 
           .C(clk32MHz), .D(n23721));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i14  (.Q(\PID_CONTROLLER.err_prev[13] ), 
           .C(clk32MHz), .D(n23720));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i15  (.Q(\PID_CONTROLLER.err_prev[14] ), 
           .C(clk32MHz), .D(n23719));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i16  (.Q(\PID_CONTROLLER.err_prev[15] ), 
           .C(clk32MHz), .D(n23718));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i17  (.Q(\PID_CONTROLLER.err_prev[16] ), 
           .C(clk32MHz), .D(n23717));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3320_11_lut (.I0(GND_net), .I1(n14558[8]), .I2(GND_net), 
            .I3(n36470), .O(n14166[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i18  (.Q(\PID_CONTROLLER.err_prev[17] ), 
           .C(clk32MHz), .D(n23716));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_3352_18 (.CI(n36192), .I0(n15112[15]), .I1(GND_net), 
            .CO(n36193));
    SB_DFF \PID_CONTROLLER.err_prev__i19  (.Q(\PID_CONTROLLER.err_prev[18] ), 
           .C(clk32MHz), .D(n23715));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_3320_11 (.CI(n36470), .I0(n14558[8]), .I1(GND_net), .CO(n36471));
    SB_DFF \PID_CONTROLLER.err_prev__i20  (.Q(\PID_CONTROLLER.err_prev[19] ), 
           .C(clk32MHz), .D(n23714));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i21  (.Q(\PID_CONTROLLER.err_prev[20] ), 
           .C(clk32MHz), .D(n23713));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3320_10_lut (.I0(GND_net), .I1(n14558[7]), .I2(GND_net), 
            .I3(n36469), .O(n14166[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i22  (.Q(\PID_CONTROLLER.err_prev[21] ), 
           .C(clk32MHz), .D(n23712));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3352_17_lut (.I0(GND_net), .I1(n15112[14]), .I2(GND_net), 
            .I3(n36191), .O(n14791[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i23  (.Q(\PID_CONTROLLER.err_prev[22] ), 
           .C(clk32MHz), .D(n23711));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_3320_10 (.CI(n36469), .I0(n14558[7]), .I1(GND_net), .CO(n36470));
    SB_DFF \PID_CONTROLLER.err_prev__i24  (.Q(\PID_CONTROLLER.err_prev[23] ), 
           .C(clk32MHz), .D(n23710));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_prev__i25  (.Q(\PID_CONTROLLER.err_prev[31] ), 
           .C(clk32MHz), .D(n23709));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 mult_14_add_1217_21_lut (.I0(GND_net), .I1(n1803[18]), .I2(GND_net), 
            .I3(n37793), .O(n1802[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3320_9_lut (.I0(GND_net), .I1(n14558[6]), .I2(GND_net), 
            .I3(n36468), .O(n14166[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_17 (.CI(n36191), .I0(n15112[14]), .I1(GND_net), 
            .CO(n36192));
    SB_CARRY add_3320_9 (.CI(n36468), .I0(n14558[6]), .I1(GND_net), .CO(n36469));
    SB_CARRY mult_14_add_1217_21 (.CI(n37793), .I0(n1803[18]), .I1(GND_net), 
            .CO(n37794));
    SB_LUT4 add_3320_8_lut (.I0(GND_net), .I1(n14558[5]), .I2(n545), .I3(n36467), 
            .O(n14166[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_16_lut (.I0(GND_net), .I1(n15112[13]), .I2(GND_net), 
            .I3(n36190), .O(n14791[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3320_8 (.CI(n36467), .I0(n14558[5]), .I1(n545), .CO(n36468));
    SB_LUT4 add_3068_7_lut (.I0(GND_net), .I1(n8329[4]), .I2(n628), .I3(n37416), 
            .O(n8311[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3059_2_lut (.I0(GND_net), .I1(n23_adj_3867), .I2(n116_adj_3868), 
            .I3(GND_net), .O(n8104[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3059_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_16 (.CI(n36190), .I0(n15112[13]), .I1(GND_net), 
            .CO(n36191));
    SB_LUT4 mult_14_add_1217_20_lut (.I0(GND_net), .I1(n1803[17]), .I2(GND_net), 
            .I3(n37792), .O(n1802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3320_7_lut (.I0(GND_net), .I1(n14558[4]), .I2(n472), .I3(n36466), 
            .O(n14166[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_15_lut (.I0(GND_net), .I1(n15112[12]), .I2(GND_net), 
            .I3(n36189), .O(n14791[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3320_7 (.CI(n36466), .I0(n14558[4]), .I1(n472), .CO(n36467));
    SB_LUT4 unary_minus_23_add_3_22_lut (.I0(\PID_CONTROLLER.result[20] ), 
            .I1(n49815), .I2(n60[20]), .I3(n36054), .O(n1_adj_3869)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3068_7 (.CI(n37416), .I0(n8329[4]), .I1(n628), .CO(n37417));
    SB_LUT4 unary_minus_17_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n79[2]), 
            .I3(n35965), .O(pwm_23__N_2960[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3387_12_lut (.I0(GND_net), .I1(n15638[9]), .I2(GND_net), 
            .I3(n37608), .O(n15397[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_15 (.CI(n36189), .I0(n15112[12]), .I1(GND_net), 
            .CO(n36190));
    SB_CARRY unary_minus_17_add_3_4 (.CI(n35965), .I0(GND_net), .I1(n79[2]), 
            .CO(n35966));
    SB_LUT4 i22079_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n37873));   // verilog/motorControl.v(43[17:23])
    defparam i22079_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF \PID_CONTROLLER.result_i1  (.Q(\PID_CONTROLLER.result [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [1]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3320_6_lut (.I0(GND_net), .I1(n14558[3]), .I2(n399_c), 
            .I3(n36465), .O(n14166[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_5_lut (.I0(GND_net), .I1(n1799[2]), .I2(n299_adj_3871), 
            .I3(n37685), .O(n1798[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_14_lut (.I0(GND_net), .I1(n15112[11]), .I2(GND_net), 
            .I3(n36188), .O(n14791[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3320_6 (.CI(n36465), .I0(n14558[3]), .I1(n399_c), .CO(n36466));
    SB_LUT4 add_3320_5_lut (.I0(GND_net), .I1(n14558[2]), .I2(n326), .I3(n36464), 
            .O(n14166[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_6_lut (.I0(GND_net), .I1(n8329[3]), .I2(n531_adj_3872), 
            .I3(n37415), .O(n8311[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n79[1]), 
            .I3(n35964), .O(pwm_23__N_2960[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3320_5 (.CI(n36464), .I0(n14558[2]), .I1(n326), .CO(n36465));
    SB_CARRY unary_minus_23_add_3_22 (.CI(n36054), .I0(n49815), .I1(n60[20]), 
            .CO(n36055));
    SB_CARRY add_3068_6 (.CI(n37415), .I0(n8329[3]), .I1(n531_adj_3872), 
            .CO(n37416));
    SB_CARRY unary_minus_17_add_3_3 (.CI(n35964), .I0(GND_net), .I1(n79[1]), 
            .CO(n35965));
    SB_LUT4 unary_minus_17_add_3_2_lut (.I0(n28894), .I1(GND_net), .I2(n79[0]), 
            .I3(VCC_net), .O(n46591)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3352_14 (.CI(n36188), .I0(n15112[11]), .I1(GND_net), 
            .CO(n36189));
    SB_LUT4 add_3320_4_lut (.I0(GND_net), .I1(n14558[1]), .I2(n253), .I3(n36463), 
            .O(n14166[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3320_4 (.CI(n36463), .I0(n14558[1]), .I1(n253), .CO(n36464));
    SB_CARRY add_3059_2 (.CI(GND_net), .I0(n23_adj_3867), .I1(n116_adj_3868), 
            .CO(n37232));
    SB_LUT4 add_3320_3_lut (.I0(GND_net), .I1(n14558[0]), .I2(n180), .I3(n36462), 
            .O(n14166[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3320_3 (.CI(n36462), .I0(n14558[0]), .I1(n180), .CO(n36463));
    SB_LUT4 add_3352_13_lut (.I0(GND_net), .I1(n15112[10]), .I2(GND_net), 
            .I3(n36187), .O(n14791[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3320_2_lut (.I0(GND_net), .I1(n35), .I2(n107), .I3(GND_net), 
            .O(n14166[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3320_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_27_lut (.I0(GND_net), .I1(n8104[24]), .I2(GND_net), 
            .I3(n37231), .O(n8076[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_20 (.CI(n37792), .I0(n1803[17]), .I1(GND_net), 
            .CO(n37793));
    SB_CARRY add_3320_2 (.CI(GND_net), .I0(n35), .I1(n107), .CO(n36462));
    SB_CARRY add_3352_13 (.CI(n36187), .I0(n15112[10]), .I1(GND_net), 
            .CO(n36188));
    SB_LUT4 add_3352_12_lut (.I0(GND_net), .I1(n15112[9]), .I2(GND_net), 
            .I3(n36186), .O(n14791[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3168_27_lut (.I0(GND_net), .I1(n11356[24]), .I2(GND_net), 
            .I3(n36461), .O(n10669[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3168_26_lut (.I0(GND_net), .I1(n11356[23]), .I2(GND_net), 
            .I3(n36460), .O(n10669[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_12 (.CI(n37608), .I0(n15638[9]), .I1(GND_net), .CO(n37609));
    SB_CARRY add_3168_26 (.CI(n36460), .I0(n11356[23]), .I1(GND_net), 
            .CO(n36461));
    SB_CARRY add_3352_12 (.CI(n36186), .I0(n15112[9]), .I1(GND_net), .CO(n36187));
    SB_LUT4 unary_minus_23_add_3_21_lut (.I0(\PID_CONTROLLER.result [19]), 
            .I1(n49815), .I2(n60[19]), .I3(n36053), .O(n452)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY unary_minus_23_add_3_21 (.CI(n36053), .I0(n49815), .I1(n60[19]), 
            .CO(n36054));
    SB_LUT4 add_3168_25_lut (.I0(GND_net), .I1(n11356[22]), .I2(GND_net), 
            .I3(n36459), .O(n10669[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n79[0]), 
            .CO(n35964));
    SB_LUT4 add_3352_11_lut (.I0(GND_net), .I1(n15112[8]), .I2(GND_net), 
            .I3(n36185), .O(n14791[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_25 (.CI(n36459), .I0(n11356[22]), .I1(GND_net), 
            .CO(n36460));
    SB_LUT4 add_3168_24_lut (.I0(GND_net), .I1(n11356[21]), .I2(GND_net), 
            .I3(n36458), .O(n10669[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_11 (.CI(n36185), .I0(n15112[8]), .I1(GND_net), .CO(n36186));
    SB_CARRY add_3168_24 (.CI(n36458), .I0(n11356[21]), .I1(GND_net), 
            .CO(n36459));
    SB_LUT4 add_3168_23_lut (.I0(GND_net), .I1(n11356[20]), .I2(GND_net), 
            .I3(n36457), .O(n10669[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_10_lut (.I0(GND_net), .I1(n15112[7]), .I2(GND_net), 
            .I3(n36184), .O(n14791[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_23 (.CI(n36457), .I0(n11356[20]), .I1(GND_net), 
            .CO(n36458));
    SB_CARRY add_3078_12 (.CI(n37526), .I0(n8470[9]), .I1(GND_net), .CO(n37527));
    SB_LUT4 add_3068_5_lut (.I0(GND_net), .I1(n8329[2]), .I2(n434_adj_3876), 
            .I3(n37414), .O(n8311[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_26_lut (.I0(GND_net), .I1(n8104[23]), .I2(GND_net), 
            .I3(n37230), .O(n8076[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3168_22_lut (.I0(GND_net), .I1(n11356[19]), .I2(GND_net), 
            .I3(n36456), .O(n10669[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_10 (.CI(n36184), .I0(n15112[7]), .I1(GND_net), .CO(n36185));
    SB_CARRY add_3168_22 (.CI(n36456), .I0(n11356[19]), .I1(GND_net), 
            .CO(n36457));
    SB_LUT4 add_3168_21_lut (.I0(GND_net), .I1(n11356[18]), .I2(GND_net), 
            .I3(n36455), .O(n10669[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_9_lut (.I0(GND_net), .I1(n15112[6]), .I2(GND_net), 
            .I3(n36183), .O(n14791[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_21 (.CI(n36455), .I0(n11356[18]), .I1(GND_net), 
            .CO(n36456));
    SB_DFF \PID_CONTROLLER.result_i2  (.Q(\PID_CONTROLLER.result [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [2]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i3  (.Q(\PID_CONTROLLER.result [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [3]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i4  (.Q(\PID_CONTROLLER.result [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [4]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i5  (.Q(\PID_CONTROLLER.result[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [5]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i6  (.Q(\PID_CONTROLLER.result [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [6]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i7  (.Q(\PID_CONTROLLER.result[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [7]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i8  (.Q(\PID_CONTROLLER.result [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [8]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i9  (.Q(\PID_CONTROLLER.result [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [9]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i10  (.Q(\PID_CONTROLLER.result [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [10]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i11  (.Q(\PID_CONTROLLER.result [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [11]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i12  (.Q(\PID_CONTROLLER.result [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [12]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i13  (.Q(\PID_CONTROLLER.result[13] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [13]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i14  (.Q(\PID_CONTROLLER.result[14] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [14]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i15  (.Q(\PID_CONTROLLER.result [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [15]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i16  (.Q(\PID_CONTROLLER.result [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [16]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i17  (.Q(\PID_CONTROLLER.result [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [17]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i18  (.Q(\PID_CONTROLLER.result [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [18]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i19  (.Q(\PID_CONTROLLER.result [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [19]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i20  (.Q(\PID_CONTROLLER.result[20] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [20]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i21  (.Q(\PID_CONTROLLER.result[21] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [21]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i22  (.Q(\PID_CONTROLLER.result [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [22]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i23  (.Q(\PID_CONTROLLER.result [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [23]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i24  (.Q(\PID_CONTROLLER.result [24]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [24]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i25  (.Q(\PID_CONTROLLER.result [25]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [25]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i26  (.Q(\PID_CONTROLLER.result [26]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [26]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i27  (.Q(\PID_CONTROLLER.result [27]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [27]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i28  (.Q(\PID_CONTROLLER.result [28]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [28]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i29  (.Q(\PID_CONTROLLER.result [29]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [29]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i30  (.Q(\PID_CONTROLLER.result [30]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [30]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.result_i31  (.Q(\PID_CONTROLLER.result [31]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_3003 [31]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err[1] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [1]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF GATES_i3 (.Q(PIN_8_c_2), .C(clk32MHz), .D(GATES_5__N_2788[2]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i4 (.Q(PIN_9_c_3), .C(clk32MHz), .D(GATES_5__N_2788[3]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i5 (.Q(PIN_10_c_4), .C(clk32MHz), .D(GATES_5__N_2788[4]));   // verilog/motorControl.v(64[10] 111[6])
    SB_DFF GATES_i6 (.Q(PIN_11_c_5), .C(clk32MHz), .D(GATES_5__N_2788[5]));   // verilog/motorControl.v(64[10] 111[6])
    SB_CARRY mult_14_add_1213_5 (.CI(n37685), .I0(n1799[2]), .I1(n299_adj_3871), 
            .CO(n37686));
    SB_LUT4 mult_14_add_1213_4_lut (.I0(GND_net), .I1(n1799[1]), .I2(n226_adj_3877), 
            .I3(n37684), .O(n1798[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_4 (.CI(n37684), .I0(n1799[1]), .I1(n226_adj_3877), 
            .CO(n37685));
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err[2] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [2]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3168_20_lut (.I0(GND_net), .I1(n11356[17]), .I2(GND_net), 
            .I3(n36454), .O(n10669[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_9 (.CI(n36183), .I0(n15112[6]), .I1(GND_net), .CO(n36184));
    SB_CARRY add_3168_20 (.CI(n36454), .I0(n11356[17]), .I1(GND_net), 
            .CO(n36455));
    SB_LUT4 add_3168_19_lut (.I0(GND_net), .I1(n11356[16]), .I2(GND_net), 
            .I3(n36453), .O(n10669[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_8_lut (.I0(GND_net), .I1(n15112[5]), .I2(n719_adj_3878), 
            .I3(n36182), .O(n14791[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_19 (.CI(n36453), .I0(n11356[16]), .I1(GND_net), 
            .CO(n36454));
    SB_CARRY add_3058_26 (.CI(n37230), .I0(n8104[23]), .I1(GND_net), .CO(n37231));
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err[3] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [3]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err[4] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [4]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [5]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [6]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [7]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err[8] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [8]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err[9] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [9]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err[10] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [10]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err[11] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [11]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err[12] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [12]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err[13] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [13]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err[14] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [14]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err[15] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [15]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err[16] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [16]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err[17] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [17]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err[18] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [18]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err[19] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [19]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err[20] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [20]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err[21] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [21]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err[22] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [22]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i24  (.Q(\PID_CONTROLLER.err[23] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [23]));   // verilog/motorControl.v(38[14] 59[8])
    SB_DFF \PID_CONTROLLER.err_i25  (.Q(\PID_CONTROLLER.err[31] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2825 [24]));   // verilog/motorControl.v(38[14] 59[8])
    SB_LUT4 add_3168_18_lut (.I0(GND_net), .I1(n11356[15]), .I2(GND_net), 
            .I3(n36452), .O(n10669[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_8 (.CI(n36182), .I0(n15112[5]), .I1(n719_adj_3878), 
            .CO(n36183));
    SB_CARRY add_3168_18 (.CI(n36452), .I0(n11356[15]), .I1(GND_net), 
            .CO(n36453));
    SB_LUT4 mult_12_i282_2_lut (.I0(\Kd[4] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n419));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3168_17_lut (.I0(GND_net), .I1(n11356[14]), .I2(GND_net), 
            .I3(n36451), .O(n10669[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_25_lut (.I0(GND_net), .I1(n8104[22]), .I2(GND_net), 
            .I3(n37229), .O(n8076[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_17 (.CI(n36451), .I0(n11356[14]), .I1(GND_net), 
            .CO(n36452));
    SB_CARRY add_3068_5 (.CI(n37414), .I0(n8329[2]), .I1(n434_adj_3876), 
            .CO(n37415));
    SB_LUT4 add_3168_16_lut (.I0(GND_net), .I1(n11356[13]), .I2(GND_net), 
            .I3(n36450), .O(n10669[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3068_4_lut (.I0(GND_net), .I1(n8329[1]), .I2(n337_adj_3879), 
            .I3(n37413), .O(n8311[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_7_lut (.I0(GND_net), .I1(n15112[4]), .I2(n622_adj_3880), 
            .I3(n36181), .O(n14791[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_16 (.CI(n36450), .I0(n11356[13]), .I1(GND_net), 
            .CO(n36451));
    SB_LUT4 add_3168_15_lut (.I0(GND_net), .I1(n11356[12]), .I2(GND_net), 
            .I3(n36449), .O(n10669[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3352_7 (.CI(n36181), .I0(n15112[4]), .I1(n622_adj_3880), 
            .CO(n36182));
    SB_CARRY add_3168_15 (.CI(n36449), .I0(n11356[12]), .I1(GND_net), 
            .CO(n36450));
    SB_LUT4 add_3168_14_lut (.I0(GND_net), .I1(n11356[11]), .I2(GND_net), 
            .I3(n36448), .O(n10669[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_6_lut (.I0(GND_net), .I1(n15112[3]), .I2(n525_adj_3881), 
            .I3(n36180), .O(n14791[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_14 (.CI(n36448), .I0(n11356[11]), .I1(GND_net), 
            .CO(n36449));
    SB_CARRY add_3068_4 (.CI(n37413), .I0(n8329[1]), .I1(n337_adj_3879), 
            .CO(n37414));
    SB_LUT4 mult_14_add_1213_3_lut (.I0(GND_net), .I1(n1799[0]), .I2(n153_adj_3882), 
            .I3(n37683), .O(n1798[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_20_lut (.I0(\PID_CONTROLLER.result [18]), 
            .I1(n49815), .I2(n60[18]), .I3(n36052), .O(n453)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mult_14_add_1213_3 (.CI(n37683), .I0(n1799[0]), .I1(n153_adj_3882), 
            .CO(n37684));
    SB_LUT4 mult_14_add_1213_2_lut (.I0(GND_net), .I1(n11_adj_3883), .I2(n80), 
            .I3(GND_net), .O(n1798[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_2 (.CI(GND_net), .I0(n11_adj_3883), .I1(n80), 
            .CO(n37683));
    SB_LUT4 mult_14_add_1212_24_lut (.I0(GND_net), .I1(n1798[21]), .I2(GND_net), 
            .I3(n37681), .O(n1797[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_24 (.CI(n37681), .I0(n1798[21]), .I1(GND_net), 
            .CO(n1687));
    SB_LUT4 mult_14_add_1212_23_lut (.I0(GND_net), .I1(n1798[20]), .I2(GND_net), 
            .I3(n37680), .O(n1797[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_25 (.CI(n37229), .I0(n8104[22]), .I1(GND_net), .CO(n37230));
    SB_CARRY unary_minus_23_add_3_20 (.CI(n36052), .I0(n49815), .I1(n60[18]), 
            .CO(n36053));
    SB_LUT4 add_3168_13_lut (.I0(GND_net), .I1(n11356[10]), .I2(GND_net), 
            .I3(n36447), .O(n10669[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_13 (.CI(n36447), .I0(n11356[10]), .I1(GND_net), 
            .CO(n36448));
    SB_CARRY add_3352_6 (.CI(n36180), .I0(n15112[3]), .I1(n525_adj_3881), 
            .CO(n36181));
    SB_LUT4 add_3168_12_lut (.I0(GND_net), .I1(n11356[9]), .I2(GND_net), 
            .I3(n36446), .O(n10669[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1013__i1 (.Q(Kd_delay_counter[1]), .C(clk32MHz), 
           .D(n70[1]));   // verilog/motorControl.v(55[27:47])
    SB_CARRY add_3168_12 (.CI(n36446), .I0(n11356[9]), .I1(GND_net), .CO(n36447));
    SB_LUT4 add_3352_5_lut (.I0(GND_net), .I1(n15112[2]), .I2(n428_adj_3884), 
            .I3(n36179), .O(n14791[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21911_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(GND_net), .O(n16635[0]));   // verilog/motorControl.v(43[17:23])
    defparam i21911_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 mult_12_i107_2_lut (.I0(\Kd[1] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n158));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i44_2_lut (.I0(\Kd[0] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n65));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i32_1_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[26]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i347_2_lut (.I0(\Kd[5] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n516_adj_3471));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i347_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3352_5 (.CI(n36179), .I0(n15112[2]), .I1(n428_adj_3884), 
            .CO(n36180));
    SB_LUT4 add_3168_11_lut (.I0(GND_net), .I1(n11356[8]), .I2(GND_net), 
            .I3(n36445), .O(n10669[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_11 (.CI(n36445), .I0(n11356[8]), .I1(GND_net), .CO(n36446));
    SB_LUT4 add_3352_4_lut (.I0(GND_net), .I1(n15112[1]), .I2(n331_adj_3885), 
            .I3(n36178), .O(n14791[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_24_lut (.I0(GND_net), .I1(n8104[21]), .I2(GND_net), 
            .I3(n37228), .O(n8076[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_19_lut (.I0(\PID_CONTROLLER.result [17]), 
            .I1(n49815), .I2(n60[17]), .I3(n36051), .O(n454)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3168_10_lut (.I0(GND_net), .I1(n11356[7]), .I2(GND_net), 
            .I3(n36444), .O(n10669[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_19 (.CI(n36051), .I0(n49815), .I1(n60[17]), 
            .CO(n36052));
    SB_LUT4 mult_14_add_1217_19_lut (.I0(GND_net), .I1(n1803[16]), .I2(GND_net), 
            .I3(n37791), .O(n1802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1013__i2 (.Q(Kd_delay_counter[2]), .C(clk32MHz), 
           .D(n70[2]));   // verilog/motorControl.v(55[27:47])
    SB_CARRY mult_14_add_1217_19 (.CI(n37791), .I0(n1803[16]), .I1(GND_net), 
            .CO(n37792));
    SB_CARRY add_3168_10 (.CI(n36444), .I0(n11356[7]), .I1(GND_net), .CO(n36445));
    SB_LUT4 add_3168_9_lut (.I0(GND_net), .I1(n11356[6]), .I2(GND_net), 
            .I3(n36443), .O(n10669[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_23 (.CI(n37680), .I0(n1798[20]), .I1(GND_net), 
            .CO(n37681));
    SB_CARRY add_3168_9 (.CI(n36443), .I0(n11356[6]), .I1(GND_net), .CO(n36444));
    SB_CARRY add_3352_4 (.CI(n36178), .I0(n15112[1]), .I1(n331_adj_3885), 
            .CO(n36179));
    SB_LUT4 add_3168_8_lut (.I0(GND_net), .I1(n11356[5]), .I2(n695_adj_3887), 
            .I3(n36442), .O(n10669[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3058_24 (.CI(n37228), .I0(n8104[21]), .I1(GND_net), .CO(n37229));
    SB_LUT4 mult_14_add_1212_22_lut (.I0(GND_net), .I1(n1798[19]), .I2(GND_net), 
            .I3(n37679), .O(n1797[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_8 (.CI(n36442), .I0(n11356[5]), .I1(n695_adj_3887), 
            .CO(n36443));
    SB_LUT4 add_3387_11_lut (.I0(GND_net), .I1(n15638[8]), .I2(GND_net), 
            .I3(n37607), .O(n15397[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_18_lut (.I0(\PID_CONTROLLER.result [16]), 
            .I1(n49815), .I2(n60[16]), .I3(n36050), .O(n455)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3168_7_lut (.I0(GND_net), .I1(n11356[4]), .I2(n598_adj_3889), 
            .I3(n36441), .O(n10669[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_23_lut (.I0(GND_net), .I1(n8104[20]), .I2(GND_net), 
            .I3(n37227), .O(n8076[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1013__i3 (.Q(Kd_delay_counter[3]), .C(clk32MHz), 
           .D(n70[3]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1013__i4 (.Q(Kd_delay_counter[4]), .C(clk32MHz), 
           .D(n70[4]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1013__i5 (.Q(Kd_delay_counter[5]), .C(clk32MHz), 
           .D(n70[5]));   // verilog/motorControl.v(55[27:47])
    SB_DFF Kd_delay_counter_1013__i6 (.Q(Kd_delay_counter[6]), .C(clk32MHz), 
           .D(n70[6]));   // verilog/motorControl.v(55[27:47])
    SB_DFF pwm_count_1014__i1 (.Q(pwm_count[1]), .C(clk32MHz), .D(n64[1]));   // verilog/motorControl.v(110[18:29])
    SB_CARRY add_3168_7 (.CI(n36441), .I0(n11356[4]), .I1(n598_adj_3889), 
            .CO(n36442));
    SB_LUT4 add_3352_3_lut (.I0(GND_net), .I1(n15112[0]), .I2(n234_adj_3890), 
            .I3(n36177), .O(n14791[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3168_6_lut (.I0(GND_net), .I1(n11356[3]), .I2(n501_adj_3891), 
            .I3(n36440), .O(n10669[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_6 (.CI(n36440), .I0(n11356[3]), .I1(n501_adj_3891), 
            .CO(n36441));
    SB_CARRY add_3352_3 (.CI(n36177), .I0(n15112[0]), .I1(n234_adj_3890), 
            .CO(n36178));
    SB_LUT4 add_3168_5_lut (.I0(GND_net), .I1(n11356[2]), .I2(n404_adj_3892), 
            .I3(n36439), .O(n10669[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3352_2_lut (.I0(GND_net), .I1(n44_adj_3893), .I2(n137_adj_3894), 
            .I3(GND_net), .O(n14791[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3352_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_18_lut (.I0(GND_net), .I1(n1803[15]), .I2(GND_net), 
            .I3(n37790), .O(n1802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3168_5 (.CI(n36439), .I0(n11356[2]), .I1(n404_adj_3892), 
            .CO(n36440));
    SB_LUT4 add_3168_4_lut (.I0(GND_net), .I1(n11356[1]), .I2(n307_adj_3895), 
            .I3(n36438), .O(n10669[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_18 (.CI(n36050), .I0(n49815), .I1(n60[16]), 
            .CO(n36051));
    SB_CARRY add_3168_4 (.CI(n36438), .I0(n11356[1]), .I1(n307_adj_3895), 
            .CO(n36439));
    SB_CARRY add_3352_2 (.CI(GND_net), .I0(n44_adj_3893), .I1(n137_adj_3894), 
            .CO(n36177));
    SB_LUT4 add_3168_3_lut (.I0(GND_net), .I1(n11356[0]), .I2(n210_adj_3896), 
            .I3(n36437), .O(n10669[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_17_lut (.I0(\PID_CONTROLLER.result [15]), 
            .I1(n49815), .I2(n60[15]), .I3(n36049), .O(n456)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3168_3 (.CI(n36437), .I0(n11356[0]), .I1(n210_adj_3896), 
            .CO(n36438));
    SB_LUT4 add_3168_2_lut (.I0(GND_net), .I1(n20_adj_3897), .I2(n113_adj_3898), 
            .I3(GND_net), .O(n10669[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_18 (.CI(n37790), .I0(n1803[15]), .I1(GND_net), 
            .CO(n37791));
    SB_LUT4 mult_14_add_1217_17_lut (.I0(GND_net), .I1(n1803[14]), .I2(GND_net), 
            .I3(n37789), .O(n1802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_22 (.CI(n37679), .I0(n1798[19]), .I1(GND_net), 
            .CO(n37680));
    SB_CARRY add_3387_11 (.CI(n37607), .I0(n15638[8]), .I1(GND_net), .CO(n37608));
    SB_LUT4 add_3078_11_lut (.I0(GND_net), .I1(n8470[8]), .I2(GND_net), 
            .I3(n37525), .O(n8446[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3078_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1014__i2 (.Q(pwm_count[2]), .C(clk32MHz), .D(n64[2]));   // verilog/motorControl.v(110[18:29])
    SB_CARRY mult_14_add_1217_17 (.CI(n37789), .I0(n1803[14]), .I1(GND_net), 
            .CO(n37790));
    SB_CARRY add_3168_2 (.CI(GND_net), .I0(n20_adj_3897), .I1(n113_adj_3898), 
            .CO(n36437));
    SB_LUT4 add_3068_3_lut (.I0(GND_net), .I1(n8329[0]), .I2(n240_adj_3899), 
            .I3(n37412), .O(n8311[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3068_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_23_add_3_17 (.CI(n36049), .I0(n49815), .I1(n60[15]), 
            .CO(n36050));
    SB_CARRY add_3058_23 (.CI(n37227), .I0(n8104[20]), .I1(GND_net), .CO(n37228));
    SB_LUT4 mult_14_add_1217_16_lut (.I0(GND_net), .I1(n1803[13]), .I2(GND_net), 
            .I3(n37788), .O(n1802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3340_12_lut (.I0(GND_net), .I1(n14910[9]), .I2(GND_net), 
            .I3(n36436), .O(n14558[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_16 (.CI(n37788), .I0(n1803[13]), .I1(GND_net), 
            .CO(n37789));
    SB_LUT4 add_3340_11_lut (.I0(GND_net), .I1(n14910[8]), .I2(GND_net), 
            .I3(n36435), .O(n14558[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3340_11 (.CI(n36435), .I0(n14910[8]), .I1(GND_net), .CO(n36436));
    SB_LUT4 mult_14_add_1217_15_lut (.I0(GND_net), .I1(n1803[12]), .I2(GND_net), 
            .I3(n37787), .O(n1802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3340_10_lut (.I0(GND_net), .I1(n14910[7]), .I2(GND_net), 
            .I3(n36434), .O(n14558[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3340_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_23_add_3_16_lut (.I0(\PID_CONTROLLER.result[14] ), 
            .I1(n49815), .I2(n60[14]), .I3(n36048), .O(n27734)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_23_add_3_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY mult_14_add_1217_15 (.CI(n37787), .I0(n1803[12]), .I1(GND_net), 
            .CO(n37788));
    SB_DFF pwm_count_1014__i3 (.Q(pwm_count[3]), .C(clk32MHz), .D(n64[3]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1014__i4 (.Q(pwm_count[4]), .C(clk32MHz), .D(n64[4]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1014__i5 (.Q(pwm_count[5]), .C(clk32MHz), .D(n64[5]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1014__i6 (.Q(pwm_count[6]), .C(clk32MHz), .D(n64[6]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1014__i7 (.Q(pwm_count[7]), .C(clk32MHz), .D(n64[7]));   // verilog/motorControl.v(110[18:29])
    SB_DFF pwm_count_1014__i8 (.Q(pwm_count[8]), .C(clk32MHz), .D(n64[8]));   // verilog/motorControl.v(110[18:29])
    SB_DFFE \PID_CONTROLLER.integral_1015__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[1]));   // verilog/motorControl.v(41[21:33])
    SB_LUT4 mult_14_add_1217_14_lut (.I0(GND_net), .I1(n1803[11]), .I2(GND_net), 
            .I3(n37786), .O(n1802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \PID_CONTROLLER.integral_1015__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[2]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1015__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[3]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1015__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[4]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1015__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[5]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1015__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[6]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1015__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[7]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1015__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[8]));   // verilog/motorControl.v(41[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1015__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(n55_adj_3726), .D(n61[9]));   // verilog/motorControl.v(41[21:33])
    SB_DFF \PID_CONTROLLER.err_prev__i1  (.Q(\PID_CONTROLLER.err_prev[0] ), 
           .C(clk32MHz), .D(n23574));   // verilog/motorControl.v(38[14] 59[8])
    SB_CARRY add_3068_3 (.CI(n37412), .I0(n8329[0]), .I1(n240_adj_3899), 
            .CO(n37413));
    SB_LUT4 add_3387_10_lut (.I0(GND_net), .I1(n15638[7]), .I2(GND_net), 
            .I3(n37606), .O(n15397[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3058_22_lut (.I0(GND_net), .I1(n8104[19]), .I2(GND_net), 
            .I3(n37226), .O(n8076[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3058_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_21_lut (.I0(GND_net), .I1(n1798[18]), .I2(GND_net), 
            .I3(n37678), .O(n1797[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_14 (.CI(n37786), .I0(n1803[11]), .I1(GND_net), 
            .CO(n37787));
    SB_CARRY add_3387_10 (.CI(n37606), .I0(n15638[7]), .I1(GND_net), .CO(n37607));
    SB_LUT4 mult_14_add_1217_13_lut (.I0(GND_net), .I1(n1803[10]), .I2(GND_net), 
            .I3(n37785), .O(n1802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_13 (.CI(n37785), .I0(n1803[10]), .I1(GND_net), 
            .CO(n37786));
    SB_LUT4 mult_14_add_1217_12_lut (.I0(GND_net), .I1(n1803[9]), .I2(GND_net), 
            .I3(n37784), .O(n1802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_12 (.CI(n37784), .I0(n1803[9]), .I1(GND_net), 
            .CO(n37785));
    SB_LUT4 mult_14_add_1217_11_lut (.I0(GND_net), .I1(n1803[8]), .I2(GND_net), 
            .I3(n37783), .O(n1802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_11 (.CI(n37783), .I0(n1803[8]), .I1(GND_net), 
            .CO(n37784));
    SB_CARRY mult_14_add_1212_21 (.CI(n37678), .I0(n1798[18]), .I1(GND_net), 
            .CO(n37679));
    SB_LUT4 add_3387_9_lut (.I0(GND_net), .I1(n15638[6]), .I2(GND_net), 
            .I3(n37605), .O(n15397[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_10_lut (.I0(GND_net), .I1(n1803[7]), .I2(GND_net), 
            .I3(n37782), .O(n1802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_10 (.CI(n37782), .I0(n1803[7]), .I1(GND_net), 
            .CO(n37783));
    SB_LUT4 mult_14_add_1217_9_lut (.I0(GND_net), .I1(n1803[6]), .I2(GND_net), 
            .I3(n37781), .O(n1802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_9 (.CI(n37605), .I0(n15638[6]), .I1(GND_net), .CO(n37606));
    SB_CARRY mult_14_add_1217_9 (.CI(n37781), .I0(n1803[6]), .I1(GND_net), 
            .CO(n37782));
    SB_LUT4 mult_14_add_1212_20_lut (.I0(GND_net), .I1(n1798[17]), .I2(GND_net), 
            .I3(n37677), .O(n1797[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3387_8_lut (.I0(GND_net), .I1(n15638[5]), .I2(n725_adj_3900), 
            .I3(n37604), .O(n15397[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_20 (.CI(n37677), .I0(n1798[17]), .I1(GND_net), 
            .CO(n37678));
    SB_CARRY add_3387_8 (.CI(n37604), .I0(n15638[5]), .I1(n725_adj_3900), 
            .CO(n37605));
    SB_LUT4 mult_14_add_1212_19_lut (.I0(GND_net), .I1(n1798[16]), .I2(GND_net), 
            .I3(n37676), .O(n1797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i412_2_lut (.I0(\Kd[6] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n613));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1217_8_lut (.I0(GND_net), .I1(n1803[5]), .I2(n530), 
            .I3(n37780), .O(n1802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_8 (.CI(n37780), .I0(n1803[5]), .I1(n530), 
            .CO(n37781));
    SB_LUT4 mult_14_add_1217_7_lut (.I0(GND_net), .I1(n1803[4]), .I2(n457), 
            .I3(n37779), .O(n1802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_7 (.CI(n37779), .I0(n1803[4]), .I1(n457), 
            .CO(n37780));
    SB_LUT4 mult_14_add_1217_6_lut (.I0(GND_net), .I1(n1803[3]), .I2(n384), 
            .I3(n37778), .O(n1802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_6 (.CI(n37778), .I0(n1803[3]), .I1(n384), 
            .CO(n37779));
    SB_LUT4 mult_14_add_1217_5_lut (.I0(GND_net), .I1(n1803[2]), .I2(n311_adj_3901), 
            .I3(n37777), .O(n1802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_5 (.CI(n37777), .I0(n1803[2]), .I1(n311_adj_3901), 
            .CO(n37778));
    SB_CARRY mult_14_add_1212_19 (.CI(n37676), .I0(n1798[16]), .I1(GND_net), 
            .CO(n37677));
    SB_LUT4 add_3387_7_lut (.I0(GND_net), .I1(n15638[4]), .I2(n628_adj_3902), 
            .I3(n37603), .O(n15397[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_18_lut (.I0(GND_net), .I1(n1798[15]), .I2(GND_net), 
            .I3(n37675), .O(n1797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_7 (.CI(n37603), .I0(n15638[4]), .I1(n628_adj_3902), 
            .CO(n37604));
    SB_CARRY add_3078_11 (.CI(n37525), .I0(n8470[8]), .I1(GND_net), .CO(n37526));
    SB_LUT4 mult_14_add_1217_4_lut (.I0(GND_net), .I1(n1803[1]), .I2(n238_adj_3903), 
            .I3(n37776), .O(n1802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_4 (.CI(n37776), .I0(n1803[1]), .I1(n238_adj_3903), 
            .CO(n37777));
    SB_LUT4 mult_14_add_1217_3_lut (.I0(GND_net), .I1(n1803[0]), .I2(n165_adj_3904), 
            .I3(n37775), .O(n1802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_3 (.CI(n37775), .I0(n1803[0]), .I1(n165_adj_3904), 
            .CO(n37776));
    SB_LUT4 mult_14_add_1217_2_lut (.I0(GND_net), .I1(n23_adj_3905), .I2(n92), 
            .I3(GND_net), .O(n1802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_2 (.CI(GND_net), .I0(n23_adj_3905), .I1(n92), 
            .CO(n37775));
    SB_LUT4 mult_14_add_1216_24_lut (.I0(GND_net), .I1(n1802[21]), .I2(GND_net), 
            .I3(n37773), .O(n1801[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_24 (.CI(n37773), .I0(n1802[21]), .I1(GND_net), 
            .CO(n1703));
    SB_LUT4 mult_14_add_1216_23_lut (.I0(GND_net), .I1(n1802[20]), .I2(GND_net), 
            .I3(n37772), .O(n1801[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_18 (.CI(n37675), .I0(n1798[15]), .I1(GND_net), 
            .CO(n37676));
    SB_LUT4 add_3387_6_lut (.I0(GND_net), .I1(n15638[3]), .I2(n531_adj_3906), 
            .I3(n37602), .O(n15397[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3387_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_17_lut (.I0(GND_net), .I1(n1798[14]), .I2(GND_net), 
            .I3(n37674), .O(n1797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3387_6 (.CI(n37602), .I0(n15638[3]), .I1(n531_adj_3906), 
            .CO(n37603));
    SB_LUT4 mult_14_i49_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n72));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i49_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[0]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i98_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n145));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i98_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_12_i477_2_lut (.I0(\Kd[7] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n710));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i172_2_lut (.I0(\Kd[2] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n255));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i147_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n218_adj_3463));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i147_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[1]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i237_2_lut (.I0(\Kd[3] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n352));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i302_2_lut (.I0(\Kd[4] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n449_c));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i367_2_lut (.I0(\Kd[5] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n546));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i432_2_lut (.I0(\Kd[6] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n643));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i497_2_lut (.I0(\Kd[7] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i71_2_lut (.I0(\Kd[1] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i8_2_lut (.I0(\Kd[0] ), .I1(n69[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3457));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i136_2_lut (.I0(\Kd[2] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n201));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i201_2_lut (.I0(\Kd[3] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n298));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i196_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n291));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i196_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i245_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n364_adj_3455));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i245_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[2]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i294_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n437_adj_3453));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i294_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_12_i266_2_lut (.I0(\Kd[4] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n395));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i343_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n510));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i343_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i392_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n583));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i392_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[3]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3451));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i331_2_lut (.I0(\Kd[5] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n492));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i89_2_lut (.I0(\Kd[1] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_3450));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i26_2_lut (.I0(\Kd[0] ), .I1(n69[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i146_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n216));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[15]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[4]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i211_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n313));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[5]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i396_2_lut (.I0(\Kd[6] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n589_adj_3446));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i276_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n410));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i154_2_lut (.I0(\Kd[2] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n228));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i341_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n507));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[6]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n604_adj_3444));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i461_2_lut (.I0(\Kd[7] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n686));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n701));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i219_2_lut (.I0(\Kd[3] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n325));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3443));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[7]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[16]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3439));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[8]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[17]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i284_2_lut (.I0(\Kd[4] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n422));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[9]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[10]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i349_2_lut (.I0(\Kd[5] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n519_adj_3434));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i109_2_lut (.I0(\Kd[1] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n161));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i46_2_lut (.I0(\Kd[0] ), .I1(n69[22]), .I2(GND_net), 
            .I3(GND_net), .O(n68));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i69_2_lut (.I0(\Kd[1] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i6_2_lut (.I0(\Kd[0] ), .I1(n69[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3433));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[18]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[11]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(n878), .I3(n17_adj_3907), 
            .O(GATES_5__N_2788[0]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i23_4_lut_4_lut.LUT_INIT = 16'h2044;
    SB_LUT4 mult_12_i134_2_lut (.I0(\Kd[2] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i199_2_lut (.I0(\Kd[3] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n295));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i505_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_3431));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[12]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[13]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i414_2_lut (.I0(\Kd[6] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n616));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i479_2_lut (.I0(\Kd[7] ), .I1(n69[11]), .I2(GND_net), 
            .I3(GND_net), .O(n713));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[14]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[19]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i78_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(GATES_5__N_3048[5]));   // verilog/motorControl.v(91[19:34])
    defparam i78_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(n42366));   // verilog/motorControl.v(86[14] 109[8])
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mult_14_i291_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n399_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i291_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1370 (.I0(n48211), .I1(pwm[21]), .I2(pwm[8]), 
            .I3(pwm_count[8]), .O(n20_adj_3908));
    defparam i5_4_lut_adj_1370.LUT_INIT = 16'hecfe;
    SB_LUT4 i11_4_lut (.I0(pwm[11]), .I1(pwm[17]), .I2(pwm[19]), .I3(pwm[15]), 
            .O(n26_adj_3909));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(pwm[16]), .I1(pwm[10]), .I2(pwm[14]), .I3(pwm[9]), 
            .O(n24_adj_3910));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(pwm[13]), .I1(n26_adj_3909), .I2(n20_adj_3908), 
            .I3(pwm[22]), .O(n28_adj_3911));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_3_lut (.I0(pwm[12]), .I1(pwm[18]), .I2(pwm[20]), .I3(GND_net), 
            .O(n23_adj_3912));
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(pwm[23]), .I1(n23_adj_3912), .I2(n28_adj_3911), 
            .I3(n24_adj_3910), .O(n17_adj_3907));   // verilog/motorControl.v(65[9:32])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_14_i340_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i340_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i162_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n240));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[11]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[12]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[13]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i389_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i389_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i73_4_lut (.I0(pwm[23]), .I1(n25), .I2(n30), .I3(n26), .O(n878));   // verilog/motorControl.v(86[19:44])
    defparam i73_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_2_lut_adj_1371 (.I0(hall3), .I1(n878), .I2(GND_net), .I3(GND_net), 
            .O(n42312));   // verilog/motorControl.v(86[14] 109[8])
    defparam i1_2_lut_adj_1371.LUT_INIT = 16'h4444;
    SB_LUT4 LessThan_22_i39_2_lut (.I0(\PID_CONTROLLER.result [19]), .I1(n67[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_3916));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i45_2_lut (.I0(\PID_CONTROLLER.result [22]), .I1(n67[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_3917));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i27570_2_lut (.I0(hall2), .I1(hall3), .I2(GND_net), .I3(GND_net), 
            .O(n43127));
    defparam i27570_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31869_3_lut (.I0(n42312), .I1(hall1), .I2(hall2), .I3(GND_net), 
            .O(n46681));   // verilog/motorControl.v(86[14] 109[8])
    defparam i31869_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 LessThan_22_i37_2_lut (.I0(\PID_CONTROLLER.result [18]), .I1(n67[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_3918));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34_4_lut (.I0(n46681), .I1(n43127), .I2(n17_adj_3907), .I3(n42366), 
            .O(n18_adj_3919));   // verilog/motorControl.v(86[14] 109[8])
    defparam i34_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i33_4_lut (.I0(n18_adj_3919), .I1(n17_adj_3907), .I2(GATES_5__N_3048[5]), 
            .I3(n42312), .O(GATES_5__N_2788[1]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i33_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 LessThan_22_i31_2_lut (.I0(\PID_CONTROLLER.result [15]), .I1(n67[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_3920));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i21_2_lut (.I0(\PID_CONTROLLER.result [10]), .I1(n67[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_3921));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i174_2_lut (.I0(\Kd[2] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i23_2_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n67[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3922));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i25_2_lut (.I0(\PID_CONTROLLER.result [12]), .I1(n67[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_3923));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n67[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3924));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n67[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3925));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n66[15]));   // verilog/motorControl.v(39[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_22_i9_2_lut (.I0(\PID_CONTROLLER.result [4]), .I1(n67[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3926));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i35_2_lut (.I0(\PID_CONTROLLER.result [17]), .I1(n67[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3927));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i33_2_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n67[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_3928));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i264_2_lut (.I0(\Kd[4] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n392));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i13_2_lut (.I0(\PID_CONTROLLER.result [6]), .I1(n67[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3929));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i329_2_lut (.I0(\Kd[5] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n489));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i329_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i394_2_lut (.I0(\Kd[6] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n586));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i239_2_lut (.I0(\Kd[3] ), .I1(n69[21]), .I2(GND_net), 
            .I3(GND_net), .O(n355));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i459_2_lut (.I0(\Kd[7] ), .I1(n69[1]), .I2(GND_net), 
            .I3(GND_net), .O(n683));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i99_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n146));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[14]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3424));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31258_4_lut (.I0(n27_adj_13), .I1(n15), .I2(n13_adj_3929), 
            .I3(n11), .O(n46817));
    defparam i31258_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_22_i12_3_lut (.I0(n413), .I1(n67[16]), .I2(n33_adj_3928), 
            .I3(GND_net), .O(n12_adj_3933));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_22_i10_3_lut (.I0(n415), .I1(n67[6]), .I2(n13_adj_3929), 
            .I3(GND_net), .O(n10_adj_3934));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_22_i30_3_lut (.I0(n12_adj_3933), .I1(n67[17]), .I2(n35_adj_3927), 
            .I3(GND_net), .O(n30_adj_3935));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32030_4_lut (.I0(n13_adj_3929), .I1(n11), .I2(n9_adj_3926), 
            .I3(n46851), .O(n47591));
    defparam i32030_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32024_4_lut (.I0(n19_adj_3925), .I1(n17_adj_3924), .I2(n15), 
            .I3(n47591), .O(n47585));
    defparam i32024_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33162_4_lut (.I0(n25_adj_3923), .I1(n23_adj_3922), .I2(n21_adj_3921), 
            .I3(n47585), .O(n48723));
    defparam i33162_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32614_4_lut (.I0(n31_adj_3920), .I1(n29_adj_14), .I2(n27_adj_13), 
            .I3(n48723), .O(n48175));
    defparam i32614_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_14_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33346_4_lut (.I0(n37_adj_3918), .I1(n35_adj_3927), .I2(n33_adj_3928), 
            .I3(n48175), .O(n48907));
    defparam i33346_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33196_3_lut (.I0(n6_adj_3937), .I1(n67[10]), .I2(n21_adj_3921), 
            .I3(GND_net), .O(n48757));   // verilog/motorControl.v(47[21:37])
    defparam i33196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33197_3_lut (.I0(n48757), .I1(n67[11]), .I2(n23_adj_3922), 
            .I3(GND_net), .O(n48758));   // verilog/motorControl.v(47[21:37])
    defparam i33197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_22_i16_3_lut (.I0(n67[9]), .I1(n399), .I2(n43), .I3(GND_net), 
            .O(n16_adj_3939));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_22_i8_3_lut (.I0(n67[4]), .I1(n67[8]), .I2(n17_adj_3924), 
            .I3(GND_net), .O(n8_adj_3940));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_22_i24_3_lut (.I0(n16_adj_3939), .I1(n67[22]), .I2(n45_adj_3917), 
            .I3(GND_net), .O(n24_adj_3941));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31267_4_lut (.I0(n21_adj_3921), .I1(n19_adj_3925), .I2(n17_adj_3924), 
            .I3(n9_adj_3926), .O(n46826));
    defparam i31267_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31234_4_lut (.I0(n43), .I1(n25_adj_3923), .I2(n23_adj_3922), 
            .I3(n46826), .O(n46793));
    defparam i31234_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33399_4_lut (.I0(n24_adj_3941), .I1(n8_adj_3940), .I2(n45_adj_3917), 
            .I3(n46791), .O(n48960));   // verilog/motorControl.v(47[21:37])
    defparam i33399_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32939_3_lut (.I0(n48758), .I1(n67[12]), .I2(n25_adj_3923), 
            .I3(GND_net), .O(n48500));   // verilog/motorControl.v(47[21:37])
    defparam i32939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_3_lut (.I0(\PID_CONTROLLER.result [30]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(n67[24]), .I3(GND_net), .O(n10_adj_3942));   // verilog/motorControl.v(47[21:37])
    defparam i3_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut (.I0(\PID_CONTROLLER.result [26]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(n67[24]), .I3(GND_net), .O(n8_adj_3943));   // verilog/motorControl.v(47[21:37])
    defparam i1_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i5_4_lut_adj_1372 (.I0(\PID_CONTROLLER.result [28]), .I1(n10_adj_3942), 
            .I2(\PID_CONTROLLER.result [25]), .I3(n67[24]), .O(n12_adj_3944));   // verilog/motorControl.v(47[21:37])
    defparam i5_4_lut_adj_1372.LUT_INIT = 16'hdffe;
    SB_LUT4 LessThan_22_i4_3_lut (.I0(n46593), .I1(n67[1]), .I2(\PID_CONTROLLER.result [1]), 
            .I3(GND_net), .O(n4_adj_3945));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33114_3_lut (.I0(n4_adj_3945), .I1(n407), .I2(n27_adj_13), 
            .I3(GND_net), .O(n48675));   // verilog/motorControl.v(47[21:37])
    defparam i33114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33115_3_lut (.I0(n48675), .I1(n406), .I2(n29_adj_14), .I3(GND_net), 
            .O(n48676));   // verilog/motorControl.v(47[21:37])
    defparam i33115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31252_4_lut (.I0(n33_adj_3928), .I1(n31_adj_3920), .I2(n29_adj_14), 
            .I3(n46817), .O(n46811));
    defparam i31252_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_21_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n60[20]));   // verilog/motorControl.v(47[28:37])
    defparam unary_minus_21_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33397_4_lut (.I0(n30_adj_3935), .I1(n10_adj_3934), .I2(n35_adj_3927), 
            .I3(n46807), .O(n48958));   // verilog/motorControl.v(47[21:37])
    defparam i33397_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32941_3_lut (.I0(n48676), .I1(n67[15]), .I2(n31_adj_3920), 
            .I3(GND_net), .O(n48502));   // verilog/motorControl.v(47[21:37])
    defparam i32941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33532_4_lut (.I0(n48502), .I1(n48958), .I2(n35_adj_3927), 
            .I3(n46811), .O(n49093));   // verilog/motorControl.v(47[21:37])
    defparam i33532_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33533_3_lut (.I0(n49093), .I1(n67[18]), .I2(n37_adj_3918), 
            .I3(GND_net), .O(n49094));   // verilog/motorControl.v(47[21:37])
    defparam i33533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33485_3_lut (.I0(n49094), .I1(n67[19]), .I2(n39_adj_3916), 
            .I3(GND_net), .O(n49046));   // verilog/motorControl.v(47[21:37])
    defparam i33485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31236_4_lut (.I0(n43), .I1(n41_adj_15), .I2(n39_adj_3916), 
            .I3(n48907), .O(n46795));
    defparam i31236_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33540_4_lut (.I0(n48500), .I1(n48960), .I2(n45_adj_3917), 
            .I3(n46793), .O(n49101));   // verilog/motorControl.v(47[21:37])
    defparam i33540_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33436_3_lut (.I0(n49046), .I1(n400), .I2(n41_adj_15), .I3(GND_net), 
            .O(n48997));   // verilog/motorControl.v(47[21:37])
    defparam i33436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33550_4_lut (.I0(n48997), .I1(n49101), .I2(n45_adj_3917), 
            .I3(n46795), .O(n49111));   // verilog/motorControl.v(47[21:37])
    defparam i33550_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6_4_lut (.I0(\PID_CONTROLLER.result [29]), .I1(n12_adj_3944), 
            .I2(n8_adj_3943), .I3(n67[24]), .O(n43881));   // verilog/motorControl.v(47[21:37])
    defparam i6_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 i33551_3_lut (.I0(n49111), .I1(n67[23]), .I2(\PID_CONTROLLER.result [23]), 
            .I3(GND_net), .O(n49112));   // verilog/motorControl.v(47[21:37])
    defparam i33551_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34256_4_lut (.I0(n49112), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n67[24]), .I3(n43881), .O(n49815));   // verilog/motorControl.v(47[21:37])
    defparam i34256_4_lut.LUT_INIT = 16'h3371;
    SB_LUT4 mult_10_i227_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n337));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n531_adj_3906));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3905));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_3904));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_3903));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n628_adj_3902));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_3901));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i487_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n725_adj_3900));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1373 (.I0(pwm_23__N_2957), .I1(n26834), .I2(PWMLimit[5]), 
            .I3(n387), .O(n24207));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1373.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1374 (.I0(pwm_23__N_2957), .I1(n1), .I2(PWMLimit[7]), 
            .I3(n387), .O(n24209));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1374.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1375 (.I0(pwm_23__N_2957), .I1(n2), .I2(PWMLimit[13]), 
            .I3(n387), .O(n24215));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1375.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1376 (.I0(pwm_23__N_2957), .I1(n27734), .I2(PWMLimit[14]), 
            .I3(n387), .O(n24216));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1376.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1377 (.I0(pwm_23__N_2957), .I1(n1_adj_3869), .I2(PWMLimit[20]), 
            .I3(n387), .O(n24222));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1377.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1378 (.I0(pwm_23__N_2957), .I1(n28362), .I2(PWMLimit[21]), 
            .I3(n387), .O(n24223));   // verilog/motorControl.v(44[10:51])
    defparam i1_4_lut_adj_1378.LUT_INIT = 16'ha088;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i37_2_lut  (.I0(deadband[18]), 
            .I1(\PID_CONTROLLER.result [18]), .I2(GND_net), .I3(GND_net), 
            .O(n37));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i37_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i39_2_lut  (.I0(deadband[19]), 
            .I1(\PID_CONTROLLER.result [19]), .I2(GND_net), .I3(GND_net), 
            .O(n39));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i39_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i31_2_lut  (.I0(deadband[15]), 
            .I1(\PID_CONTROLLER.result [15]), .I2(GND_net), .I3(GND_net), 
            .O(n31_adj_3406));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i31_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i162_2_lut (.I0(\Kd[2] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n240_adj_3899));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i7_2_lut  (.I0(deadband[3]), .I1(\PID_CONTROLLER.result [3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3948));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i7_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i35_2_lut  (.I0(deadband[17]), 
            .I1(\PID_CONTROLLER.result [17]), .I2(GND_net), .I3(GND_net), 
            .O(n35_adj_3416));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i35_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3898));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i33_2_lut  (.I0(deadband[16]), 
            .I1(\PID_CONTROLLER.result [16]), .I2(GND_net), .I3(GND_net), 
            .O(n33));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i33_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3897));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i142_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n210_adj_3896));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i207_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n307_adj_3895));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i13_2_lut  (.I0(deadband[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3949));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i13_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i93_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n137_adj_3894));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3893));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i272_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n404_adj_3892));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i337_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n501_adj_3891));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i158_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n234_adj_3890));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i45_2_lut  (.I0(deadband[22]), 
            .I1(\PID_CONTROLLER.result [22]), .I2(GND_net), .I3(GND_net), 
            .O(n45));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i45_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n598_adj_3889));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n695_adj_3887));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i23_2_lut  (.I0(deadband[11]), 
            .I1(\PID_CONTROLLER.result [11]), .I2(GND_net), .I3(GND_net), 
            .O(n23_adj_3950));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i23_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i25_2_lut  (.I0(deadband[12]), 
            .I1(\PID_CONTROLLER.result [12]), .I2(GND_net), .I3(GND_net), 
            .O(n25_c));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i25_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i223_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n331_adj_3885));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i288_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n428_adj_3884));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i9_2_lut  (.I0(deadband[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3951));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i9_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i17_2_lut  (.I0(deadband[8]), .I1(\PID_CONTROLLER.result [8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3952));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i17_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i19_2_lut  (.I0(deadband[9]), .I1(\PID_CONTROLLER.result [9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3953));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i19_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i21_2_lut  (.I0(deadband[10]), 
            .I1(\PID_CONTROLLER.result [10]), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_3954));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i21_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i39_2_lut (.I0(PWMLimit[19]), .I1(\PID_CONTROLLER.result [19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_3955));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i45_2_lut (.I0(PWMLimit[22]), .I1(\PID_CONTROLLER.result [22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_3956));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i37_2_lut (.I0(PWMLimit[18]), .I1(\PID_CONTROLLER.result [18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_3957));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i31_2_lut (.I0(PWMLimit[15]), .I1(\PID_CONTROLLER.result [15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_3958));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3883));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i23_2_lut (.I0(PWMLimit[11]), .I1(\PID_CONTROLLER.result [11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3959));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i25_2_lut (.I0(PWMLimit[12]), .I1(\PID_CONTROLLER.result [12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_3960));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_3882));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i35_2_lut (.I0(PWMLimit[17]), .I1(\PID_CONTROLLER.result [17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3961));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n525_adj_3881));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i33_2_lut (.I0(PWMLimit[16]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_3962));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i9_2_lut (.I0(PWMLimit[4]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3963));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i17_2_lut (.I0(PWMLimit[8]), .I1(\PID_CONTROLLER.result [8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3964));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i19_2_lut (.I0(PWMLimit[9]), .I1(\PID_CONTROLLER.result [9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3965));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i21_2_lut (.I0(PWMLimit[10]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_3966));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_20_i13_2_lut (.I0(PWMLimit[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_3967));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31334_4_lut (.I0(n21_adj_3966), .I1(n19_adj_3965), .I2(n17_adj_3964), 
            .I3(n9_adj_3963), .O(n46893));
    defparam i31334_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31328_4_lut (.I0(n27_adj_16), .I1(n15_adj_17), .I2(n13_adj_3967), 
            .I3(n11_adj_18), .O(n46887));
    defparam i31328_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_20_i30_3_lut (.I0(n12_adj_3971), .I1(\PID_CONTROLLER.result [17]), 
            .I2(n35_adj_3961), .I3(GND_net), .O(n30_adj_3972));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32116_4_lut (.I0(n13_adj_3967), .I1(n11_adj_18), .I2(n9_adj_3963), 
            .I3(n46916), .O(n47677));
    defparam i32116_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32112_4_lut (.I0(n19_adj_3965), .I1(n17_adj_3964), .I2(n15_adj_17), 
            .I3(n47677), .O(n47673));
    defparam i32112_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33184_4_lut (.I0(n25_adj_3960), .I1(n23_adj_3959), .I2(n21_adj_3966), 
            .I3(n47673), .O(n48745));
    defparam i33184_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32640_4_lut (.I0(n31_adj_3958), .I1(n29_adj_19), .I2(n27_adj_16), 
            .I3(n48745), .O(n48201));
    defparam i32640_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33350_4_lut (.I0(n37_adj_3957), .I1(n35_adj_3961), .I2(n33_adj_3962), 
            .I3(n48201), .O(n48911));
    defparam i33350_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33120_3_lut (.I0(n6_adj_3974), .I1(\PID_CONTROLLER.result [10]), 
            .I2(n21_adj_3966), .I3(GND_net), .O(n48681));   // verilog/motorControl.v(45[12:27])
    defparam i33120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33121_3_lut (.I0(n48681), .I1(\PID_CONTROLLER.result [11]), 
            .I2(n23_adj_3959), .I3(GND_net), .O(n48682));   // verilog/motorControl.v(45[12:27])
    defparam i33121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_20_i24_3_lut (.I0(n16_adj_3975), .I1(\PID_CONTROLLER.result [22]), 
            .I2(n45_adj_3956), .I3(GND_net), .O(n24_adj_3976));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31299_4_lut (.I0(n43_adj_20), .I1(n25_adj_3960), .I2(n23_adj_3959), 
            .I3(n46893), .O(n46858));
    defparam i31299_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32936_4_lut (.I0(n24_adj_3976), .I1(n8_adj_3978), .I2(n45_adj_3956), 
            .I3(n46854), .O(n48497));   // verilog/motorControl.v(45[12:27])
    defparam i32936_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32931_3_lut (.I0(n48682), .I1(\PID_CONTROLLER.result [12]), 
            .I2(n25_adj_3960), .I3(GND_net), .O(n48492));   // verilog/motorControl.v(45[12:27])
    defparam i32931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33118_3_lut (.I0(n4_adj_3979), .I1(\PID_CONTROLLER.result[13] ), 
            .I2(n27_adj_16), .I3(GND_net), .O(n48679));   // verilog/motorControl.v(45[12:27])
    defparam i33118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33119_3_lut (.I0(n48679), .I1(\PID_CONTROLLER.result[14] ), 
            .I2(n29_adj_19), .I3(GND_net), .O(n48680));   // verilog/motorControl.v(45[12:27])
    defparam i33119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31319_4_lut (.I0(n33_adj_3962), .I1(n31_adj_3958), .I2(n29_adj_19), 
            .I3(n46887), .O(n46878));
    defparam i31319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33395_4_lut (.I0(n30_adj_3972), .I1(n10_adj_3980), .I2(n35_adj_3961), 
            .I3(n46875), .O(n48956));   // verilog/motorControl.v(45[12:27])
    defparam i33395_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32933_3_lut (.I0(n48680), .I1(\PID_CONTROLLER.result [15]), 
            .I2(n31_adj_3958), .I3(GND_net), .O(n48494));   // verilog/motorControl.v(45[12:27])
    defparam i32933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33530_4_lut (.I0(n48494), .I1(n48956), .I2(n35_adj_3961), 
            .I3(n46878), .O(n49091));   // verilog/motorControl.v(45[12:27])
    defparam i33530_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33531_3_lut (.I0(n49091), .I1(\PID_CONTROLLER.result [18]), 
            .I2(n37_adj_3957), .I3(GND_net), .O(n49092));   // verilog/motorControl.v(45[12:27])
    defparam i33531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33487_3_lut (.I0(n49092), .I1(\PID_CONTROLLER.result [19]), 
            .I2(n39_adj_3955), .I3(GND_net), .O(n49048));   // verilog/motorControl.v(45[12:27])
    defparam i33487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31301_4_lut (.I0(n43_adj_20), .I1(n41_adj_21), .I2(n39_adj_3955), 
            .I3(n48911), .O(n46860));
    defparam i31301_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33192_4_lut (.I0(n48492), .I1(n48497), .I2(n45_adj_3956), 
            .I3(n46858), .O(n48753));   // verilog/motorControl.v(45[12:27])
    defparam i33192_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33434_3_lut (.I0(n49048), .I1(\PID_CONTROLLER.result[20] ), 
            .I2(n41_adj_21), .I3(GND_net), .O(n40_adj_3982));   // verilog/motorControl.v(45[12:27])
    defparam i33434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33194_4_lut (.I0(n40_adj_3982), .I1(n48753), .I2(n45_adj_3956), 
            .I3(n46860), .O(n48755));   // verilog/motorControl.v(45[12:27])
    defparam i33194_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33195_3_lut (.I0(n48755), .I1(\PID_CONTROLLER.result [23]), 
            .I2(PWMLimit[23]), .I3(GND_net), .O(n48_adj_3983));   // verilog/motorControl.v(45[12:27])
    defparam i33195_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i3_4_lut_adj_1379 (.I0(\PID_CONTROLLER.result [26]), .I1(n48_adj_3983), 
            .I2(\PID_CONTROLLER.result [24]), .I3(\PID_CONTROLLER.result [25]), 
            .O(n44079));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_1379.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1380 (.I0(\PID_CONTROLLER.result [26]), .I1(n48_adj_3983), 
            .I2(\PID_CONTROLLER.result [24]), .I3(\PID_CONTROLLER.result [25]), 
            .O(n44083));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_1380.LUT_INIT = 16'h8000;
    SB_LUT4 i3_4_lut_adj_1381 (.I0(\PID_CONTROLLER.result [30]), .I1(n56_adj_3984), 
            .I2(\PID_CONTROLLER.result [28]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n44134));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_1381.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1382 (.I0(\PID_CONTROLLER.result [30]), .I1(n56_adj_3984), 
            .I2(\PID_CONTROLLER.result [28]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n44139));   // verilog/motorControl.v(45[12:27])
    defparam i3_4_lut_adj_1382.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1383 (.I0(PWMLimit[23]), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n44139), .I3(n44134), .O(n387));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut_adj_1383.LUT_INIT = 16'hb3a2;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n622_adj_3880));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i227_2_lut (.I0(\Kd[3] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n337_adj_3879));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32369_3_lut (.I0(n25_c), .I1(n23_adj_3950), .I2(n21_adj_3954), 
            .I3(GND_net), .O(n47930));
    defparam i32369_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i32281_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [26]), 
            .I2(\PID_CONTROLLER.result [27]), .I3(n47930), .O(n47842));
    defparam i32281_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i31644_4_lut (.I0(n21_adj_3954), .I1(n19_adj_3953), .I2(n17_adj_3952), 
            .I3(n9_adj_3951), .O(n47205));
    defparam i31644_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31578_4_lut (.I0(n43_adj_22), .I1(n25_c), .I2(n23_adj_3950), 
            .I3(n47205), .O(n47139));
    defparam i31578_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32718_4_lut (.I0(deadband[23]), .I1(n45), .I2(\PID_CONTROLLER.result [23]), 
            .I3(n47139), .O(n48279));
    defparam i32718_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i33250_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\PID_CONTROLLER.result [25]), .I3(n48279), .O(n48811));
    defparam i33250_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32287_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [26]), 
            .I2(\PID_CONTROLLER.result [27]), .I3(n48811), .O(n47848));
    defparam i32287_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i31481_4_lut (.I0(\PID_CONTROLLER.result [6]), .I1(pwm_23__N_2960[5]), 
            .I2(pwm_23__N_2960[6]), .I3(\PID_CONTROLLER.result[5] ), .O(n47041));
    defparam i31481_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i32245_3_lut (.I0(pwm_23__N_2960[7]), .I1(n47041), .I2(\PID_CONTROLLER.result[7] ), 
            .I3(GND_net), .O(n47806));
    defparam i32245_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i32223_4_lut (.I0(\pwm_23__N_2960[14] ), .I1(n50261), .I2(\PID_CONTROLLER.result[14] ), 
            .I3(n47806), .O(n47784));
    defparam i32223_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 pwm_23__I_819_i31_rep_273_2_lut (.I0(\PID_CONTROLLER.result [15]), 
            .I1(pwm_23__N_2960[15]), .I2(GND_net), .I3(GND_net), .O(n50255));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i31_rep_273_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_819_i12_3_lut (.I0(pwm_23__N_2960[7]), .I1(pwm_23__N_2960[16]), 
            .I2(\PID_CONTROLLER.result [16]), .I3(GND_net), .O(n12_adj_3986));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31435_4_lut (.I0(\PID_CONTROLLER.result [16]), .I1(pwm_23__N_2960[7]), 
            .I2(pwm_23__N_2960[16]), .I3(\PID_CONTROLLER.result[7] ), .O(n46995));
    defparam i31435_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 pwm_23__I_819_i10_3_lut (.I0(pwm_23__N_2960[5]), .I1(pwm_23__N_2960[6]), 
            .I2(\PID_CONTROLLER.result [6]), .I3(GND_net), .O(n10));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 pwm_23__I_819_i30_3_lut (.I0(n12_adj_3986), .I1(pwm_23__N_2960[17]), 
            .I2(\PID_CONTROLLER.result [17]), .I3(GND_net), .O(n30_c));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i483_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n719_adj_3878));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31493_4_lut (.I0(\PID_CONTROLLER.result [3]), .I1(\PID_CONTROLLER.result [2]), 
            .I2(pwm_23__N_2960[3]), .I3(pwm_23__N_2960[2]), .O(n47053));
    defparam i31493_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 pwm_23__I_819_i9_rep_308_2_lut (.I0(\PID_CONTROLLER.result [4]), 
            .I1(pwm_23__N_2960[4]), .I2(GND_net), .I3(GND_net), .O(n50290));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i9_rep_308_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_14_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_3877));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31487_4_lut (.I0(pwm_23__N_2960[5]), .I1(n50290), .I2(\PID_CONTROLLER.result[5] ), 
            .I3(n47053), .O(n47047));
    defparam i31487_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 pwm_23__I_819_i13_rep_337_2_lut (.I0(\PID_CONTROLLER.result [6]), 
            .I1(pwm_23__N_2960[6]), .I2(GND_net), .I3(GND_net), .O(n50319));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i13_rep_337_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i24_4_lut (.I0(GATES_5__N_3048[4]), .I1(GATES_5__N_3048[5]), 
            .I2(n17_adj_3907), .I3(n878), .O(GATES_5__N_2788[5]));   // verilog/motorControl.v(86[14] 109[8])
    defparam i24_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i32688_4_lut (.I0(pwm_23__N_2960[7]), .I1(n50319), .I2(\PID_CONTROLLER.result[7] ), 
            .I3(n47047), .O(n48249));
    defparam i32688_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i2_4_lut_adj_1384 (.I0(hall1), .I1(GATES_5__N_3048[5]), .I2(hall2), 
            .I3(hall3), .O(GATES_5__N_3048[4]));   // verilog/motorControl.v(70[16] 85[10])
    defparam i2_4_lut_adj_1384.LUT_INIT = 16'h1050;
    SB_LUT4 GATES_5__I_0_i5_4_lut (.I0(n878), .I1(GATES_5__N_3048[4]), .I2(n17_adj_3907), 
            .I3(GATES_5__N_3048[5]), .O(GATES_5__N_2788[4]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i5_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 pwm_23__I_819_i17_rep_311_2_lut (.I0(\PID_CONTROLLER.result [8]), 
            .I1(pwm_23__N_2960[8]), .I2(GND_net), .I3(GND_net), .O(n50293));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i17_rep_311_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1385 (.I0(pwm_count[8]), .I1(n865), .I2(n868), 
            .I3(n16), .O(n19_adj_3988));
    defparam i3_4_lut_adj_1385.LUT_INIT = 16'h0223;
    SB_LUT4 i28798_3_lut (.I0(n866), .I1(n21), .I2(n853), .I3(GND_net), 
            .O(n44357));
    defparam i28798_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i28794_4_lut (.I0(n862), .I1(n864), .I2(n859), .I3(n861), 
            .O(n44353));
    defparam i28794_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28796_4_lut (.I0(n867), .I1(n863), .I2(n856), .I3(n860), 
            .O(n44355));
    defparam i28796_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32243_4_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n50293), 
            .I2(pwm_23__N_2960[9]), .I3(n48249), .O(n47804));
    defparam i32243_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i13_4_lut_adj_1386 (.I0(n44357), .I1(n19_adj_3988), .I2(n855), 
            .I3(n857), .O(n29_adj_3989));
    defparam i13_4_lut_adj_1386.LUT_INIT = 16'h0004;
    SB_LUT4 pwm_23__I_819_i21_rep_325_2_lut (.I0(\PID_CONTROLLER.result [10]), 
            .I1(pwm_23__N_2960[10]), .I2(GND_net), .I3(GND_net), .O(n50307));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i21_rep_325_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1387 (.I0(n29_adj_3989), .I1(hall3), .I2(n44355), 
            .I3(n44353), .O(n6_adj_3990));
    defparam i2_4_lut_adj_1387.LUT_INIT = 16'h333b;
    SB_LUT4 i33023_4_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n50307), 
            .I2(pwm_23__N_2960[11]), .I3(n47804), .O(n48584));
    defparam i33023_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 GATES_5__I_0_i4_4_lut (.I0(n5_adj_3549), .I1(GATES_5__N_3048[3]), 
            .I2(n17_adj_3907), .I3(n6_adj_3990), .O(GATES_5__N_2788[3]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i4_4_lut.LUT_INIT = 16'h0c5c;
    SB_LUT4 pwm_23__I_819_i25_rep_320_2_lut (.I0(\PID_CONTROLLER.result [12]), 
            .I1(pwm_23__N_2960[12]), .I2(GND_net), .I3(GND_net), .O(n50302));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i25_rep_320_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(hall2), .I1(GATES_5__N_3048[5]), .I2(hall3), 
            .I3(GND_net), .O(GATES_5__N_3048[3]));   // verilog/motorControl.v(70[16] 85[10])
    defparam i2_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i31450_4_lut (.I0(\pwm_23__N_2960[13] ), .I1(n50302), .I2(\PID_CONTROLLER.result[13] ), 
            .I3(n48584), .O(n47010));
    defparam i31450_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 GATES_5__I_0_i3_4_lut (.I0(n46652), .I1(hall2), .I2(n17_adj_3907), 
            .I3(hall3), .O(GATES_5__N_2788[2]));   // verilog/motorControl.v(86[14] 109[8])
    defparam GATES_5__I_0_i3_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 mult_12_i292_2_lut (.I0(\Kd[4] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n434_adj_3876));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32676_4_lut (.I0(\PID_CONTROLLER.result [15]), .I1(n50258), 
            .I2(pwm_23__N_2960[15]), .I3(n47010), .O(n48237));
    defparam i32676_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 unary_minus_17_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[0]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pwm_23__I_819_i33_rep_331_2_lut (.I0(\PID_CONTROLLER.result [16]), 
            .I1(pwm_23__N_2960[16]), .I2(GND_net), .I3(GND_net), .O(n50313));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i33_rep_331_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_17_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[1]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i357_2_lut (.I0(\Kd[5] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n531_adj_3872));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33232_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(n50313), 
            .I2(pwm_23__N_2960[17]), .I3(n48237), .O(n48793));
    defparam i33232_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_14_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_3871));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_819_i37_rep_267_2_lut (.I0(\PID_CONTROLLER.result [18]), 
            .I1(pwm_23__N_2960[18]), .I2(GND_net), .I3(GND_net), .O(n50249));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i37_rep_267_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33443_4_lut (.I0(\PID_CONTROLLER.result [19]), .I1(n50249), 
            .I2(pwm_23__N_2960[19]), .I3(n48793), .O(n49004));
    defparam i33443_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 pwm_23__I_819_i16_3_lut (.I0(pwm_23__N_2960[9]), .I1(pwm_23__N_2960[21]), 
            .I2(\PID_CONTROLLER.result[21] ), .I3(GND_net), .O(n16_adj_3991));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31390_4_lut (.I0(pwm_23__N_2960[21]), .I1(\PID_CONTROLLER.result [9]), 
            .I2(\PID_CONTROLLER.result[21] ), .I3(pwm_23__N_2960[9]), .O(n46950));
    defparam i31390_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 pwm_23__I_819_i8_3_lut (.I0(pwm_23__N_2960[4]), .I1(pwm_23__N_2960[8]), 
            .I2(\PID_CONTROLLER.result [8]), .I3(GND_net), .O(n8_adj_3992));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 pwm_23__I_819_i24_3_lut (.I0(n16_adj_3991), .I1(pwm_23__N_2960[22]), 
            .I2(\PID_CONTROLLER.result [22]), .I3(GND_net), .O(n24_adj_3993));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_17_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[2]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31471_4_lut (.I0(\PID_CONTROLLER.result [8]), .I1(\PID_CONTROLLER.result [4]), 
            .I2(pwm_23__N_2960[8]), .I3(pwm_23__N_2960[4]), .O(n47031));
    defparam i31471_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i32239_3_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n47031), 
            .I2(pwm_23__N_2960[9]), .I3(GND_net), .O(n47800));
    defparam i32239_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 pwm_23__I_819_i6_3_lut (.I0(pwm_23__N_2960[2]), .I1(pwm_23__N_2960[3]), 
            .I2(\PID_CONTROLLER.result [3]), .I3(GND_net), .O(n6_adj_3994));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32898_3_lut (.I0(n6_adj_3994), .I1(pwm_23__N_2960[10]), .I2(\PID_CONTROLLER.result [10]), 
            .I3(GND_net), .O(n48459));   // verilog/motorControl.v(44[31:51])
    defparam i32898_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i79_2_lut (.I0(\Kd[1] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_3868));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32899_3_lut (.I0(n48459), .I1(pwm_23__N_2960[11]), .I2(\PID_CONTROLLER.result [11]), 
            .I3(GND_net), .O(n48460));   // verilog/motorControl.v(44[31:51])
    defparam i32899_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i16_2_lut (.I0(\Kd[0] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3867));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32235_4_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n50307), 
            .I2(pwm_23__N_2960[11]), .I3(n47800), .O(n47796));
    defparam i32235_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i31393_4_lut (.I0(pwm_23__N_2960[21]), .I1(n50302), .I2(\PID_CONTROLLER.result[21] ), 
            .I3(n47796), .O(n46953));
    defparam i31393_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_12_i422_2_lut (.I0(\Kd[6] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n628));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 pwm_23__I_819_i45_rep_257_2_lut (.I0(\PID_CONTROLLER.result [22]), 
            .I1(pwm_23__N_2960[22]), .I2(GND_net), .I3(GND_net), .O(n50239));   // verilog/motorControl.v(44[31:51])
    defparam pwm_23__I_819_i45_rep_257_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33393_4_lut (.I0(n24_adj_3993), .I1(n8_adj_3992), .I2(n50239), 
            .I3(n46950), .O(n48954));   // verilog/motorControl.v(44[31:51])
    defparam i33393_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32103_3_lut (.I0(n48460), .I1(pwm_23__N_2960[12]), .I2(\PID_CONTROLLER.result [12]), 
            .I3(GND_net), .O(n47664));   // verilog/motorControl.v(44[31:51])
    defparam i32103_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31626_4_lut (.I0(n27), .I1(n15_adj_23), .I2(n13_adj_3949), 
            .I3(n11_adj_24), .O(n47187));
    defparam i31626_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i30_3_lut  (.I0(n12_adj_3997), 
            .I1(\PID_CONTROLLER.result [17]), .I2(n35_adj_3416), .I3(GND_net), 
            .O(n30_adj_3414));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i32399_4_lut (.I0(n9_adj_3951), .I1(n7_adj_3948), .I2(deadband[2]), 
            .I3(\PID_CONTROLLER.result [2]), .O(n47960));
    defparam i32399_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i32762_4_lut (.I0(n15_adj_23), .I1(n13_adj_3949), .I2(n11_adj_24), 
            .I3(n47960), .O(n48323));
    defparam i32762_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32756_4_lut (.I0(n21_adj_3954), .I1(n19_adj_3953), .I2(n17_adj_3952), 
            .I3(n48323), .O(n48317));
    defparam i32756_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31630_4_lut (.I0(n27), .I1(n25_c), .I2(n23_adj_3950), .I3(n48317), 
            .O(n47191));
    defparam i31630_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33049_4_lut (.I0(n33), .I1(n31_adj_3406), .I2(n29), .I3(n47191), 
            .O(n48610));
    defparam i33049_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33464_4_lut (.I0(n39), .I1(n37), .I2(n35_adj_3416), .I3(n48610), 
            .O(n49025));
    defparam i33464_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32317_4_lut (.I0(n45), .I1(n43_adj_22), .I2(n41), .I3(n49025), 
            .O(n47878));
    defparam i32317_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33039_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [23]), 
            .I2(\PID_CONTROLLER.result [24]), .I3(n47878), .O(n48600));
    defparam i33039_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33381_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [25]), 
            .I2(\PID_CONTROLLER.result [26]), .I3(n48600), .O(n48942));
    defparam i33381_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33520_4_lut (.I0(deadband[23]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\PID_CONTROLLER.result [28]), .I3(n48942), .O(n49081));
    defparam i33520_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i31357_3_lut_4_lut (.I0(PWMLimit[3]), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(PWMLimit[2]), .O(n46916));   // verilog/motorControl.v(45[12:27])
    defparam i31357_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i5_4_lut_adj_1388 (.I0(Kd_delay_counter[5]), .I1(Kd_delay_counter[3]), 
            .I2(Kd_delay_counter[6]), .I3(Kd_delay_counter[4]), .O(n12_adj_3998));   // verilog/motorControl.v(56[10:29])
    defparam i5_4_lut_adj_1388.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1389 (.I0(Kd_delay_counter[1]), .I1(n12_adj_3998), 
            .I2(Kd_delay_counter[2]), .I3(Kd_delay_counter[0]), .O(n43357));   // verilog/motorControl.v(56[10:29])
    defparam i6_4_lut_adj_1389.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_20_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(GND_net), .O(n6_adj_3974));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3866));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3865));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i140_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n207_adj_3864));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i2_2_lut (.I0(\Kd[0] ), .I1(n69[0]), .I2(GND_net), 
            .I3(GND_net), .O(n191[0]));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i205_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n304_adj_3863));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i144_2_lut (.I0(\Kd[2] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n213_adj_3862));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i270_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n401_adj_3861));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i97_2_lut (.I0(\Kd[1] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n143));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i487_2_lut (.I0(\Kd[7] ), .I1(n69[15]), .I2(GND_net), 
            .I3(GND_net), .O(n725));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i335_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n498_adj_3860));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i6_3_lut_3_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n67[3]), 
            .I2(n67[2]), .I3(GND_net), .O(n6_adj_3937));   // verilog/motorControl.v(47[21:37])
    defparam LessThan_22_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i31292_3_lut_4_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n67[3]), 
            .I2(n67[2]), .I3(\PID_CONTROLLER.result [2]), .O(n46851));   // verilog/motorControl.v(47[21:37])
    defparam i31292_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n595_adj_3859));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i34_2_lut (.I0(\Kd[0] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[3]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3857));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3856));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3854));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3852));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n692_adj_3850));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[4]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i209_2_lut (.I0(\Kd[3] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n310_adj_3846));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_3845));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[5]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i113_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n167_adj_3839));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[6]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i178_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n264_adj_3837));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i274_2_lut (.I0(\Kd[4] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n407_adj_3836));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i339_2_lut (.I0(\Kd[5] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n504_adj_3835));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[7]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i243_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n361_adj_3833));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[8]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n458_adj_3831));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[9]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i404_2_lut (.I0(\Kd[6] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n601_adj_3829));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n555_adj_3828));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i469_2_lut (.I0(\Kd[7] ), .I1(n69[6]), .I2(GND_net), 
            .I3(GND_net), .O(n698_adj_3827));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i438_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n652_adj_3826));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i503_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_3825));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[10]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3820));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_3819));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[11]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[12]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[13]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i95_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n140_adj_3814));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3813));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[14]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3811));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[15]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[16]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3807));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3806));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_3805));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[17]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i203_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n301_adj_3803));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i268_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n398_adj_3802));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22241_3_lut_4_lut (.I0(n10844[2]), .I1(\Kd[4] ), .I2(n69[25]), 
            .I3(n6_adj_3999), .O(n8_adj_4000));   // verilog/motorControl.v(43[26:45])
    defparam i22241_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kd[5] ), .I1(n69[25]), .I2(\Kd[4] ), 
            .I3(n6_adj_3999), .O(n8_adj_4001));   // verilog/motorControl.v(43[26:45])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hb748;
    SB_LUT4 i22200_3_lut_4_lut (.I0(n10844[1]), .I1(\Kd[3] ), .I2(n69[25]), 
            .I3(n4_adj_3545), .O(n6_adj_3999));   // verilog/motorControl.v(43[26:45])
    defparam i22200_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i22137_2_lut_3_lut (.I0(\Kd[0] ), .I1(n69[25]), .I2(\Kd[1] ), 
            .I3(GND_net), .O(n35689));   // verilog/motorControl.v(43[26:45])
    defparam i22137_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_1390 (.I0(n10844[2]), .I1(\Kd[4] ), .I2(n69[25]), 
            .I3(n6_adj_3999), .O(n10109[3]));   // verilog/motorControl.v(43[26:45])
    defparam i1_3_lut_4_lut_adj_1390.LUT_INIT = 16'h956a;
    SB_LUT4 LessThan_4_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4002));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i333_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n495_adj_3801));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[18]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i160_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n237_adj_3799));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n592_adj_3798));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n689_adj_3797));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[19]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[20]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[21]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i225_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n334_adj_3793));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31574_2_lut_4_lut (.I0(deadband[21]), .I1(\PID_CONTROLLER.result[21] ), 
            .I2(deadband[9]), .I3(\PID_CONTROLLER.result [9]), .O(n47135));
    defparam i31574_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_14_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_3792));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i290_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n431_adj_3789));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i99_2_lut (.I0(\Kd[1] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n146_adj_3786));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i36_2_lut (.I0(\Kd[0] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_3785));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i16_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [9]), 
            .I1(\PID_CONTROLLER.result[21] ), .I2(deadband[21]), .I3(GND_net), 
            .O(n16_c));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i16_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i164_2_lut (.I0(\Kd[2] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n243_adj_3784));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n528_adj_3783));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[22]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n58[0]));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n282[0]));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[5] ), 
            .I1(\PID_CONTROLLER.result [6]), .I2(deadband[6]), .I3(GND_net), 
            .O(n10_adj_3415));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 i31606_2_lut_4_lut (.I0(deadband[16]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(deadband[7]), .I3(\PID_CONTROLLER.result[7] ), .O(n47167));
    defparam i31606_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i12_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[7] ), 
            .I1(\PID_CONTROLLER.result [16]), .I2(deadband[16]), .I3(GND_net), 
            .O(n12_adj_3997));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i12_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_12_i229_2_lut (.I0(\Kd[3] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n340_adj_3779));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31458_2_lut_4_lut (.I0(hall2), .I1(GATES_5__N_3048[5]), .I2(hall3), 
            .I3(n878), .O(n46652));   // verilog/motorControl.v(86[14] 109[8])
    defparam i31458_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 mult_14_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3778));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i32_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[31]));   // verilog/motorControl.v(44[41:50])
    defparam unary_minus_17_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i111_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n164_adj_3776));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i48_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n71_adj_3775));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i176_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n261_adj_3774));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i241_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n358_adj_3773));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i294_2_lut (.I0(\Kd[4] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n437_adj_3772));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i359_2_lut (.I0(\Kd[5] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n534_adj_3771));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n455_adj_3770));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_3769));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n552_adj_3768));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i105_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n155_adj_3767));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_3766));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n625_adj_3765));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i424_2_lut (.I0(\Kd[6] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n631_adj_3764));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i170_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n252_adj_3763));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[0]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i489_2_lut (.I0(\Kd[7] ), .I1(n69[16]), .I2(GND_net), 
            .I3(GND_net), .O(n728_adj_3760));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[1]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i436_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n649_adj_3757));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i485_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n722_adj_3756));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i501_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_3755));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[2]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i235_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n349_adj_3752));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n446_adj_3751));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_3750));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i91_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n134_adj_3748));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3747));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[3]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[4]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i156_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n231_adj_3742));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i81_2_lut (.I0(\Kd[1] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_3741));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i18_2_lut (.I0(\Kd[0] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_3740));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[5]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_3737));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i221_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n328_adj_3735));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[6]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_4_lut_adj_1391 (.I0(\PID_CONTROLLER.result [27]), .I1(PWMLimit[23]), 
            .I2(n44083), .I3(n44079), .O(n56_adj_3984));   // verilog/motorControl.v(45[12:27])
    defparam i1_4_lut_4_lut_adj_1391.LUT_INIT = 16'hb3a2;
    SB_LUT4 mult_10_i286_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n425_adj_3732));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_20_i4_4_lut_4_lut (.I0(\PID_CONTROLLER.result [0]), .I1(\PID_CONTROLLER.result [1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_3979));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i4_4_lut_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 LessThan_20_i8_3_lut_3_lut (.I0(\PID_CONTROLLER.result [4]), .I1(\PID_CONTROLLER.result [8]), 
            .I2(PWMLimit[8]), .I3(GND_net), .O(n8_adj_3978));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31295_2_lut_4_lut (.I0(PWMLimit[21]), .I1(\PID_CONTROLLER.result[21] ), 
            .I2(PWMLimit[9]), .I3(\PID_CONTROLLER.result [9]), .O(n46854));
    defparam i31295_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_20_i16_3_lut_3_lut (.I0(\PID_CONTROLLER.result [9]), 
            .I1(\PID_CONTROLLER.result[21] ), .I2(PWMLimit[21]), .I3(GND_net), 
            .O(n16_adj_3975));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_20_i10_3_lut_3_lut (.I0(\PID_CONTROLLER.result[5] ), 
            .I1(\PID_CONTROLLER.result [6]), .I2(PWMLimit[6]), .I3(GND_net), 
            .O(n10_adj_3980));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31316_2_lut_4_lut (.I0(PWMLimit[16]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(PWMLimit[7]), .I3(\PID_CONTROLLER.result[7] ), .O(n46875));
    defparam i31316_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_20_i12_3_lut_3_lut (.I0(\PID_CONTROLLER.result[7] ), 
            .I1(\PID_CONTROLLER.result [16]), .I2(PWMLimit[16]), .I3(GND_net), 
            .O(n12_adj_3971));   // verilog/motorControl.v(45[12:27])
    defparam LessThan_20_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15417_1_lut (.I0(pwm_count[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n28817));   // verilog/motorControl.v(110[18:29])
    defparam i15417_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i1_1_lut (.I0(pwm[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[0]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3730));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3729));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n522_adj_3728));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i2_1_lut (.I0(pwm[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[1]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31232_2_lut_4_lut (.I0(n399), .I1(\PID_CONTROLLER.result[21] ), 
            .I2(\PID_CONTROLLER.result [9]), .I3(n67[9]), .O(n46791));
    defparam i31232_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i4_2_lut (.I0(n19_adj_3683), .I1(n25_adj_3634), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4003));   // verilog/motorControl.v(40[38:63])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n33_adj_3607), .I1(n43_adj_3566), .I2(n27_adj_3626), 
            .I3(n35_adj_3603), .O(n24_adj_4004));   // verilog/motorControl.v(40[38:63])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n41_adj_3576), .I1(n45_adj_3539), .I2(n31_adj_3609), 
            .I3(n23_adj_3640), .O(n22_adj_4005));   // verilog/motorControl.v(40[38:63])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n29_adj_3612), .I1(n24_adj_4004), .I2(n18_adj_4003), 
            .I3(n37_adj_3594), .O(n26_adj_4006));   // verilog/motorControl.v(40[38:63])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1392 (.I0(n21_adj_3669), .I1(n26_adj_4006), .I2(n22_adj_4005), 
            .I3(n39_adj_3590), .O(n43653));   // verilog/motorControl.v(40[38:63])
    defparam i13_4_lut_adj_1392.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_4_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(IntegralLimit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4007));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(IntegralLimit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4008));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(IntegralLimit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4009));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32495_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4009), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4008), .O(n48056));
    defparam i32495_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32493_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[10]), 
            .I2(IntegralLimit[11]), .I3(n48056), .O(n48054));
    defparam i32493_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i31696_4_lut (.I0(n11_adj_3738), .I1(n9_adj_3743), .I2(n7_adj_3745), 
            .I3(n5_adj_3753), .O(n47257));
    defparam i31696_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_4_i13_rep_559_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n50541));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i13_rep_559_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32509_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n50541), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4007), .O(n48070));
    defparam i32509_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32477_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n48070), .O(n48038));
    defparam i32477_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i31742_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n47303));
    defparam i31742_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_4_i35_rep_547_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n50529));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i35_rep_547_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31248_2_lut_4_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n67[16]), 
            .I2(n413), .I3(\PID_CONTROLLER.result[7] ), .O(n46807));
    defparam i31248_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_4_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4010));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_4_i30_4_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[16]), .O(n30_adj_4011));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_4_i5_2_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(IntegralLimit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4012));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32499_4_lut (.I0(n9_adj_4008), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n5_adj_4012), .I3(IntegralLimit[3]), .O(n48060));
    defparam i32499_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i31797_4_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n11_adj_4007), 
            .I2(IntegralLimit[6]), .I3(n48060), .O(n47358));
    defparam i31797_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i31789_4_lut (.I0(n17_adj_4009), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n47358), .I3(IntegralLimit[7]), .O(n47350));
    defparam i31789_4_lut.LUT_INIT = 16'haeab;
    SB_LUT4 i32808_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[9]), 
            .I2(IntegralLimit[10]), .I3(n47350), .O(n48369));
    defparam i32808_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33282_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[11]), 
            .I2(IntegralLimit[12]), .I3(n48369), .O(n48843));
    defparam i33282_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32483_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n48843), .O(n48044));
    defparam i32483_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i33067_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n48044), .O(n48628));
    defparam i33067_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33389_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[17]), 
            .I2(IntegralLimit[18]), .I3(n48628), .O(n48950));
    defparam i33389_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33524_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[19]), 
            .I2(IntegralLimit[20]), .I3(n48950), .O(n49085));
    defparam i33524_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_4_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4013));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31899_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(IntegralLimit[9]), .O(n47460));
    defparam i31899_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 LessThan_4_i24_4_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[21]), .O(n24_adj_4014));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i24_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i32920_3_lut (.I0(n6_adj_4013), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48481));   // verilog/motorControl.v(40[10:34])
    defparam i32920_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31714_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[12]), 
            .I2(IntegralLimit[21]), .I3(n48054), .O(n47275));
    defparam i31714_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_4_i45_rep_512_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n50494));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i45_rep_512_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32924_3_lut (.I0(n24_adj_4014), .I1(n8_adj_4002), .I2(n47460), 
            .I3(GND_net), .O(n48485));   // verilog/motorControl.v(40[10:34])
    defparam i32924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32077_4_lut (.I0(n48481), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[11]), .O(n47638));   // verilog/motorControl.v(40[10:34])
    defparam i32077_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_6_i4_4_lut (.I0(n73[0]), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3_adj_3758), .I3(\PID_CONTROLLER.integral [0]), .O(n4_adj_4015));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i4_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i32914_3_lut (.I0(n4_adj_4015), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n11_adj_3738), .I3(GND_net), .O(n48475));   // verilog/motorControl.v(40[38:63])
    defparam i32914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32915_3_lut (.I0(n48475), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n13_adj_3733), .I3(GND_net), .O(n48476));   // verilog/motorControl.v(40[38:63])
    defparam i32915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i8_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n17_adj_3698), .I3(GND_net), .O(n8_adj_4016));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31680_2_lut (.I0(n17_adj_3698), .I1(n9_adj_3743), .I2(GND_net), 
            .I3(GND_net), .O(n47241));
    defparam i31680_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_6_i6_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n7_adj_3745), .I3(GND_net), .O(n6_adj_4017));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i16_3_lut (.I0(n8_adj_4016), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n43653), .I3(GND_net), .O(n16_adj_4018));   // verilog/motorControl.v(40[38:63])
    defparam LessThan_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31686_4_lut (.I0(n17_adj_3698), .I1(n15_adj_3702), .I2(n13_adj_3733), 
            .I3(n47257), .O(n47247));
    defparam i31686_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33021_4_lut (.I0(n16_adj_4018), .I1(n6_adj_4017), .I2(n43653), 
            .I3(n47241), .O(n48582));   // verilog/motorControl.v(40[38:63])
    defparam i33021_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32087_3_lut (.I0(n48476), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n15_adj_3702), .I3(GND_net), .O(n47648));   // verilog/motorControl.v(40[38:63])
    defparam i32087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33354_4_lut (.I0(n47648), .I1(n48582), .I2(n43653), .I3(n47247), 
            .O(n48915));   // verilog/motorControl.v(40[38:63])
    defparam i33354_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_4_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(IntegralLimit[1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), .O(n4_adj_4019));   // verilog/motorControl.v(40[10:34])
    defparam LessThan_4_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i32918_3_lut (.I0(n4_adj_4019), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48479));   // verilog/motorControl.v(40[10:34])
    defparam i32918_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31746_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n48038), .O(n47307));
    defparam i31746_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i33314_4_lut (.I0(n30_adj_4011), .I1(n10_adj_4010), .I2(n50529), 
            .I3(n47303), .O(n48875));   // verilog/motorControl.v(40[10:34])
    defparam i33314_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32079_4_lut (.I0(n48479), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[14]), .O(n47640));   // verilog/motorControl.v(40[10:34])
    defparam i32079_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33488_4_lut (.I0(n47640), .I1(n48875), .I2(n50529), .I3(n47307), 
            .O(n49049));   // verilog/motorControl.v(40[10:34])
    defparam i33488_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33489_3_lut (.I0(n49049), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n49050));   // verilog/motorControl.v(40[10:34])
    defparam i33489_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32441_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(n49085), .O(n48002));
    defparam i32441_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i33186_4_lut (.I0(n47638), .I1(n48485), .I2(n50494), .I3(n47275), 
            .O(n48747));   // verilog/motorControl.v(40[10:34])
    defparam i33186_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32085_4_lut (.I0(n49050), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[19]), .O(n47646));   // verilog/motorControl.v(40[10:34])
    defparam i32085_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33355_3_lut (.I0(n48915), .I1(n73[23]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48916));   // verilog/motorControl.v(40[38:63])
    defparam i33355_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33352_3_lut (.I0(n47646), .I1(n48747), .I2(n48002), .I3(GND_net), 
            .O(n48913));   // verilog/motorControl.v(40[10:34])
    defparam i33352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1393 (.I0(n48913), .I1(n48916), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[23]), .O(n55_adj_3726));   // verilog/motorControl.v(40[10:63])
    defparam i8_4_lut_adj_1393.LUT_INIT = 16'h80c8;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n543_adj_3725));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i3_1_lut (.I0(pwm[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[2]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i430_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n640_adj_3723));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i136_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n201_adj_3722));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i201_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n298_adj_3721));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n619_adj_3720));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i481_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n716_adj_3719));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i266_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n395_adj_3718));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i146_2_lut (.I0(\Kd[2] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n216_adj_3717));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i211_2_lut (.I0(\Kd[3] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n313_adj_3716));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i276_2_lut (.I0(\Kd[4] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n410_adj_3715));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i341_2_lut (.I0(\Kd[5] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n507_adj_3714));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i495_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_3713));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i406_2_lut (.I0(\Kd[6] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n604_adj_3712));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_c));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i471_2_lut (.I0(\Kd[7] ), .I1(n69[7]), .I2(GND_net), 
            .I3(GND_net), .O(n701_adj_3709));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i4_1_lut (.I0(pwm[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[3]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i331_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n492_adj_3707));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n589_adj_3706));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i5_1_lut (.I0(pwm[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[4]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n686_adj_3704));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[7]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i6_1_lut (.I0(pwm[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[5]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[8]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i101_2_lut (.I0(\Kd[1] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n149_adj_3697));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i38_2_lut (.I0(\Kd[0] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_3696));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i7_1_lut (.I0(pwm[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[6]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i103_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n152_adj_3694));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i40_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n59_adj_3693));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i168_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n249_adj_3692));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i166_2_lut (.I0(\Kd[2] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n246_adj_3691));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i231_2_lut (.I0(\Kd[3] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n343_adj_3690));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i296_2_lut (.I0(\Kd[4] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n440_adj_3689));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i233_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n346_adj_3688));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i361_2_lut (.I0(\Kd[5] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n537_adj_3687));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n443_adj_3686));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i8_1_lut (.I0(pwm[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[7]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[9]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i426_2_lut (.I0(\Kd[6] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n634_adj_3682));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_3681));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3680));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i154_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n228_adj_3679));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i219_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n325_adj_3678));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n540_adj_3677));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i491_2_lut (.I0(\Kd[7] ), .I1(n69[17]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_3676));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i9_1_lut (.I0(pwm[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[8]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3674));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3673));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i284_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n422_adj_3672));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i428_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n637_adj_3671));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[10]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n519_adj_3668));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n616_adj_3667));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i10_1_lut (.I0(pwm[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n76[9]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i479_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n713_adj_3665));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3664));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3663));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3662));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i199_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n295_adj_3661));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i83_2_lut (.I0(\Kd[1] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_3660));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i20_2_lut (.I0(\Kd[0] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3659));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i264_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n392_adj_3658));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i329_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n489_adj_3657));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i329_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n586_adj_3656));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n683_adj_3655));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i148_2_lut (.I0(\Kd[2] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n219_adj_3654));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_3653));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i493_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_3652));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_3651));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i109_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n161_adj_3649));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i46_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n68_adj_3648));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i174_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n258_adj_3647));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i239_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n355_adj_3646));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i213_2_lut (.I0(\Kd[3] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n316_adj_3645));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n452_adj_3644));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i278_2_lut (.I0(\Kd[4] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n413_adj_3643));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i343_2_lut (.I0(\Kd[5] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n510_adj_3642));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[11]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i408_2_lut (.I0(\Kd[6] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n607_adj_3638));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n549_adj_3637));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i11_1_lut (.I0(pwm[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[10]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[12]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i434_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n646_adj_3633));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i473_2_lut (.I0(\Kd[7] ), .I1(n69[8]), .I2(GND_net), 
            .I3(GND_net), .O(n704_adj_3632));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i499_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_3631));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i12_1_lut (.I0(pwm[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[11]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i13_1_lut (.I0(pwm[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[12]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i14_1_lut (.I0(pwm[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[13]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[13]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i87_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n128_adj_3625));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3624));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i152_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n225_adj_3623));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i15_1_lut (.I0(pwm[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[14]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i217_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n322_adj_3621));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i282_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n419_adj_3620));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i16_1_lut (.I0(pwm[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[15]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n516_adj_3618));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n613_adj_3617));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i477_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n710_adj_3616));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i17_1_lut (.I0(pwm[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[16]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[14]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i18_1_lut (.I0(pwm[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[17]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[15]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[16]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i19_1_lut (.I0(pwm[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[18]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i20_1_lut (.I0(pwm[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[19]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[17]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i21_1_lut (.I0(pwm[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[20]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i103_2_lut (.I0(\Kd[1] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n152_adj_3601));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i40_2_lut (.I0(\Kd[0] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i22_1_lut (.I0(pwm[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[21]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i23_1_lut (.I0(pwm[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[22]));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3597));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3596));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[18]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i24_1_lut (.I0(pwm[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(GATES_5__N_3055));   // verilog/motorControl.v(86[38:44])
    defparam unary_minus_70_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3593));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[19]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3589));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3588));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i197_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n292_adj_3587));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i150_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n222_adj_3585));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i168_2_lut (.I0(\Kd[2] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n249));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i262_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n389_adj_3583));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i1_1_lut (.I0(\PID_CONTROLLER.err[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[0]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i327_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n486_adj_3581));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i233_2_lut (.I0(\Kd[3] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n346));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i215_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n319_adj_3580));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i392_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n583_adj_3579));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[20]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i280_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n416_adj_3575));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n680_adj_3574));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i298_2_lut (.I0(\Kd[4] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n443_adj_3572));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i2_1_lut (.I0(\PID_CONTROLLER.err[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[1]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n513_adj_3570));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i3_1_lut (.I0(\PID_CONTROLLER.err[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[2]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[21]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i363_2_lut (.I0(\Kd[5] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n540));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i117_2_lut (.I0(\Kd[1] ), .I1(n69[25]), .I2(GND_net), 
            .I3(GND_net), .O(n182_adj_3565));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i117_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i182_2_lut (.I0(\Kd[2] ), .I1(n69[25]), .I2(GND_net), 
            .I3(GND_net), .O(n276_adj_3564));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i182_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i85_2_lut (.I0(\Kd[1] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i22_2_lut (.I0(\Kd[0] ), .I1(n69[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_3562));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i428_2_lut (.I0(\Kd[6] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n637));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i101_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n149));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i150_2_lut (.I0(\Kd[2] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n222_adj_3560));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i493_2_lut (.I0(\Kd[7] ), .I1(n69[18]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n610_adj_3559));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i215_2_lut (.I0(\Kd[3] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n319));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i166_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n246_adj_3558));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i280_2_lut (.I0(\Kd[4] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n416_adj_3557));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i345_2_lut (.I0(\Kd[5] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n513));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i231_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n343));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3555));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3554));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1394 (.I0(\Kd[2] ), .I1(\Kd[0] ), .I2(n69[25]), 
            .I3(\Kd[1] ), .O(n4_adj_3545));   // verilog/motorControl.v(43[26:45])
    defparam i2_4_lut_adj_1394.LUT_INIT = 16'ha080;
    SB_LUT4 mult_12_i247_2_lut (.I0(\Kd[3] ), .I1(n69[25]), .I2(GND_net), 
            .I3(GND_net), .O(n370_adj_3544));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22161_3_lut (.I0(n69[25]), .I1(n35689), .I2(n35704), .I3(GND_net), 
            .O(n10844[1]));   // verilog/motorControl.v(43[26:45])
    defparam i22161_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_12_i312_2_lut (.I0(\Kd[4] ), .I1(n69[25]), .I2(GND_net), 
            .I3(GND_net), .O(n464_adj_3563));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i379_2_lut (.I0(\Kd[5] ), .I1(n69[25]), .I2(GND_net), 
            .I3(GND_net), .O(n564));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i379_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i442_2_lut (.I0(\Kd[6] ), .I1(n69[25]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_3553));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1395 (.I0(n35689), .I1(n7_adj_3546), .I2(n8_adj_4000), 
            .I3(n8_adj_4001), .O(n43988));   // verilog/motorControl.v(43[26:45])
    defparam i5_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i475_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n707_adj_3552));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i410_2_lut (.I0(\Kd[6] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n610));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n440));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i475_2_lut (.I0(\Kd[7] ), .I1(n69[9]), .I2(GND_net), 
            .I3(GND_net), .O(n707));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [4]), 
            .I1(\PID_CONTROLLER.result [8]), .I2(deadband[8]), .I3(GND_net), 
            .O(n8));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n4_adj_4020), .I3(n37873), .O(n7_adj_3822));   // verilog/motorControl.v(43[17:23])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h78b4;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n4_adj_4020), .I3(n16635[1]), .O(n16635[2]));   // verilog/motorControl.v(43[17:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_12_i105_2_lut (.I0(\Kd[1] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i42_2_lut (.I0(\Kd[0] ), .I1(n69[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i170_2_lut (.I0(\Kd[2] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n252));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n537));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i235_2_lut (.I0(\Kd[3] ), .I1(n69[19]), .I2(GND_net), 
            .I3(GND_net), .O(n349));   // verilog/motorControl.v(43[26:45])
    defparam mult_12_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i426_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n634));   // verilog/motorControl.v(43[17:23])
    defparam mult_10_i426_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_3543));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i4_1_lut (.I0(\PID_CONTROLLER.err[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[3]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[22]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_3538));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i5_1_lut (.I0(\PID_CONTROLLER.err[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[4]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(43[48:59])
    defparam mult_14_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21934_3_lut_4_lut (.I0(n16635[2]), .I1(\Kp[4] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n6_adj_4021), .O(n8_adj_3823));   // verilog/motorControl.v(43[17:23])
    defparam i21934_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_3_lut_4_lut_adj_1396 (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[4] ), .I3(n6_adj_4021), .O(n8_adj_3824));   // verilog/motorControl.v(43[17:23])
    defparam i2_3_lut_4_lut_adj_1396.LUT_INIT = 16'hb748;
    SB_LUT4 i21926_3_lut_4_lut (.I0(n16635[1]), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n4_adj_4020), .O(n6_adj_4021));   // verilog/motorControl.v(43[17:23])
    defparam i21926_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[23]));   // verilog/motorControl.v(40[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i6_1_lut (.I0(\PID_CONTROLLER.err[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n63[5]));   // verilog/motorControl.v(43[31:45])
    defparam sub_11_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21918_4_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n16635[0]), .I3(n35561), .O(n4_adj_4020));   // verilog/motorControl.v(43[17:23])
    defparam i21918_4_lut_4_lut.LUT_INIT = 16'hf8a0;
    SB_LUT4 i21906_2_lut_3_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[1] ), .I3(GND_net), .O(n35561));   // verilog/motorControl.v(43[17:23])
    defparam i21906_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_1397 (.I0(n16635[2]), .I1(\Kp[4] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n6_adj_4021), .O(n16635[3]));   // verilog/motorControl.v(43[17:23])
    defparam i1_3_lut_4_lut_adj_1397.LUT_INIT = 16'h956a;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1398 (.I0(\Kd[3] ), .I1(n69[25]), .I2(n4_adj_3545), 
            .I3(n10844[1]), .O(n10844[2]));   // verilog/motorControl.v(43[26:45])
    defparam i1_2_lut_3_lut_4_lut_adj_1398.LUT_INIT = 16'h8778;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i18_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [10]), 
            .I1(\PID_CONTROLLER.result [11]), .I2(deadband[11]), .I3(GND_net), 
            .O(n18));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i18_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [2]), 
            .I1(\PID_CONTROLLER.result [3]), .I2(deadband[3]), .I3(GND_net), 
            .O(n6));   // verilog/motorControl.v(44[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n24202, encoder1_position, clk32MHz, 
            n24201, n24200, n24199, n24198, n24197, n24196, n24195, 
            n24194, n24193, n24192, n24191, n24190, n24189, n24188, 
            n24187, n24186, n24185, n24184, n24183, n24182, n24181, 
            n24170, data_o, n2226, GND_net, n23577, count_enable, 
            n24231, reg_B, n43884, PIN_18_c_1, PIN_19_c_0, n23580) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n24202;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n24201;
    input n24200;
    input n24199;
    input n24198;
    input n24197;
    input n24196;
    input n24195;
    input n24194;
    input n24193;
    input n24192;
    input n24191;
    input n24190;
    input n24189;
    input n24188;
    input n24187;
    input n24186;
    input n24185;
    input n24184;
    input n24183;
    input n24182;
    input n24181;
    input n24170;
    output [1:0]data_o;
    output [23:0]n2226;
    input GND_net;
    input n23577;
    output count_enable;
    input n24231;
    output [1:0]reg_B;
    output n43884;
    input PIN_18_c_1;
    input PIN_19_c_0;
    input n23580;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire B_delayed, A_delayed, n2216, n36081, n36080, n36079, n36078, 
        n36077, n36076, n36075, n36074, n36073, n36072, n36071, 
        n36070, n36069, n36068, n36067, n36066, n36065, n36064, 
        n36063, n36062, n36061, n36060, n36059, count_direction, 
        n36058;
    
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n24202));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n24201));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n24200));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n24199));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n24198));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n24197));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n24196));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n24195));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n24194));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n24193));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n24192));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n24191));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n24190));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n24189));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n24188));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n24187));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n24186));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n24185));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n24184));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n24183));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n24182));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n24181));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n24170));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_507_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2216), 
            .I3(n36081), .O(n2226[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_507_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2216), 
            .I3(n36080), .O(n2226[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_24 (.CI(n36080), .I0(encoder1_position[22]), .I1(n2216), 
            .CO(n36081));
    SB_LUT4 add_507_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2216), 
            .I3(n36079), .O(n2226[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_23 (.CI(n36079), .I0(encoder1_position[21]), .I1(n2216), 
            .CO(n36080));
    SB_LUT4 add_507_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2216), 
            .I3(n36078), .O(n2226[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_22 (.CI(n36078), .I0(encoder1_position[20]), .I1(n2216), 
            .CO(n36079));
    SB_LUT4 add_507_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2216), 
            .I3(n36077), .O(n2226[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_21 (.CI(n36077), .I0(encoder1_position[19]), .I1(n2216), 
            .CO(n36078));
    SB_LUT4 add_507_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2216), 
            .I3(n36076), .O(n2226[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_20 (.CI(n36076), .I0(encoder1_position[18]), .I1(n2216), 
            .CO(n36077));
    SB_LUT4 add_507_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2216), 
            .I3(n36075), .O(n2226[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_19 (.CI(n36075), .I0(encoder1_position[17]), .I1(n2216), 
            .CO(n36076));
    SB_LUT4 add_507_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2216), 
            .I3(n36074), .O(n2226[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_18 (.CI(n36074), .I0(encoder1_position[16]), .I1(n2216), 
            .CO(n36075));
    SB_LUT4 add_507_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2216), 
            .I3(n36073), .O(n2226[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_17 (.CI(n36073), .I0(encoder1_position[15]), .I1(n2216), 
            .CO(n36074));
    SB_LUT4 add_507_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2216), 
            .I3(n36072), .O(n2226[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_16 (.CI(n36072), .I0(encoder1_position[14]), .I1(n2216), 
            .CO(n36073));
    SB_LUT4 add_507_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2216), 
            .I3(n36071), .O(n2226[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_15 (.CI(n36071), .I0(encoder1_position[13]), .I1(n2216), 
            .CO(n36072));
    SB_LUT4 add_507_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2216), 
            .I3(n36070), .O(n2226[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_14 (.CI(n36070), .I0(encoder1_position[12]), .I1(n2216), 
            .CO(n36071));
    SB_LUT4 add_507_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2216), 
            .I3(n36069), .O(n2226[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_13 (.CI(n36069), .I0(encoder1_position[11]), .I1(n2216), 
            .CO(n36070));
    SB_LUT4 add_507_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2216), 
            .I3(n36068), .O(n2226[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_12 (.CI(n36068), .I0(encoder1_position[10]), .I1(n2216), 
            .CO(n36069));
    SB_LUT4 add_507_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2216), 
            .I3(n36067), .O(n2226[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_11 (.CI(n36067), .I0(encoder1_position[9]), .I1(n2216), 
            .CO(n36068));
    SB_LUT4 add_507_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2216), 
            .I3(n36066), .O(n2226[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_10 (.CI(n36066), .I0(encoder1_position[8]), .I1(n2216), 
            .CO(n36067));
    SB_LUT4 add_507_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2216), 
            .I3(n36065), .O(n2226[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_9 (.CI(n36065), .I0(encoder1_position[7]), .I1(n2216), 
            .CO(n36066));
    SB_LUT4 add_507_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2216), 
            .I3(n36064), .O(n2226[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_8 (.CI(n36064), .I0(encoder1_position[6]), .I1(n2216), 
            .CO(n36065));
    SB_LUT4 add_507_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2216), 
            .I3(n36063), .O(n2226[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_7 (.CI(n36063), .I0(encoder1_position[5]), .I1(n2216), 
            .CO(n36064));
    SB_LUT4 add_507_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2216), 
            .I3(n36062), .O(n2226[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_6 (.CI(n36062), .I0(encoder1_position[4]), .I1(n2216), 
            .CO(n36063));
    SB_LUT4 add_507_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2216), 
            .I3(n36061), .O(n2226[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_5 (.CI(n36061), .I0(encoder1_position[3]), .I1(n2216), 
            .CO(n36062));
    SB_LUT4 add_507_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2216), 
            .I3(n36060), .O(n2226[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_4 (.CI(n36060), .I0(encoder1_position[2]), .I1(n2216), 
            .CO(n36061));
    SB_LUT4 add_507_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2216), 
            .I3(n36059), .O(n2226[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_3 (.CI(n36059), .I0(encoder1_position[1]), .I1(n2216), 
            .CO(n36060));
    SB_LUT4 add_507_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n36058), .O(n2226[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_507_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_507_2 (.CI(n36058), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n36059));
    SB_CARRY add_507_1 (.CI(GND_net), .I0(n2216), .I1(n2216), .CO(n36058));
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n23577));   // quad.v(35[10] 41[6])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i773_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2216));   // quad.v(37[5] 40[8])
    defparam i773_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    \grp_debouncer(2,5)  debounce (.n24231(n24231), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .reg_B({reg_B}), .n43884(n43884), .GND_net(GND_net), .PIN_18_c_1(PIN_18_c_1), 
            .PIN_19_c_0(PIN_19_c_0), .n23580(n23580)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n24231, data_o, clk32MHz, reg_B, n43884, 
            GND_net, PIN_18_c_1, PIN_19_c_0, n23580) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24231;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    output n43884;
    input GND_net;
    input PIN_18_c_1;
    input PIN_19_c_0;
    input n23580;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    wire cnt_next_2__N_3113, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24231));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n43884));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFFSR cnt_reg_1017__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_18_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_19_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23580));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1017__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1017__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22289_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22289_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22282_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22282_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n43884), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22280_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22280_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=47, LSE_LCOL=12, LSE_RCOL=39, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, gearBoxRatio, GND_net, n24099, \data_in[0] , 
            n24098, n24097, n24096, n24095, n24094, n24093, n24092, 
            \data_in[1] , n24091, n24090, n24089, n24088, n24087, 
            n24086, n24085, n24084, \data_in[2] , n24083, n24082, 
            n24081, n24080, n24079, n24078, n24077, deadband, n24258, 
            setpoint, n24257, n24256, n24255, n24254, n24253, n24252, 
            n24251, n24250, n24249, n24248, n24247, n24246, n24245, 
            n24244, n24243, n24242, n24241, n24240, n24239, n24238, 
            n24237, n24236, VCC_net, IntegralLimit, n24063, \data_out_frame[5][2] , 
            rx_data, n24076, \data_in[3] , n24075, n24074, n24073, 
            rx_data_ready, n24072, \Kd[7] , n24071, n23930, \data_in_frame[1] , 
            n23929, n23928, n23927, n23926, n23925, n23924, n23923, 
            n23914, \data_in_frame[3] , n23913, n23912, n23911, n23910, 
            n23909, n23908, n23907, \FRAME_MATCHER.state , \FRAME_MATCHER.state[2] , 
            n23898, \data_in_frame[5] , n23897, n23896, n23895, n23894, 
            n23893, n23892, n23891, \Kp[1] , \data_in_frame[6][1] , 
            n23882, \data_in_frame[7] , n23881, n23880, n23879, n23878, 
            n23877, n23876, n23875, \data_in_frame[8] , \data_in_frame[8][2] , 
            \Kp[2] , n22501, n2, n42614, \Kp[3] , \Kp[4] , n5, 
            n23866, \data_in_frame[9] , n43935, \Kp[5] , n23865, n42406, 
            n23864, n23863, n23862, n23861, n23860, n23859, \data_in_frame[12][4] , 
            n23858, \data_in_frame[10] , n23857, n23856, n23855, n23854, 
            n23853, n23852, n23851, n23850, \data_in_frame[11] , n23849, 
            \Kp[6] , n20435, \data_in_frame[12][1] , \data_out_frame[0][4] , 
            n42421, n23848, n24070, \Kp[7] , n22289, \Ki[1] , \Ki[2] , 
            \Ki[3] , n23847, n22303, n23846, n28374, n23844, n23843, 
            n63, n20088, n23834, \data_in_frame[13] , n23833, n23832, 
            n23831, n23830, n26846, n23828, n23827, n23818, \data_in_frame[15] , 
            n124, n23817, n23816, n23815, n23814, n23813, n23812, 
            n23811, n2857, n89, n22424, n23802, \data_in_frame[17] , 
            n23801, n23800, n23799, n24069, n23798, n23797, n23796, 
            n23795, n23786, \data_in_frame[19] , n23785, n23784, n23783, 
            n23782, n23781, n23780, n23779, n23770, \data_in_frame[21] , 
            n23769, n23768, n23767, n23766, n23765, n23764, n23763, 
            control_mode, n20195, \Ki[4] , n42422, n20420, n43035, 
            PWMLimit, n49980, n49981, n43032, \Ki[5] , n43011, n24068, 
            \data_out_frame[0][2] , n24067, \data_out_frame[0][3] , n24066, 
            \Ki[6] , \Ki[7] , \Kd[1] , \Kd[2] , \Kd[3] , \Kd[4] , 
            \Kd[5] , \Kd[6] , LED_c, n22277, encoder1_position, n38879, 
            n23013, n22538, n3346, encoder0_position, n22589, n23584, 
            n41786, n23570, \Kd[0] , \Ki[0] , \Kp[0] , n42896, n42559, 
            n42920, displacement, n42621, pwm, n20471, n42418, n3790, 
            n407, \PID_CONTROLLER.result[13] , n27, n3791, n3792, 
            n3793, n3794, n5017, n3795, n3796, n3797, n3798, n3799, 
            r_SM_Main, n3800, n27_adj_3, n3801, n27_adj_4, n3802, 
            n3803, \pwm_23__N_2960[13] , n50261, n23444, n3804, n3805, 
            n3806, n123, n740, n16810, \FRAME_MATCHER.state_31__N_1989[1] , 
            n3807, n3808, n3809, n3810, n3811, n3812, n3813, n22296, 
            n22422, n3761, n2103, n22309, \FRAME_MATCHER.state_31__N_1861[2] , 
            n7, n22908, n42400, n42424, n42405, n42413, n23609, 
            \r_Clock_Count[8] , n23612, \r_Clock_Count[7] , n23615, 
            \r_Clock_Count[6] , n23618, \r_Clock_Count[5] , n23621, 
            \r_Clock_Count[4] , n23624, \r_Clock_Count[3] , n23627, 
            \r_Clock_Count[2] , n23630, \r_Clock_Count[1] , n23634, 
            r_Bit_Index, n23637, n24235, n23680, n313, n314, n315, 
            n316, n317, n318, \r_SM_Main_2__N_2753[1] , n319, n320, 
            n23629, n23463, n23547, n4032, o_Tx_Serial_N_2784, n49982, 
            n23583, n23581, tx_o, n49, tx_enable, n23640, r_Bit_Index_adj_12, 
            n23643, n28961, \r_SM_Main[1]_adj_8 , n23683, n24171, 
            r_Rx_Data, PIN_13_N_26, n46671, n46670, \r_SM_Main[2]_adj_9 , 
            n23457, n23545, n4010, n23650, n23649, n23648, n23647, 
            n23646, n23645, n23644, n23579, n22411, n4, n28925, 
            n1, n28462, n4_adj_10, n4_adj_11, n22416) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    output [23:0]gearBoxRatio;
    input GND_net;
    input n24099;
    output [7:0]\data_in[0] ;
    input n24098;
    input n24097;
    input n24096;
    input n24095;
    input n24094;
    input n24093;
    input n24092;
    output [7:0]\data_in[1] ;
    input n24091;
    input n24090;
    input n24089;
    input n24088;
    input n24087;
    input n24086;
    input n24085;
    input n24084;
    output [7:0]\data_in[2] ;
    input n24083;
    input n24082;
    input n24081;
    input n24080;
    input n24079;
    input n24078;
    input n24077;
    output [23:0]deadband;
    input n24258;
    output [23:0]setpoint;
    input n24257;
    input n24256;
    input n24255;
    input n24254;
    input n24253;
    input n24252;
    input n24251;
    input n24250;
    input n24249;
    input n24248;
    input n24247;
    input n24246;
    input n24245;
    input n24244;
    input n24243;
    input n24242;
    input n24241;
    input n24240;
    input n24239;
    input n24238;
    input n24237;
    input n24236;
    input VCC_net;
    output [23:0]IntegralLimit;
    input n24063;
    output \data_out_frame[5][2] ;
    output [7:0]rx_data;
    input n24076;
    output [7:0]\data_in[3] ;
    input n24075;
    input n24074;
    input n24073;
    output rx_data_ready;
    input n24072;
    output \Kd[7] ;
    input n24071;
    input n23930;
    output [7:0]\data_in_frame[1] ;
    input n23929;
    input n23928;
    input n23927;
    input n23926;
    input n23925;
    input n23924;
    input n23923;
    input n23914;
    output [7:0]\data_in_frame[3] ;
    input n23913;
    input n23912;
    input n23911;
    input n23910;
    input n23909;
    input n23908;
    input n23907;
    output [31:0]\FRAME_MATCHER.state ;
    output \FRAME_MATCHER.state[2] ;
    input n23898;
    output [7:0]\data_in_frame[5] ;
    input n23897;
    input n23896;
    input n23895;
    input n23894;
    input n23893;
    input n23892;
    input n23891;
    output \Kp[1] ;
    output \data_in_frame[6][1] ;
    input n23882;
    output [7:0]\data_in_frame[7] ;
    input n23881;
    input n23880;
    input n23879;
    input n23878;
    input n23877;
    input n23876;
    input n23875;
    output [7:0]\data_in_frame[8] ;
    output \data_in_frame[8][2] ;
    output \Kp[2] ;
    output n22501;
    output n2;
    output n42614;
    output \Kp[3] ;
    output \Kp[4] ;
    output n5;
    input n23866;
    output [7:0]\data_in_frame[9] ;
    output n43935;
    output \Kp[5] ;
    input n23865;
    output n42406;
    input n23864;
    input n23863;
    input n23862;
    input n23861;
    input n23860;
    input n23859;
    output \data_in_frame[12][4] ;
    input n23858;
    output [7:0]\data_in_frame[10] ;
    input n23857;
    input n23856;
    input n23855;
    input n23854;
    input n23853;
    input n23852;
    input n23851;
    input n23850;
    output [7:0]\data_in_frame[11] ;
    input n23849;
    output \Kp[6] ;
    output n20435;
    output \data_in_frame[12][1] ;
    output \data_out_frame[0][4] ;
    output n42421;
    input n23848;
    input n24070;
    output \Kp[7] ;
    output n22289;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    input n23847;
    output n22303;
    input n23846;
    input n28374;
    input n23844;
    input n23843;
    output n63;
    output n20088;
    input n23834;
    output [7:0]\data_in_frame[13] ;
    input n23833;
    input n23832;
    input n23831;
    input n23830;
    input n26846;
    input n23828;
    input n23827;
    input n23818;
    output [7:0]\data_in_frame[15] ;
    output n124;
    input n23817;
    input n23816;
    input n23815;
    input n23814;
    input n23813;
    input n23812;
    input n23811;
    output n2857;
    output n89;
    output n22424;
    input n23802;
    output [7:0]\data_in_frame[17] ;
    input n23801;
    input n23800;
    input n23799;
    input n24069;
    input n23798;
    input n23797;
    input n23796;
    input n23795;
    input n23786;
    output [7:0]\data_in_frame[19] ;
    input n23785;
    input n23784;
    input n23783;
    input n23782;
    input n23781;
    input n23780;
    input n23779;
    input n23770;
    output [7:0]\data_in_frame[21] ;
    input n23769;
    input n23768;
    input n23767;
    input n23766;
    input n23765;
    input n23764;
    input n23763;
    output [7:0]control_mode;
    output n20195;
    output \Ki[4] ;
    output n42422;
    output n20420;
    input n43035;
    output [23:0]PWMLimit;
    input n49980;
    input n49981;
    input n43032;
    output \Ki[5] ;
    input n43011;
    input n24068;
    output \data_out_frame[0][2] ;
    input n24067;
    output \data_out_frame[0][3] ;
    input n24066;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Kd[1] ;
    output \Kd[2] ;
    output \Kd[3] ;
    output \Kd[4] ;
    output \Kd[5] ;
    output \Kd[6] ;
    output LED_c;
    output n22277;
    input [23:0]encoder1_position;
    input n38879;
    output n23013;
    output n22538;
    output n3346;
    input [23:0]encoder0_position;
    input n22589;
    input n23584;
    input n41786;
    input n23570;
    output \Kd[0] ;
    output \Ki[0] ;
    output \Kp[0] ;
    input n42896;
    input n42559;
    output n42920;
    input [23:0]displacement;
    input n42621;
    input [23:0]pwm;
    output n20471;
    output n42418;
    output n3790;
    input n407;
    input \PID_CONTROLLER.result[13] ;
    output n27;
    output n3791;
    output n3792;
    output n3793;
    output n3794;
    output n5017;
    output n3795;
    output n3796;
    output n3797;
    output n3798;
    output n3799;
    output [2:0]r_SM_Main;
    output n3800;
    output n27_adj_3;
    output n3801;
    output n27_adj_4;
    output n3802;
    output n3803;
    input \pwm_23__N_2960[13] ;
    output n50261;
    output n23444;
    output n3804;
    output n3805;
    output n3806;
    output n123;
    output n740;
    output n16810;
    output \FRAME_MATCHER.state_31__N_1989[1] ;
    output n3807;
    output n3808;
    output n3809;
    output n3810;
    output n3811;
    output n3812;
    output n3813;
    output n22296;
    output n22422;
    output n3761;
    output n2103;
    output n22309;
    output \FRAME_MATCHER.state_31__N_1861[2] ;
    output n7;
    output n22908;
    output n42400;
    output n42424;
    output n42405;
    output n42413;
    input n23609;
    output \r_Clock_Count[8] ;
    input n23612;
    output \r_Clock_Count[7] ;
    input n23615;
    output \r_Clock_Count[6] ;
    input n23618;
    output \r_Clock_Count[5] ;
    input n23621;
    output \r_Clock_Count[4] ;
    input n23624;
    output \r_Clock_Count[3] ;
    input n23627;
    output \r_Clock_Count[2] ;
    input n23630;
    output \r_Clock_Count[1] ;
    input n23634;
    output [2:0]r_Bit_Index;
    input n23637;
    input n24235;
    input n23680;
    output n313;
    output n314;
    output n315;
    output n316;
    output n317;
    output n318;
    output \r_SM_Main_2__N_2753[1] ;
    output n319;
    output n320;
    output n23629;
    output n23463;
    output n23547;
    output n4032;
    output o_Tx_Serial_N_2784;
    input n49982;
    input n23583;
    input n23581;
    output tx_o;
    output n49;
    output tx_enable;
    input n23640;
    output [2:0]r_Bit_Index_adj_12;
    input n23643;
    input n28961;
    output \r_SM_Main[1]_adj_8 ;
    input n23683;
    input n24171;
    output r_Rx_Data;
    input PIN_13_N_26;
    output n46671;
    output n46670;
    output \r_SM_Main[2]_adj_9 ;
    output n23457;
    output n23545;
    output n4010;
    input n23650;
    input n23649;
    input n23648;
    input n23647;
    input n23646;
    input n23645;
    input n23644;
    input n23579;
    output n22411;
    output n4;
    output n28925;
    output n1;
    output n28462;
    output n4_adj_10;
    output n4_adj_11;
    output n22416;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n24028;
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    
    wire n24027, n24026, n24025;
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    
    wire n24024, n24023, n24022, n24103, n24102, n24101, n24100, 
        n24021, n35873;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n35874, n35861, n35862, n24020, n24019, n24018, n2_c, 
        n35872, n1498, n24017;
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    
    wire n24016, n24015, n24014, n24013, n24012, n24011, n24010, 
        n24009;
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    
    wire n24008, n24282, n24281, n24280, n24279, n24278, n24277, 
        n24276, n24275, n24274, n24273, n24272, n24271, n24270, 
        n24269, n24268, n24267, n24266, n24265, n24264, n24263, 
        n24262, n24261, n24259, n24234;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire n23653, n23656, n23659, n23662, n23665, n23668, n24177, 
        n24169, n24168, n24167, n24166, n24165, n24164, n24163, 
        n24162, n24161, n24160, n24159, n24158, n24157, n24156, 
        n24155, n24007, n24064;
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    
    wire n24006, n24005, n24062, n24004, n24061, n24003, n24060, 
        n24002, n24059, n24001;
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    
    wire n24058, n24000, n24057;
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    
    wire n23999, n24056, n23998, n24055, n23997, n24054, n23996, 
        n24053, n23995, n24052, n23994, n24051, n23993;
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    
    wire n24050, n24049;
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    
    wire n24048, n24047, n24046, n24045, n24044, n24043, n24042, 
        n24041;
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    
    wire n24040, n24118, n24117, n24116, n24115, n24114, n24113, 
        n24112, n24039, n24038, n24037, n24036, n24035, n24034, 
        n23992, n23991, n24033, n24032, n23990, n24111, n23989, 
        n23988, n10, n42399;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    
    wire n23915, n23987, n23916, n23986, n23985;
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    
    wire n23984, n23983, n23982, n23981, n23980, n23979, n23978, 
        n23977;
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    
    wire n23976, n23975, n23974, n23973, n23972, n23971, n23970, 
        n23969;
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    
    wire n23968, \FRAME_MATCHER.rx_data_ready_prev , n23967, n23966, 
        n23965, n23964, n23963, n23962, n23961;
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    
    wire n24123, n24122, n24110, n24151, n23960, n23959, n23958, 
        n23957, n23956, n23955, n24150, n24149, n23954, n24148, 
        n24147, n23953;
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    
    wire n23952, n23951, n23950, n23949, n23948, n23947, n23946, 
        n23945;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    
    wire n23944, n23943, n23942, n23941, n23940, n23939, n23938, 
        n23937;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire n23936, n23935, n23934, n23917, n23933, n23932, n23931, 
        n23922, n23921, n23920, n23919, n23918, n24146, n23906;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    
    wire n23905, n23904, n23903;
    wire [31:0]\FRAME_MATCHER.state_c ;   // verilog/coms.v(110[11:16])
    
    wire n45, n23902, n23901, n23900, n23899, n43207, n28433, 
        n6, n28987, n28413, n22274, n3831, n23890;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    
    wire n24145, n24144, n24143, n2_adj_3117, n35860, n23889, n23888, 
        n23887, n23886, n23885, n2_adj_3118, n35871, n23884, n23883, 
        n24031, n24030, n23874, n23873;
    wire [7:0]\data_in_frame[8]_c ;   // verilog/coms.v(94[12:25])
    
    wire n23872, n23871, n23870, n23869, n23868, n23867, n24142, 
        n28411, Kp_23__N_152, n31, n43149, n22777, n15, n8, n22554, 
        n16, n24141, n24140, n23042, n22941, n1_c, n8_adj_3120, 
        n19, n22657, n22, n13, n18, n38403, n19790, n24139, 
        n30654, n35924, n8_adj_3121, n42411;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    
    wire n23835, n23836, n23837, n19_adj_3122, n35923, n42403, n23838, 
        n23839, n23840, n23663, n35922, n24138, n23841, n23660, 
        n35921, n23842, n23657, n35920, n49962, n49965, n2_adj_3123, 
        n35859, n42419, n23654, n35919, n8_adj_3124;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    
    wire n23819, n23820, n23651, n35918, n23821, n23822, n23823, 
        n23824, n23825, n2_adj_3125, n35870, n23826, n8_adj_3126;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n23803, n23804;
    wire [7:0]n2236;
    
    wire tx_transmit_N_2648, n23805, n23806, n23807, n23808, n23809, 
        n28404, n23810, n22342, n22175, n10_adj_3127;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    
    wire n23787, n23788, n23789, n23790, n23791, n23792, n23793, 
        n23794, n61, n1_adj_3128, n37, n28837, n2_adj_3129, n35869, 
        n28839, n24137, n28841, n28843, n28845, n19_adj_3130, n46706, 
        n49968, n8_adj_3131, n8_adj_3132, n8_adj_3133, n41708, n22421, 
        n41714, n8_adj_3134, n24136, n24135, n24134, n2_adj_3135, 
        n35868, n22294, n28564, n8_adj_3136, n2_adj_3137, n35858, 
        n8_adj_3138, n2_adj_3139, n35867, n8_adj_3140, n2_adj_3141, 
        n35857, n2_adj_3142, n35866, n63_c, n63_adj_3143, n17, n16_adj_3145, 
        n49971, n46688, n5_adj_3146, n49956, n49959, n49950, n49953, 
        n49944, n49947, n49938, n49941, n49932, n49935, n49926, 
        n49929, n49920, n49923, n49914, n49917, n49908, n49911, 
        n7_c, n42390, n2_adj_3147, n35865, n49902, n53, n32579, 
        n2_adj_3148, n35856, n49905, n42971, n21986, n7_adj_3149, 
        n2_adj_3150, n35886, n42430, n42770, n42846, n42377, n41780, 
        n42375, n41732, n7_adj_3151, n7_adj_3152, n7_adj_3153, n42376, 
        n41726, n42384, n41728, n7_adj_3154, n42388, n41782, n7_adj_3155, 
        n42380, n41784, n42378, n41730, n7_adj_3156, n7_adj_3157, 
        n42386, n41788, n7_adj_3158, n28432, n28430, n42383, n41790, 
        n42387, n41724, n42382, n42374, n28428, n42379, n41792, 
        n42381, n41794, n42389, n41796, n42385, n41722, n41720, 
        n41950, n43887, n23438;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    
    wire n22077, n38954, n10_adj_3159, n1506, n39131, n42549, n43836, 
        n42464, n43657, n43874, n43873, n42734, n42735, n44064;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n43976, n43972, n42492, n43853, n43560, n43845, n43454, 
        n23194, n10_adj_3160, n42480, n42646, n3, n42471, n42806, 
        n2_adj_3161, n35885, n2_adj_3162, n35864, n23004, n42803, 
        n23247, n42584, n43500, n43803, n3_adj_3163, n2_adj_3164, 
        n3_adj_3165, n2_adj_3166, n3_adj_3167, n2_adj_3168, n3_adj_3169, 
        n2_adj_3170, n3_adj_3171, n2_adj_3172, n3_adj_3173, n2_adj_3174, 
        n3_adj_3175, n2_adj_3176, n3_adj_3177, n2_adj_3178, n3_adj_3179, 
        n2_adj_3180, n3_adj_3181, n2_adj_3182, n3_adj_3183, n2_adj_3184, 
        n3_adj_3185, n2_adj_3186, n3_adj_3187, n3_adj_3188, n3_adj_3189, 
        n3_adj_3190, n3_adj_3191, n3_adj_3192, n3_adj_3193, n3_adj_3194, 
        n3_adj_3195, n3_adj_3196, n2_adj_3197, n3_adj_3198, n2_adj_3199, 
        n3_adj_3200, n2_adj_3201, n3_adj_3202, n3_adj_3203, n3_adj_3204, 
        n3_adj_3205, n3_adj_3206, n3_adj_3207, n10_adj_3208, n42688, 
        n39144, n42849, n35884, n24121, n24120, n24119, n49896, 
        n49899, n35883, n49890, n23778;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    
    wire n23777, n23776, n23775, n35882, n23774, n23773, n23772, 
        n23771, n35881, n23762, n35880, n24133, n49893, n23761, 
        n23760, n23064, n42717, n49884, n42926, n7_adj_3209, n10_adj_3210, 
        n38377, n23759, n23758, n23757, n23756, n23755, n23754, 
        n23753, n23752, n26838, n23750, n23749, n23748, n23747, 
        n23746, n23745, n23744, n27693, n27746, n23741, n23740, 
        n23739, n23738, n23737, n28334, n28366, n23734, n23733, 
        n35879, n22745, n42742, n10_adj_3211, n42941, n22611, n14, 
        n43038, n42843, n42793, n39163, n42910, n26, n23244, n24, 
        n49887, n49878, n49881, n49872, n49875, n49866, n49869, 
        n49860, n49863, n49854, n49857, n22723, n38367, n25, n24132, 
        n23, n42796, n49848, n49851, n46769;
    wire [2:0]r_SM_Main_2__N_2756;
    
    wire n42202, n24109, n42536, n43029, n6_adj_3212, n43745, n42923, 
        n22993, n12, n35878, n24065, n24108, n35863, n24131, n38426, 
        n42678, n42545, n43056, n10_adj_3213, n39117, n49836, n42591, 
        n42953, n8_adj_3214, n42840, n42947, n39161, n24130, n24129, 
        n24128, n24127, n24126, n24125, n24124, n22299, n43084, 
        n8_adj_3215, n43008, n43069, n39133, n49839, n42879, n42998, 
        n42812, n43673, n42980, n43002, n20947, n12_adj_3216, Kp_23__N_176, 
        n22464, n42959, Kp_23__N_786, n42457, n44171, n28478, n48, 
        n46, n47, n42831, n42587, n45_adj_3217, n35877, n42799, 
        n42474, n44, n43, Kp_23__N_193, n54, n49_c, n35876, n49986, 
        n43005, n4_c, n43059, n42666, n38429, n24107, n22701, 
        n2_adj_3218, n164, n24106, n24105, n6_adj_3219, n24104, 
        n35875, n3_adj_3220, n23585, n24029, n23573, n23572, n23571, 
        n23569, n23568, n23567, n23566, n23565, n23105, n38473, 
        n23229, n42530, n42834, n12_adj_3221, n42983, n23178, n42494, 
        n22960, Kp_23__N_866, n23007, n22698, n42505, n42889, n39, 
        n42886, n51, n56, n42855, n42675, n42681, n42608, n54_adj_3222, 
        n22954, n55, n42861, n53_adj_3223, n50, n58, n62, n42858, 
        n49_adj_3224, n6_adj_3225, n43044, n42466, n42956, n28, 
        n32, n42819, n30, n42867, n31_adj_3226, n42524, n29, n39122, 
        n42995, n10_adj_3227, n42864, n42747, n42522, n42575, n12_adj_3228, 
        Kp_23__N_459, n42508, n22594, n42784, n6_adj_3229, Kp_23__N_379, 
        n42974, n6_adj_3230, n42736, n42611, n42567, n23049, n23309, 
        n6_adj_3231, n12_adj_3232, n23324, n12_adj_3233, n12_adj_3234, 
        n42516, n42708, n42572, n42892, n44074, n12_adj_3235, n42562, 
        n8_adj_3236, n23238, n20914, n42852, n42443, n4_adj_3237, 
        n22824, n5_adj_3238, n42870, Kp_23__N_326, n42899, n18_adj_3239, 
        n30_adj_3240, n42787, n22629, n28_adj_3241, n29_adj_3242, 
        n27_c, n22837, n42815, n10_adj_3243, n19_adj_3244, n46920, 
        n5_adj_3245, n44416, n44417, n44388, n44390, n42663, n44389, 
        n42649, n42630, n12_adj_3246, n38982, n12_adj_3247, n42828, 
        n22560, n14_adj_3248, n14_adj_3249, n13_adj_3250, n13_adj_3251, 
        n10_adj_3252, n43318, n10_adj_3253, n42686, n12_adj_3254, 
        n43047, n8_adj_3255, n42950, n43516, n12_adj_3256, n43674, 
        n43338, n42460, n44317, n42753, n10_adj_3257, n43536, n6_adj_3258, 
        n43313, n44313, n22_adj_3259, n44315, n21, n14_adj_3260, 
        n15_adj_3261, n43672, n18_adj_3262, n26_adj_3263, n30_adj_3264, 
        n17_adj_3265, n63_adj_3266, n49830, n49833, n49824, n23411, 
        tx_active, n23582, n19_adj_3269, n47082, n5_adj_3270, n44386, 
        n44387, n45253, n44412, n44414, n44413, n19_adj_3271, n47075, 
        n5_adj_3272, n44383, n44384, n44409, n44411, n44410, n19_adj_3274, 
        n47070, n5_adj_3275, n44380, n49827, n44381, n44406, n44408, 
        n44407, n19_adj_3276, n44377, n48799, n49821, n44378, n48803;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    wire n46666, n6_adj_3277, n5_adj_3278, n44397, n44399, n44398, 
        n46663, n19_adj_3279, n6_adj_3280, n5_adj_3281, n44422, n44423, 
        n44394, n44396, n44395, n19_adj_3282, n47051, n5_adj_3283, 
        n44419, n44420, n44391, n44393, n44392, n28971, n28985, 
        n4_adj_3284, n5019;
    wire [31:0]\FRAME_MATCHER.state_31__N_1925 ;
    
    wire n44365, n38, n39_adj_3285, n37_adj_3286, n44361, n46_adj_3287, 
        n44363, n42691, n6_adj_3288, n38418, n42902, n38867, n38351, 
        n12_adj_3289, n43017, n23136, n1716, n42758, n6_adj_3290, 
        n42491, n23295, n42550, n22668, n10_adj_3291, n44169, n42731, 
        n23267, n1444, n1695, n12_adj_3292, n42477, n42723, n1509, 
        n42598, n1595, n38210, n6_adj_3293, n22520, n42917, n39149, 
        n12_adj_3294, n43026, n42595, n42533, n42932, n42944, n22779, 
        n12_adj_3295, n43041, n39125, n28_adj_3296, n43065, n42876, 
        n43020, n31_adj_3297, n38811, n42751, n23251, n30_adj_3298, 
        n34, n22674, n29_adj_3299, n23345, n42929, n22019, n42720, 
        n42764, n16_adj_3300, n42542, n42761, n42694, n17_adj_3301, 
        n21999, n14_adj_3302, n15_adj_3303, n23114, n38353, n22017, 
        n39189, n14_adj_3304, n43050, n42977, n15_adj_3305, n42704, 
        n22926, n42781, n42434, n22445, n12_adj_3306, n42809, n22458, 
        n1515, n42822, n10_adj_3307, n42992, n20, n42883, n19_adj_3308, 
        n21_adj_3309, n44021, n18_adj_3310, n42905, n20_adj_3311, 
        n15_adj_3312, n38601, n22793, n35, n6_adj_3313, n12_adj_3314, 
        n42938, n42669, n43023, n42450, n22937, n22482, n22843, 
        n18_adj_3315, n16_adj_3316, n20_adj_3317, n42935, n42453, 
        n42672, n38668, n23274, n42711, n10_adj_3318, n42659, n42642, 
        n42700, n22853, n23111, n6_adj_3319, n18_adj_3320, n30_adj_3321, 
        n42498, n42986, n28_adj_3322, n42539, n29_adj_3323, n43053, 
        n27_adj_3324, n20_adj_3325, n19_adj_3326, n21_adj_3327, n42913, 
        n42641, n42965, n10_adj_3328, n42463, n39102, n42655, n38948, 
        n23271, n42837, n42989, n10_adj_3329, n7_adj_3330, n42501, 
        n42774, n14_adj_3331, n10_adj_3332, n42968, n6_adj_3333, n42778, 
        n42825, n42605, n12_adj_3334, n12_adj_3335, n18_adj_3336, 
        n16_adj_3337, n20_adj_3338, n6_adj_3339, n3_adj_3340, n11, 
        n22297, n12_adj_3341, n42373, n7_adj_3342, n42371, n20078, 
        n30621, n5_adj_3343, n8_adj_3344, n14_adj_3345, n13_adj_3346, 
        n20_adj_3347, n19_adj_3348, n32_adj_3349, n30_adj_3350, n31_adj_3351, 
        n29_adj_3352, n14_adj_3353, n22408, n15_adj_3354, n22195, 
        n16_adj_3355, n17_adj_3356, n22280, n10_adj_3357, n14_adj_3358, 
        n9, n22316, n18_adj_3359, n20_adj_3360, n15_adj_3361, n16_adj_3362, 
        n17_adj_3363, n20_adj_3364, n19_adj_3365, n44367, n4_adj_3366, 
        n43205, n49818;
    
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n24028));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n24027));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n24026));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n24025));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n24024));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n24023));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n24022));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n24103));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n24102));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n24101));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n24100));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n24021));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_20 (.CI(n35873), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n35874));
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n24099));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_8 (.CI(n35861), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n35862));
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n24098));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n24097));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n24020));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n24019));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n24018));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_19_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n35872), .O(n2_c)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n24017));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n24096));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n24016));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n24015));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n24014));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n24013));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n24012));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n24011));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n24010));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n24009));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n24095));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n24094));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n24093));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n24092));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n24091));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n24090));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n24089));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n24088));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n24087));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n24086));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n24085));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n24084));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n24083));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n24082));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n24081));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n24080));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n24079));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n24078));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n24077));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n24008));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i23 (.Q(deadband[23]), .C(clk32MHz), .D(n24282));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i22 (.Q(deadband[22]), .C(clk32MHz), .D(n24281));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i21 (.Q(deadband[21]), .C(clk32MHz), .D(n24280));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i20 (.Q(deadband[20]), .C(clk32MHz), .D(n24279));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i19 (.Q(deadband[19]), .C(clk32MHz), .D(n24278));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i18 (.Q(deadband[18]), .C(clk32MHz), .D(n24277));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i17 (.Q(deadband[17]), .C(clk32MHz), .D(n24276));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i16 (.Q(deadband[16]), .C(clk32MHz), .D(n24275));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i15 (.Q(deadband[15]), .C(clk32MHz), .D(n24274));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i14 (.Q(deadband[14]), .C(clk32MHz), .D(n24273));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i13 (.Q(deadband[13]), .C(clk32MHz), .D(n24272));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i12 (.Q(deadband[12]), .C(clk32MHz), .D(n24271));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i11 (.Q(deadband[11]), .C(clk32MHz), .D(n24270));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i10 (.Q(deadband[10]), .C(clk32MHz), .D(n24269));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i9 (.Q(deadband[9]), .C(clk32MHz), .D(n24268));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i8 (.Q(deadband[8]), .C(clk32MHz), .D(n24267));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i7 (.Q(deadband[7]), .C(clk32MHz), .D(n24266));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i6 (.Q(deadband[6]), .C(clk32MHz), .D(n24265));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i5 (.Q(deadband[5]), .C(clk32MHz), .D(n24264));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i4 (.Q(deadband[4]), .C(clk32MHz), .D(n24263));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i3 (.Q(deadband[3]), .C(clk32MHz), .D(n24262));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i2 (.Q(deadband[2]), .C(clk32MHz), .D(n24261));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i1 (.Q(deadband[1]), .C(clk32MHz), .D(n24259));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n24258));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n24257));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n24256));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n24255));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n24254));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n24253));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n24252));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n24251));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n24250));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n24249));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n24248));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n24247));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n24246));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n24245));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n24244));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n24243));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n24242));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n24241));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n24240));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n24239));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n24238));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n24237));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n24236));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(VCC_net), .D(n24234));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
           .D(n23653));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
           .D(n23656));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
           .D(n23659));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
           .D(n23662));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
           .D(n23665));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
           .D(n23668));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
           .D(n24177));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n24169));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n24168));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n24167));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n24166));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n24165));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n24164));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n24163));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n24162));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n24161));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n24160));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n24159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n24158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n24157));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n24156));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n24155));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n24007));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n24064));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n24006));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5][2] ), .C(clk32MHz), 
           .D(n24063));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n24005));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n24062));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n24004));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n24061));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n24003));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n24060));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n24002));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n24059));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n24001));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n24058));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n24000));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n24057));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n23999));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n24056));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n23998));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n24055));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n23997));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n24054));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n23996));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n24053));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n23995));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n24052));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n23994));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n24051));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n23993));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n24050));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n24049));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n24048));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n24047));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n24046));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n24045));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n24044));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n24043));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n24042));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n24041));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n24040));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n24118));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n24117));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n24116));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n24115));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n24114));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n24113));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n24112));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n24039));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n24038));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n24037));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n24036));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n24035));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n24034));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n23992));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n23991));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n24033));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n24032));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n23990));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n24111));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n23989));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n23988));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10501_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n23915));
    defparam i10501_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n24076));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n23987));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10502_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n23916));
    defparam i10502_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n23986));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n23985));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n23984));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n23983));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n23982));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n24075));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n23981));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n23980));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n23979));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n23978));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n23977));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n23976));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n23975));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n24074));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n24073));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n23974));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n23973));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n23972));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n23971));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n23970));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n23969));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n23968));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3228  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n23967));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n23966));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n23965));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n23964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n23963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n23962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n24072));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n23961));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i7 (.Q(\Kd[7] ), .C(clk32MHz), .D(n24123));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n24122));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n24110));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n24071));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n24151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n23960));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n23959));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n23958));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n23957));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n23956));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n23955));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n24150));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n24149));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n23954));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n24148));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n24147));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n23953));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n23952));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n23951));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n23950));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n23949));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n23948));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n23947));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n23946));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n23945));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n23944));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n23943));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n23942));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n23941));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n23940));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n23939));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n23938));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n23937));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n23936));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n23935));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n23934));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10503_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n23917));
    defparam i10503_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n23933));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n23932));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n23931));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n23930));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n23929));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n23928));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n23927));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n23926));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n23925));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n23924));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n23923));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n23922));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n23921));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n23920));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n23919));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n23918));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n23917));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n23916));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n23915));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n23914));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n23913));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n23912));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n23911));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n24146));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n23910));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n23909));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n23908));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n23907));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n23906));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n23905));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n23904));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n23903));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/coms.v(110[11:16])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n23902));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n23901));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n23900));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n23899));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut (.I0(n43207), .I1(n28433), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(\FRAME_MATCHER.state[2] ), .O(n6));
    defparam i2_4_lut.LUT_INIT = 16'h5d55;
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n23898));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n23897));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut (.I0(n28987), .I1(n6), .I2(n28413), .I3(n22274), 
            .O(n3831));
    defparam i3_4_lut.LUT_INIT = 16'hfeee;
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n23896));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10504_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n23918));
    defparam i10504_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10505_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n23919));
    defparam i10505_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n23895));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n23894));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n23893));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n23892));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n23891));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n23890));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n24145));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_19 (.CI(n35872), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n35873));
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n24144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n24143));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_7_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n35860), .O(n2_adj_3117)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6][1] ), .C(clk32MHz), 
           .D(n23889));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n23888));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n23887));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n23886));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n23885));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_18_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n35871), .O(n2_adj_3118)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n23884));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n23883));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n23882));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n23881));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n24031));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10506_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n23920));
    defparam i10506_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n24030));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n23880));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n23879));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n23878));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n23877));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n23876));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n23875));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n23874));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8]_c [1]), .C(clk32MHz), 
           .D(n23873));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8][2] ), .C(clk32MHz), 
           .D(n23872));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8]_c [3]), .C(clk32MHz), 
           .D(n23871));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8]_c [4]), .C(clk32MHz), 
           .D(n23870));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8]_c [5]), .C(clk32MHz), 
           .D(n23869));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8]_c [6]), .C(clk32MHz), 
           .D(n23868));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8]_c [7]), .C(clk32MHz), 
           .D(n23867));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10507_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n23921));
    defparam i10507_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n24142));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i27592_4_lut (.I0(n28411), .I1(Kp_23__N_152), .I2(n31), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n43149));
    defparam i27592_4_lut.LUT_INIT = 16'hfabb;
    SB_LUT4 i3_3_lut (.I0(n22501), .I1(n22777), .I2(n15), .I3(GND_net), 
            .O(n8));   // verilog/coms.v(230[9:81])
    defparam i3_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i4_4_lut (.I0(n2), .I1(n22554), .I2(n8), .I3(n42614), .O(n16));   // verilog/coms.v(230[9:81])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n24141));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n24140));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i7_4_lut (.I0(n23042), .I1(n22941), .I2(n1_c), .I3(n8_adj_3120), 
            .O(n19));   // verilog/coms.v(230[9:81])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n19), .I1(n22657), .I2(n16), .I3(n5), .O(n22));   // verilog/coms.v(230[9:81])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n13), .I1(n22), .I2(n18), .I3(n38403), .O(n31));   // verilog/coms.v(230[9:81])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15022_2_lut (.I0(n31), .I1(n28411), .I2(GND_net), .I3(GND_net), 
            .O(n28413));
    defparam i15022_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n23866));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_3_lut_adj_828 (.I0(n43149), .I1(n19790), .I2(n28987), .I3(GND_net), 
            .O(n43935));
    defparam i3_3_lut_adj_828.LUT_INIT = 16'hfbfb;
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n24139));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_18 (.CI(n35871), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n35872));
    SB_LUT4 i10508_3_lut_4_lut (.I0(n10), .I1(n42399), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n23922));
    defparam i10508_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_547_9_lut (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[7]), 
            .I2(n3831), .I3(n35924), .O(n30654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_9_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i10421_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n23835));
    defparam i10421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10422_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n23836));
    defparam i10422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n23865));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10423_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n23837));
    defparam i10423_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_547_8_lut (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[6]), 
            .I2(n3831), .I3(n35923), .O(n19_adj_3122)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42403), .I3(\FRAME_MATCHER.i [0]), .O(n42406));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n23864));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n23863));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n23862));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n23861));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n23860));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n23859));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10424_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[4]), 
            .I3(\data_in_frame[12][4] ), .O(n23838));
    defparam i10424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10425_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n23839));
    defparam i10425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n23858));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n23857));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n23856));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_547_8 (.CI(n35923), .I0(byte_transmit_counter[6]), .I1(n3831), 
            .CO(n35924));
    SB_LUT4 i10426_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n23840));
    defparam i10426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n23855));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n23854));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_547_7_lut (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[5]), 
            .I2(n3831), .I3(n35922), .O(n23663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_7_lut.LUT_INIT = 16'hA3AC;
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n23853));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n23852));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n23851));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n23850));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n23849));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n24138));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_547_7 (.CI(n35922), .I0(byte_transmit_counter[5]), .I1(n3831), 
            .CO(n35923));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_829 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42411), .I3(\FRAME_MATCHER.i [0]), .O(n20435));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_829.LUT_INIT = 16'hfdff;
    SB_LUT4 i10427_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[1]), 
            .I3(\data_in_frame[12][1] ), .O(n23841));
    defparam i10427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_7 (.CI(n35860), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n35861));
    SB_LUT4 add_547_6_lut (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[4]), 
            .I2(n3831), .I3(n35921), .O(n23660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_547_6 (.CI(n35921), .I0(byte_transmit_counter[4]), .I1(n3831), 
            .CO(n35922));
    SB_LUT4 i10428_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42411), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n23842));
    defparam i10428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_547_5_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[3]), 
            .I2(n3831), .I3(n35920), .O(n23657)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 n49962_bdd_4_lut_4_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(n49962), .O(n49965));
    defparam n49962_bdd_4_lut_4_lut.LUT_INIT = 16'hfc02;
    SB_CARRY add_547_5 (.CI(n35920), .I0(byte_transmit_counter[3]), .I1(n3831), 
            .CO(n35921));
    SB_LUT4 add_44_6_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n35859), .O(n2_adj_3123)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_830 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42419), .I3(\FRAME_MATCHER.i [0]), .O(n42421));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_830.LUT_INIT = 16'hfdff;
    SB_LUT4 add_547_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[2]), 
            .I2(n3831), .I3(n35919), .O(n23654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i10405_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n23819));
    defparam i10405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10406_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n23820));
    defparam i10406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_547_4 (.CI(n35919), .I0(byte_transmit_counter[2]), .I1(n3831), 
            .CO(n35920));
    SB_LUT4 add_547_3_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[1]), 
            .I2(n3831), .I3(n35918), .O(n23651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i10407_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n23821));
    defparam i10407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10408_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n23822));
    defparam i10408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10409_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n23823));
    defparam i10409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10410_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n23824));
    defparam i10410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10411_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n23825));
    defparam i10411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_17_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n35870), .O(n2_adj_3125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10412_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42411), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n23826));
    defparam i10412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10389_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n23803));
    defparam i10389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10390_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n23804));
    defparam i10390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_547_3 (.CI(n35918), .I0(byte_transmit_counter[1]), .I1(n3831), 
            .CO(n35919));
    SB_LUT4 add_547_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_2648), .I3(GND_net), .O(n2236[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_547_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10391_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n23805));
    defparam i10391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n23848));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10392_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n23806));
    defparam i10392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10393_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n23807));
    defparam i10393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10394_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n23808));
    defparam i10394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10395_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n23809));
    defparam i10395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n28404), .O(n42399));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i10396_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42419), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n23810));
    defparam i10396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_831 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n22342), .I3(\FRAME_MATCHER.i [4]), .O(n22175));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_831.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(GND_net), .O(n10_adj_3127));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i10373_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n23787));
    defparam i10373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10374_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n23788));
    defparam i10374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10375_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n23789));
    defparam i10375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10376_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n23790));
    defparam i10376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n24070));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10377_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n23791));
    defparam i10377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10378_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n23792));
    defparam i10378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_17 (.CI(n35870), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n35871));
    SB_LUT4 i10379_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n23793));
    defparam i10379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10380_3_lut_4_lut (.I0(n10_adj_3127), .I1(n42399), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n23794));
    defparam i10380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_6 (.CI(n35859), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n35860));
    SB_LUT4 i15436_2_lut_4_lut (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [8]), .O(n28837));
    defparam i15436_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 add_44_16_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n35869), .O(n2_adj_3129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut (.I0(n61), .I1(n1_adj_3128), .I2(n37), .I3(\FRAME_MATCHER.state_c [9]), 
            .O(n28839));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n24137));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i15438_2_lut_4_lut (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [10]), .O(n28841));
    defparam i15438_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i15439_2_lut_4_lut (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [13]), .O(n28843));
    defparam i15439_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i15440_2_lut_4_lut (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [14]), .O(n28845));
    defparam i15440_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_3130), .I2(n46706), .I3(byte_transmit_counter[2]), 
            .O(n49968));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_832 (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [15]), .O(n8_adj_3131));
    defparam i1_2_lut_4_lut_adj_832.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_833 (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [17]), .O(n8_adj_3132));
    defparam i1_2_lut_4_lut_adj_833.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_834 (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [18]), .O(n8_adj_3133));
    defparam i1_2_lut_4_lut_adj_834.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_835 (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [21]), .O(n41708));
    defparam i1_2_lut_4_lut_adj_835.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_836 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n28987), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(GND_net), .O(n22289));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_3_lut_adj_836.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_837 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n28987), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(GND_net), .O(n22421));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_3_lut_adj_837.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_4_lut_adj_838 (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [23]), .O(n41714));
    defparam i1_2_lut_4_lut_adj_838.LUT_INIT = 16'hfe00;
    SB_CARRY add_547_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_2648), 
            .CO(n35918));
    SB_CARRY add_44_16 (.CI(n35869), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n35870));
    SB_LUT4 i1_2_lut_4_lut_adj_839 (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [26]), .O(n8_adj_3134));
    defparam i1_2_lut_4_lut_adj_839.LUT_INIT = 16'hfe00;
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n24136));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n24135));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n24134));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n23847));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_15_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n35868), .O(n2_adj_3135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_840 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n28987), 
            .I2(n22294), .I3(n22303), .O(n28564));   // verilog/coms.v(152[5:27])
    defparam i2_3_lut_4_lut_adj_840.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_841 (.I0(n61), .I1(n1_adj_3128), .I2(n37), 
            .I3(\FRAME_MATCHER.state_c [27]), .O(n8_adj_3136));
    defparam i1_2_lut_4_lut_adj_841.LUT_INIT = 16'hfe00;
    SB_LUT4 add_44_5_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n35858), .O(n2_adj_3137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_15 (.CI(n35868), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n35869));
    SB_LUT4 i78_2_lut_4_lut (.I0(n61), .I1(n1_adj_3128), .I2(n37), .I3(\FRAME_MATCHER.state_c [28]), 
            .O(n8_adj_3138));
    defparam i78_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 add_44_14_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n35867), .O(n2_adj_3139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_14 (.CI(n35867), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n35868));
    SB_LUT4 i68_2_lut_4_lut (.I0(n61), .I1(n1_adj_3128), .I2(n37), .I3(\FRAME_MATCHER.state_c [31]), 
            .O(n8_adj_3140));
    defparam i68_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_CARRY add_44_5 (.CI(n35858), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n35859));
    SB_LUT4 add_44_4_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n35857), .O(n2_adj_3141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n23846));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n28374));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n23844));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n23843));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_13_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n35866), .O(n2_adj_3142)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10485_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n23899));
    defparam i10485_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_842 (.I0(n63_c), .I1(n63_adj_3143), .I2(n63), 
            .I3(GND_net), .O(n20088));
    defparam i1_2_lut_3_lut_adj_842.LUT_INIT = 16'h8080;
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n23842));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49968_bdd_4_lut (.I0(n49968), .I1(n17), .I2(n16_adj_3145), 
            .I3(byte_transmit_counter[2]), .O(n49971));
    defparam n49968_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12][1] ), .C(clk32MHz), 
           .D(n23841));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n23840));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_34384 (.I0(byte_transmit_counter[1]), 
            .I1(n46688), .I2(n5_adj_3146), .I3(byte_transmit_counter[2]), 
            .O(n49962));
    defparam byte_transmit_counter_1__bdd_4_lut_34384.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n23839));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12][4] ), .C(clk32MHz), 
           .D(n23838));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n23837));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n49956));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n23836));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49956_bdd_4_lut (.I0(n49956), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n49959));
    defparam n49956_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n23835));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n23834));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34375 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n49950));
    defparam byte_transmit_counter_0__bdd_4_lut_34375.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n23833));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49950_bdd_4_lut (.I0(n49950), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n49953));
    defparam n49950_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n23832));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n23831));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34370 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n49944));
    defparam byte_transmit_counter_0__bdd_4_lut_34370.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n23830));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49944_bdd_4_lut (.I0(n49944), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n49947));
    defparam n49944_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n26846));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n23828));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34365 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n49938));
    defparam byte_transmit_counter_0__bdd_4_lut_34365.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n23827));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49938_bdd_4_lut (.I0(n49938), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n49941));
    defparam n49938_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n23826));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n23825));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34360 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n49932));
    defparam byte_transmit_counter_0__bdd_4_lut_34360.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n23824));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49932_bdd_4_lut (.I0(n49932), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n49935));
    defparam n49932_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n23823));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n23822));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34355 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n49926));
    defparam byte_transmit_counter_0__bdd_4_lut_34355.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n23821));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49926_bdd_4_lut (.I0(n49926), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n49929));
    defparam n49926_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n23820));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n23819));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34350 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n49920));
    defparam byte_transmit_counter_0__bdd_4_lut_34350.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n23818));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i15305_2_lut_3_lut (.I0(n63_c), .I1(n63_adj_3143), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n124));
    defparam i15305_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n49920_bdd_4_lut (.I0(n49920), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n49923));
    defparam n49920_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n23817));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n23816));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34345 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n49914));
    defparam byte_transmit_counter_0__bdd_4_lut_34345.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n23815));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49914_bdd_4_lut (.I0(n49914), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n49917));
    defparam n49914_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n23814));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n23813));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34340 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n49908));
    defparam byte_transmit_counter_0__bdd_4_lut_34340.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n23812));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49908_bdd_4_lut (.I0(n49908), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n49911));
    defparam n49908_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n23811));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_13 (.CI(n35866), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n35867));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_843 (.I0(n2857), .I1(n20088), .I2(\FRAME_MATCHER.state [0]), 
            .I3(\FRAME_MATCHER.state[2] ), .O(n7_c));   // verilog/coms.v(221[6] 223[9])
    defparam i1_2_lut_3_lut_4_lut_adj_843.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_3_lut_adj_844 (.I0(n2857), .I1(n20088), .I2(n22303), 
            .I3(GND_net), .O(n61));   // verilog/coms.v(221[6] 223[9])
    defparam i1_2_lut_3_lut_adj_844.LUT_INIT = 16'h0404;
    SB_LUT4 i10486_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n23900));
    defparam i10486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_845 (.I0(n89), .I1(n20088), .I2(\FRAME_MATCHER.state [0]), 
            .I3(\FRAME_MATCHER.state[2] ), .O(n42390));
    defparam i1_2_lut_3_lut_4_lut_adj_845.LUT_INIT = 16'h8000;
    SB_LUT4 i10487_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n23901));
    defparam i10487_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n23810));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10488_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n23902));
    defparam i10488_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_12_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n35865), .O(n2_adj_3147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10489_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n23903));
    defparam i10489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_4 (.CI(n35857), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n35858));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34335 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n49902));
    defparam byte_transmit_counter_0__bdd_4_lut_34335.LUT_INIT = 16'he4aa;
    SB_LUT4 i76_3_lut_4_lut (.I0(n89), .I1(n20088), .I2(n53), .I3(n22424), 
            .O(n32579));
    defparam i76_3_lut_4_lut.LUT_INIT = 16'hf0f8;
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n23809));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n23808));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n23807));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n23806));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_12 (.CI(n35865), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n35866));
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n23805));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_3_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n35856), .O(n2_adj_3148)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n23804));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n23803));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49902_bdd_4_lut (.I0(n49902), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n49905));
    defparam n49902_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n23802));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n23801));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n23800));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n23799));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n24069));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n23798));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n23797));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n23796));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n23795));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n23794));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_846 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n42971), .I3(GND_net), .O(n21986));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_846.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n23793));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n23792));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n23791));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(clk32MHz), 
            .D(n7_adj_3149), .S(n8_adj_3140));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10490_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n23904));
    defparam i10490_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_33_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n35886), .O(n2_adj_3150)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_847 (.I0(n42430), .I1(n42770), .I2(\data_out_frame[15] [6]), 
            .I3(\data_out_frame[15] [7]), .O(n42846));
    defparam i2_3_lut_4_lut_adj_847.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(clk32MHz), 
            .D(n42377), .S(n41780));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(clk32MHz), 
            .D(n42375), .S(n41732));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(clk32MHz), 
            .D(n7_adj_3151), .S(n8_adj_3138));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(clk32MHz), 
            .D(n7_adj_3152), .S(n8_adj_3136));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(clk32MHz), 
            .D(n7_adj_3153), .S(n8_adj_3134));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(clk32MHz), 
            .D(n42376), .S(n41726));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(clk32MHz), 
            .D(n42384), .S(n41728));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(clk32MHz), 
            .D(n7_adj_3154), .S(n41714));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(clk32MHz), 
            .D(n42388), .S(n41782));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(clk32MHz), 
            .D(n7_adj_3155), .S(n41708));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(clk32MHz), 
            .D(n42380), .S(n41784));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(clk32MHz), 
            .D(n42378), .S(n41730));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(clk32MHz), 
            .D(n7_adj_3156), .S(n8_adj_3133));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(clk32MHz), 
            .D(n7_adj_3157), .S(n8_adj_3132));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(clk32MHz), 
            .D(n42386), .S(n41788));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(clk32MHz), 
            .D(n7_adj_3158), .S(n8_adj_3131));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(clk32MHz), 
            .D(n28432), .S(n28845));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(clk32MHz), 
            .D(n28430), .S(n28843));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(clk32MHz), 
            .D(n42383), .S(n41790));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(clk32MHz), 
            .D(n42387), .S(n41724));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(clk32MHz), 
            .D(n42382), .S(n28841));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(clk32MHz), 
            .D(n42374), .S(n28839));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(clk32MHz), 
            .D(n28428), .S(n28837));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(clk32MHz), 
            .D(n42379), .S(n41792));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(clk32MHz), 
            .D(n42381), .S(n41794));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(clk32MHz), 
            .D(n42389), .S(n41796));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(clk32MHz), 
            .D(n42385), .S(n41722));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state_c [3]), .C(clk32MHz), 
            .D(n41720), .S(n41950));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n23790));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n23789));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n23438), .D(n43887));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(n22077), .I1(n38954), .I2(n10_adj_3159), 
            .I3(n1506), .O(n39131));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_848 (.I0(n22077), .I1(n38954), .I2(\data_out_frame[12] [5]), 
            .I3(GND_net), .O(n42549));
    defparam i1_2_lut_3_lut_adj_848.LUT_INIT = 16'h9696;
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n23438), .D(n43836));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n23438), .D(n42464));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n23438), .D(n43657));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n23438), .D(n43874));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n23438), .D(n43873));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n23438), .D(n42734));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n23438), .D(n42735));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n23438), .D(n44064));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n23438), .D(n43976));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n23438), .D(n43972));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n23438), .D(n42492));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n23438), .D(n43853));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n23438), .D(n43560));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n23438), .D(n43845));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n23438), .D(n43454));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_4_lut_adj_849 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(n23194), .I3(n10_adj_3160), .O(n42480));   // verilog/coms.v(71[16:34])
    defparam i5_3_lut_4_lut_adj_849.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n23788));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_850 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n42646));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_3_lut_adj_850.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n23787));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3150), .S(n3));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10491_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n23905));
    defparam i10491_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_851 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(n42471), .I3(n42806), .O(n22077));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_4_lut_adj_851.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_852 (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n22294));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_adj_852.LUT_INIT = 16'hbbbb;
    SB_LUT4 add_44_32_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n35885), .O(n2_adj_3161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15171_1_lut (.I0(n28564), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1498));
    defparam i15171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_44_11_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n35864), .O(n2_adj_3162)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_853 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(n42471), .I3(n23004), .O(n42803));   // verilog/coms.v(69[16:62])
    defparam i1_2_lut_4_lut_adj_853.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_854 (.I0(\data_out_frame[17] [4]), .I1(n23247), 
            .I2(n42584), .I3(n43500), .O(n43803));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_854.LUT_INIT = 16'h9669;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3161), .S(n3_adj_3163));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3164), .S(n3_adj_3165));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3166), .S(n3_adj_3167));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3168), .S(n3_adj_3169));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3170), .S(n3_adj_3171));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3172), .S(n3_adj_3173));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3174), .S(n3_adj_3175));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3176), .S(n3_adj_3177));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3178), .S(n3_adj_3179));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3180), .S(n3_adj_3181));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3182), .S(n3_adj_3183));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3184), .S(n3_adj_3185));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3186), .S(n3_adj_3187));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_c), .S(n3_adj_3188));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3118), .S(n3_adj_3189));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3125), .S(n3_adj_3190));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3129), .S(n3_adj_3191));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3135), .S(n3_adj_3192));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3139), .S(n3_adj_3193));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3142), .S(n3_adj_3194));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3147), .S(n3_adj_3195));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3162), .S(n3_adj_3196));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3197), .S(n3_adj_3198));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3199), .S(n3_adj_3200));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3201), .S(n3_adj_3202));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3117), .S(n3_adj_3203));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3123), .S(n3_adj_3204));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3137), .S(n3_adj_3205));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3141), .S(n3_adj_3206));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3148), .S(n3_adj_3207));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n23786));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_32 (.CI(n35885), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n35886));
    SB_LUT4 i1_2_lut_4_lut_adj_855 (.I0(\data_out_frame[5] [7]), .I1(n10_adj_3208), 
            .I2(\data_out_frame[9] [7]), .I3(n42688), .O(n39144));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_4_lut_adj_855.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_856 (.I0(\data_out_frame[5] [7]), .I1(n10_adj_3208), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[16] [7]), .O(n42849));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_4_lut_adj_856.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_31_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n35884), .O(n2_adj_3164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n24121));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n23785));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n24120));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n23784));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n24119));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n23783));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n23782));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n23781));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34330 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n49896));
    defparam byte_transmit_counter_0__bdd_4_lut_34330.LUT_INIT = 16'he4aa;
    SB_CARRY add_44_31 (.CI(n35884), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n35885));
    SB_LUT4 n49896_bdd_4_lut (.I0(n49896), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n49899));
    defparam n49896_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n23780));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_30_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n35883), .O(n2_adj_3166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10492_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42403), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n23906));
    defparam i10492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_30 (.CI(n35883), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n35884));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34325 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n49890));
    defparam byte_transmit_counter_0__bdd_4_lut_34325.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n23779));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n23778));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n23777));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n23776));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n23775));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_29_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n35882), .O(n2_adj_3168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_29 (.CI(n35882), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n35883));
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n23774));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n23773));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n23772));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n23771));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n23770));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n23769));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n23768));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n23767));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n23766));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n23765));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n23764));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_28_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n35881), .O(n2_adj_3170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 equal_63_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3121));   // verilog/coms.v(154[7:23])
    defparam equal_63_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n23763));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n23762));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_28 (.CI(n35881), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n35882));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_857 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42403), .I3(\FRAME_MATCHER.i [0]), .O(n20195));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_857.LUT_INIT = 16'hfbff;
    SB_LUT4 add_44_27_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n35880), .O(n2_adj_3172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n24133));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49890_bdd_4_lut (.I0(n49890), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n49893));
    defparam n49890_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_858 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42419), .I3(\FRAME_MATCHER.i [0]), .O(n42422));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_858.LUT_INIT = 16'hfbff;
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n23761));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_859 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42411), .I3(\FRAME_MATCHER.i [0]), .O(n20420));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_859.LUT_INIT = 16'hfbff;
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n23760));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_27 (.CI(n35880), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n35881));
    SB_LUT4 i1_2_lut_adj_860 (.I0(\data_in_frame[15] [4]), .I1(n23064), 
            .I2(GND_net), .I3(GND_net), .O(n42717));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_860.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34320 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n49884));
    defparam byte_transmit_counter_0__bdd_4_lut_34320.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_861 (.I0(n42926), .I1(n7_adj_3209), .I2(\data_in_frame[12] [2]), 
            .I3(n43035), .O(n10_adj_3210));
    defparam i4_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[8] [0]), .I1(n10_adj_3210), .I2(\data_in_frame[10] [0]), 
            .I3(GND_net), .O(n38377));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n23759));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_11 (.CI(n35864), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n35865));
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n23758));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n23757));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n23756));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n23755));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n23754));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n23753));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n23752));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n26838));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n23750));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n23749));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n23748));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n23747));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n23746));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n23745));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n23744));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n27693));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n27746));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n23741));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n23740));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n23739));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n23738));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n23737));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n28334));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n28366));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n23734));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n23733));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_26_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n35879), .O(n2_adj_3174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_862 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[17] [0]), 
            .I2(n22745), .I3(\data_in_frame[16] [6]), .O(n42742));
    defparam i3_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state_c [1]), .C(clk32MHz), 
           .D(n49980));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state[2] ), .C(clk32MHz), 
           .D(n49981));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10357_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n23771));
    defparam i10357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut (.I0(\data_in_frame[12] [6]), .I1(n42742), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3211));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut (.I0(\data_in_frame[17] [1]), .I1(n38377), .I2(n42941), 
            .I3(n22611), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_863 (.I0(\data_in_frame[19] [2]), .I1(n14), .I2(n10_adj_3211), 
            .I3(n43038), .O(n42843));
    defparam i7_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i10358_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n23772));
    defparam i10358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_864 (.I0(\data_in_frame[8]_c [1]), .I1(n42793), 
            .I2(n39163), .I3(n42910), .O(n26));
    defparam i11_4_lut_adj_864.LUT_INIT = 16'h9669;
    SB_CARRY add_44_26 (.CI(n35879), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n35880));
    SB_LUT4 i9_4_lut (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[18] [7]), 
            .I2(n23244), .I3(\data_in_frame[12][4] ), .O(n24));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10359_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n23773));
    defparam i10359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49884_bdd_4_lut (.I0(n49884), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n49887));
    defparam n49884_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34315 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n49878));
    defparam byte_transmit_counter_0__bdd_4_lut_34315.LUT_INIT = 16'he4aa;
    SB_LUT4 n49878_bdd_4_lut (.I0(n49878), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n49881));
    defparam n49878_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34310 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n49872));
    defparam byte_transmit_counter_0__bdd_4_lut_34310.LUT_INIT = 16'he4aa;
    SB_LUT4 n49872_bdd_4_lut (.I0(n49872), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n49875));
    defparam n49872_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34305 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n49866));
    defparam byte_transmit_counter_0__bdd_4_lut_34305.LUT_INIT = 16'he4aa;
    SB_LUT4 n49866_bdd_4_lut (.I0(n49866), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n49869));
    defparam n49866_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34300 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n49860));
    defparam byte_transmit_counter_0__bdd_4_lut_34300.LUT_INIT = 16'he4aa;
    SB_LUT4 n49860_bdd_4_lut (.I0(n49860), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n49863));
    defparam n49860_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34295 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n49854));
    defparam byte_transmit_counter_0__bdd_4_lut_34295.LUT_INIT = 16'he4aa;
    SB_LUT4 n49854_bdd_4_lut (.I0(n49854), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n49857));
    defparam n49854_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10_4_lut_adj_865 (.I0(n22723), .I1(n43032), .I2(n7_adj_3209), 
            .I3(n38367), .O(n25));
    defparam i10_4_lut_adj_865.LUT_INIT = 16'h6996;
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n24132));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i8_3_lut (.I0(n42742), .I1(\data_in_frame[19] [1]), .I2(n43011), 
            .I3(GND_net), .O(n23));
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut (.I0(n23), .I1(n25), .I2(n24), .I3(n26), .O(n42796));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34290 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n49848));
    defparam byte_transmit_counter_0__bdd_4_lut_34290.LUT_INIT = 16'he4aa;
    SB_DFF data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk32MHz), 
           .D(n24068));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n49848_bdd_4_lut (.I0(n49848), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n49851));
    defparam n49848_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk32MHz), 
           .D(n24067));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSR tx_transmit_3227 (.Q(r_SM_Main_2__N_2756[0]), .C(clk32MHz), 
            .D(n46769), .R(n42202));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n24109));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk32MHz), 
           .D(n24066));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_866 (.I0(\data_in_frame[10] [3]), .I1(n42536), 
            .I2(n43029), .I3(n6_adj_3212), .O(n43745));
    defparam i4_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n43745), .I1(n42923), .I2(\data_in_frame[16] [7]), 
            .I3(n22993), .O(n12));   // verilog/coms.v(76[16:27])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_44_3 (.CI(n35856), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n35857));
    SB_LUT4 add_44_25_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n35878), .O(n2_adj_3176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n24065));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n24108));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10360_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n23774));
    defparam i10360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_10_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n35863), .O(n2_adj_3197)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n24131));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_867 (.I0(n38426), .I1(n12), .I2(\data_in_frame[19] [3]), 
            .I3(n42678), .O(n42545));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_867.LUT_INIT = 16'h6996;
    SB_LUT4 i10361_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n23775));
    defparam i10361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_868 (.I0(\data_in_frame[16] [4]), .I1(n43056), 
            .I2(\data_in_frame[16] [6]), .I3(\data_in_frame[19] [0]), .O(n10_adj_3213));
    defparam i4_4_lut_adj_868.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_869 (.I0(\data_in_frame[14] [3]), .I1(n10_adj_3213), 
            .I2(n43038), .I3(GND_net), .O(n39117));
    defparam i5_3_lut_adj_869.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34285 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n49836));
    defparam byte_transmit_counter_0__bdd_4_lut_34285.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_870 (.I0(n42591), .I1(n42796), .I2(n42953), .I3(n42843), 
            .O(n8_adj_3214));
    defparam i3_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_871 (.I0(n42545), .I1(n8_adj_3214), .I2(n42840), 
            .I3(n42947), .O(n39161));
    defparam i4_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n24130));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_10 (.CI(n35863), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n35864));
    SB_CARRY add_44_25 (.CI(n35878), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n35879));
    SB_DFF Kd_i1 (.Q(\Kd[1] ), .C(clk32MHz), .D(n24129));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i2 (.Q(\Kd[2] ), .C(clk32MHz), .D(n24128));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i3 (.Q(\Kd[3] ), .C(clk32MHz), .D(n24127));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i4 (.Q(\Kd[4] ), .C(clk32MHz), .D(n24126));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i5 (.Q(\Kd[5] ), .C(clk32MHz), .D(n24125));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i6 (.Q(\Kd[6] ), .C(clk32MHz), .D(n24124));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE LED_3230 (.Q(LED_c), .C(clk32MHz), .E(n43084), .D(n22299));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10362_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n23776));
    defparam i10362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10363_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n23777));
    defparam i10363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_872 (.I0(\data_in_frame[13] [5]), .I1(n8_adj_3215), 
            .I2(n43008), .I3(n43069), .O(n39133));
    defparam i4_4_lut_adj_872.LUT_INIT = 16'h9669;
    SB_LUT4 n49836_bdd_4_lut (.I0(n49836), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n49839));
    defparam n49836_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_873 (.I0(n42879), .I1(n42998), .I2(GND_net), 
            .I3(GND_net), .O(n43056));
    defparam i1_2_lut_adj_873.LUT_INIT = 16'h6666;
    SB_LUT4 i10364_3_lut_4_lut (.I0(n8_adj_3121), .I1(n42419), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n23778));
    defparam i10364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10613_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[22]), .I3(\data_out_frame[9] [6]), .O(n24027));
    defparam i10613_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[7] [3]), 
            .I2(n42812), .I3(GND_net), .O(n43673));   // verilog/coms.v(77[16:35])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_874 (.I0(n42980), .I1(n43002), .I2(\data_in_frame[13] [7]), 
            .I3(n20947), .O(n12_adj_3216));
    defparam i5_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_875 (.I0(n38879), .I1(n12_adj_3216), .I2(n23013), 
            .I3(n43673), .O(Kp_23__N_176));
    defparam i6_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_876 (.I0(\data_in_frame[16] [3]), .I1(Kp_23__N_176), 
            .I2(GND_net), .I3(GND_net), .O(n22464));
    defparam i1_2_lut_adj_876.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_877 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42959));
    defparam i1_2_lut_adj_877.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_18__7__I_0_3252_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_786));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_18__7__I_0_3252_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_878 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23013));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_878.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_879 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42793));
    defparam i1_2_lut_adj_879.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_880 (.I0(n39163), .I1(n42793), .I2(n42457), .I3(\data_in_frame[16] [5]), 
            .O(n44171));
    defparam i3_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i15084_2_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28478));
    defparam i15084_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut (.I0(\FRAME_MATCHER.state_c [15]), .I1(\FRAME_MATCHER.state_c [5]), 
            .I2(\FRAME_MATCHER.state_c [21]), .I3(\FRAME_MATCHER.state_c [18]), 
            .O(n48));   // verilog/coms.v(152[5:27])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.state_c [24]), .I1(\FRAME_MATCHER.state_c [8]), 
            .I2(\FRAME_MATCHER.state_c [4]), .I3(\FRAME_MATCHER.state_c [7]), 
            .O(n46));   // verilog/coms.v(152[5:27])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.state_c [17]), .I1(\FRAME_MATCHER.state_c [20]), 
            .I2(\FRAME_MATCHER.state_c [10]), .I3(\FRAME_MATCHER.state_c [19]), 
            .O(n47));   // verilog/coms.v(152[5:27])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10648_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(control_mode[3]), .I3(\data_out_frame[5] [3]), .O(n24062));
    defparam i10648_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_881 (.I0(n23244), .I1(n42831), .I2(n42587), .I3(n44171), 
            .O(n38367));
    defparam i3_4_lut_adj_881.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.state_c [9]), .I1(\FRAME_MATCHER.state_c [11]), 
            .I2(\FRAME_MATCHER.state_c [26]), .I3(\FRAME_MATCHER.state_c [27]), 
            .O(n45_adj_3217));   // verilog/coms.v(152[5:27])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_44_24_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n35877), .O(n2_adj_3178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_882 (.I0(n22538), .I1(n42799), .I2(n42474), .I3(\data_in_frame[8][2] ), 
            .O(n22745));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.state_c [16]), .I1(\FRAME_MATCHER.state_c [12]), 
            .I2(\FRAME_MATCHER.state_c [23]), .I3(\FRAME_MATCHER.state_c [13]), 
            .O(n44));   // verilog/coms.v(152[5:27])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.state_c [28]), .I1(\FRAME_MATCHER.state_c [30]), 
            .I2(\FRAME_MATCHER.state_c [14]), .I3(\FRAME_MATCHER.state_c [25]), 
            .O(n43));   // verilog/coms.v(152[5:27])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 data_in_frame_12__7__I_0_3248_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_193));   // verilog/coms.v(69[16:27])
    defparam data_in_frame_12__7__I_0_3248_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i26_4_lut (.I0(n45_adj_3217), .I1(n47), .I2(n46), .I3(n48), 
            .O(n54));   // verilog/coms.v(152[5:27])
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(\FRAME_MATCHER.state_c [31]), .I1(\FRAME_MATCHER.state_c [6]), 
            .I2(\FRAME_MATCHER.state_c [22]), .I3(\FRAME_MATCHER.state_c [29]), 
            .O(n49_c));   // verilog/coms.v(152[5:27])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_c), .I1(n54), .I2(n43), .I3(n44), .O(n28987));   // verilog/coms.v(152[5:27])
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_44_24 (.CI(n35877), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n35878));
    SB_LUT4 i1_2_lut_adj_883 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42678));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_883.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_23_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n35876), .O(n2_adj_3180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n22274));
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h2222;
    SB_LUT4 i15_rep_4_2_lut (.I0(\FRAME_MATCHER.state_c [3]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49986));
    defparam i15_rep_4_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_885 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43005));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n49986), .I1(n28987), .I2(n4_c), .I3(n28478), 
            .O(n3346));
    defparam i1_4_lut.LUT_INIT = 16'h3032;
    SB_LUT4 i10626_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[1]), .I3(\data_out_frame[8] [1]), .O(n24040));
    defparam i10626_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10623_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[4]), .I3(\data_out_frame[8] [4]), .O(n24037));
    defparam i10623_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_886 (.I0(n22501), .I1(\data_in_frame[8]_c [3]), 
            .I2(\data_in_frame[6][1] ), .I3(GND_net), .O(n43059));   // verilog/coms.v(94[12:25])
    defparam i2_3_lut_adj_886.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_887 (.I0(n42666), .I1(n42910), .I2(GND_net), 
            .I3(GND_net), .O(n38426));
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_888 (.I0(n22589), .I1(n38426), .I2(\data_in_frame[14] [5]), 
            .I3(GND_net), .O(n38429));
    defparam i2_3_lut_adj_888.LUT_INIT = 16'h9696;
    SB_CARRY add_44_23 (.CI(n35876), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n35877));
    SB_LUT4 add_44_9_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n35862), .O(n2_adj_3199)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n24107));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_889 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n22701));
    defparam i1_2_lut_adj_889.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_2_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [0]), .I2(n164), 
            .I3(GND_net), .O(n2_adj_3218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n24106));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n24105));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_890 (.I0(\data_in_frame[8]_c [1]), .I1(n43035), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3219));
    defparam i1_2_lut_adj_890.LUT_INIT = 16'h6666;
    SB_CARRY add_44_9 (.CI(n35862), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n35863));
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n24104));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i10624_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[3]), .I3(\data_out_frame[8] [3]), .O(n24038));
    defparam i10624_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_891 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[9] [7]), 
            .I2(n38403), .I3(n6_adj_3219), .O(n42666));
    defparam i4_4_lut_adj_891.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_22_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n35875), .O(n2_adj_3182)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10583_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[12]), .I3(\data_out_frame[13] [4]), .O(n23997));
    defparam i10583_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_44_22 (.CI(n35875), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n35876));
    SB_LUT4 add_44_21_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n35874), .O(n2_adj_3184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10625_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[2]), .I3(\data_out_frame[8] [2]), .O(n24039));
    defparam i10625_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_CARRY add_44_21 (.CI(n35874), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n35875));
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n164), 
            .CO(n35856));
    SB_LUT4 add_44_20_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n35873), .O(n2_adj_3186)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3218), .S(n3_adj_3220));   // verilog/coms.v(126[12] 289[6])
    SB_DFF deadband_i0_i0 (.Q(deadband[0]), .C(clk32MHz), .D(n23585));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n23584));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
           .D(n41786));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n24029));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n23573));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n23572));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n23571));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n23570));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n23569));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kd_i0 (.Q(\Kd[0] ), .C(clk32MHz), .D(n23568));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n23567));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n23566));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n23565));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_8_lut (.I0(n1498), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n35861), .O(n2_adj_3201)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_892 (.I0(\data_in_frame[14] [1]), .I1(n42998), 
            .I2(n2), .I3(\data_in_frame[11] [5]), .O(n42812));
    defparam i3_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_893 (.I0(n23105), .I1(n38473), .I2(GND_net), 
            .I3(GND_net), .O(n43069));
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_894 (.I0(\data_in_frame[13] [3]), .I1(n23229), 
            .I2(\data_in_frame[10] [7]), .I3(GND_net), .O(n42530));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_adj_894.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_895 (.I0(n13), .I1(n23042), .I2(\data_in_frame[6] [5]), 
            .I3(\data_in_frame[8]_c [7]), .O(n42834));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_896 (.I0(n42614), .I1(n42834), .I2(\data_in_frame[11] [3]), 
            .I3(\data_in_frame[7] [1]), .O(n12_adj_3221));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_897 (.I0(\data_in_frame[9] [1]), .I1(n12_adj_3221), 
            .I2(n42983), .I3(n23178), .O(n23105));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42494));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_899 (.I0(n22960), .I1(n23105), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_866));
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_900 (.I0(n23007), .I1(n42834), .I2(n42530), .I3(n22960), 
            .O(n22698));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_901 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42923));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_902 (.I0(n42505), .I1(n42889), .I2(\data_in_frame[7] [2]), 
            .I3(\data_in_frame[4] [6]), .O(n39));
    defparam i7_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_903 (.I0(n43069), .I1(n42812), .I2(n42886), 
            .I3(n42666), .O(n51));
    defparam i19_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(\data_in_frame[12][4] ), .I1(n22701), .I2(\data_in_frame[13] [1]), 
            .I3(n38429), .O(n56));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n42855), .I1(n42675), .I2(n42681), .I3(n42608), 
            .O(n54_adj_3222));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10627_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[0]), .I3(\data_out_frame[8] [0]), .O(n24041));
    defparam i10627_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10628_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[15]), .I3(\data_out_frame[7] [7]), .O(n24042));
    defparam i10628_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i23_4_lut (.I0(n42530), .I1(n22954), .I2(n42494), .I3(\data_in_frame[4] [6]), 
            .O(n55));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_904 (.I0(\data_in_frame[15] [0]), .I1(n42896), 
            .I2(n43059), .I3(n42861), .O(n53_adj_3223));
    defparam i21_4_lut_adj_904.LUT_INIT = 16'h6996;
    SB_LUT4 i10629_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[14]), .I3(\data_out_frame[7] [6]), .O(n24043));
    defparam i10629_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i18_4_lut_adj_905 (.I0(n43005), .I1(\data_in_frame[9] [2]), 
            .I2(n42678), .I3(\data_in_frame[12] [2]), .O(n50));
    defparam i18_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut_adj_906 (.I0(n51), .I1(n39), .I2(Kp_23__N_193), 
            .I3(\data_in_frame[13] [0]), .O(n58));
    defparam i26_4_lut_adj_906.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n53_adj_3223), .I1(n55), .I2(n54_adj_3222), 
            .I3(n56), .O(n62));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10630_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[13]), .I3(\data_out_frame[7] [5]), .O(n24044));
    defparam i10630_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i17_4_lut_adj_907 (.I0(\data_in_frame[15] [2]), .I1(n42858), 
            .I2(n42559), .I3(\data_in_frame[12] [0]), .O(n49_adj_3224));
    defparam i17_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n49_adj_3224), .I1(n62), .I2(n58), .I3(n50), 
            .O(n39163));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_908 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22723));   // verilog/coms.v(83[17:63])
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_909 (.I0(n23244), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3225));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_910 (.I0(n43044), .I1(n42466), .I2(\data_in_frame[18] [2]), 
            .I3(n6_adj_3225), .O(n42956));   // verilog/coms.v(72[16:43])
    defparam i4_4_lut_adj_910.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_911 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[17] [5]), 
            .I2(n42956), .I3(n42457), .O(n28));
    defparam i10_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_912 (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n22421), .I3(GND_net), .O(n22424));
    defparam i1_2_lut_3_lut_adj_912.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_913 (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n22289), .I3(GND_net), .O(n22303));
    defparam i1_2_lut_3_lut_adj_913.LUT_INIT = 16'hf7f7;
    SB_LUT4 i14_3_lut (.I0(\data_in_frame[17] [7]), .I1(n28), .I2(n38367), 
            .I3(GND_net), .O(n32));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut (.I0(n39163), .I1(n42819), .I2(\data_in_frame[18] [3]), 
            .I3(n42923), .O(n30));
    defparam i12_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[16] [5]), .I1(n42867), .I2(\data_in_frame[17] [0]), 
            .I3(\data_in_frame[17] [6]), .O(n31_adj_3226));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_914 (.I0(Kp_23__N_786), .I1(n42524), .I2(n42959), 
            .I3(n44171), .O(n29));
    defparam i11_4_lut_adj_914.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_915 (.I0(n29), .I1(n31_adj_3226), .I2(n30), 
            .I3(n32), .O(n39122));
    defparam i17_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i10633_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[10]), .I3(\data_out_frame[7] [2]), .O(n24047));
    defparam i10633_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10634_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[9]), .I3(\data_out_frame[7] [1]), .O(n24048));
    defparam i10634_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_916 (.I0(\data_in_frame[19] [6]), .I1(n42995), 
            .I2(Kp_23__N_193), .I3(n22745), .O(n10_adj_3227));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_917 (.I0(n42864), .I1(n10_adj_3227), .I2(\data_in_frame[17] [4]), 
            .I3(GND_net), .O(n42747));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_917.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_918 (.I0(n39122), .I1(n42995), .I2(n42522), .I3(n42575), 
            .O(n12_adj_3228));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_918.LUT_INIT = 16'h6996;
    SB_LUT4 i17_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/coms.v(153[9:50])
    defparam i17_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_919 (.I0(\data_in_frame[15] [5]), .I1(n12_adj_3228), 
            .I2(\data_in_frame[19] [7]), .I3(n42861), .O(n42591));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i10636_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[23]), .I3(\data_out_frame[6] [7]), .O(n24050));
    defparam i10636_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 equal_1011_i7_2_lut (.I0(Kp_23__N_459), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3209));   // verilog/coms.v(230[9:81])
    defparam equal_1011_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10635_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[8]), .I3(\data_out_frame[7] [0]), .O(n24049));
    defparam i10635_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_920 (.I0(\data_in_frame[1] [3]), .I1(n42508), .I2(\data_in_frame[5] [5]), 
            .I3(GND_net), .O(n22501));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_920.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_921 (.I0(n28404), .I1(n10), .I2(GND_net), .I3(GND_net), 
            .O(n42403));
    defparam i1_2_lut_adj_921.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_922 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n22594));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_922.LUT_INIT = 16'h6666;
    SB_LUT4 i10579_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[0]), .I3(\data_out_frame[14] [0]), .O(n23993));
    defparam i10579_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_923 (.I0(n42575), .I1(n42784), .I2(n23007), .I3(n6_adj_3229), 
            .O(n42864));   // verilog/coms.v(72[16:43])
    defparam i4_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(Kp_23__N_379), .I1(\data_in_frame[5] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3120));   // verilog/coms.v(94[12:25])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_924 (.I0(n22589), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[15] [0]), .I3(GND_net), .O(n42941));
    defparam i2_3_lut_adj_924.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_925 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[5] [6]), 
            .I2(Kp_23__N_459), .I3(\data_in_frame[10] [4]), .O(n42799));   // verilog/coms.v(83[17:70])
    defparam i3_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_in_frame[12] [5]), .I1(n42799), 
            .I2(GND_net), .I3(GND_net), .O(n42974));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_927 (.I0(Kp_23__N_379), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n42920));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_927.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_928 (.I0(\data_in_frame[14] [7]), .I1(n42974), 
            .I2(\data_in_frame[10] [5]), .I3(\data_in_frame[15] [1]), .O(n42675));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i10637_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[22]), .I3(\data_out_frame[6] [6]), .O(n24051));
    defparam i10637_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10580_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[15]), .I3(\data_out_frame[13] [7]), .O(n23994));
    defparam i10580_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_929 (.I0(\data_in_frame[8]_c [4]), .I1(\data_in_frame[13] [2]), 
            .I2(\data_in_frame[8]_c [6]), .I3(n6_adj_3230), .O(n42886));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_929.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_930 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22954));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_930.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_931 (.I0(\data_in_frame[4] [1]), .I1(n42736), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[2] [0]), .O(n22554));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_932 (.I0(n22554), .I1(\data_in_frame[6] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n42536));
    defparam i1_2_lut_adj_932.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_933 (.I0(\data_in_frame[8]_c [3]), .I1(Kp_23__N_379), 
            .I2(\data_in_frame[5] [7]), .I3(n42536), .O(n42474));
    defparam i3_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_934 (.I0(n42608), .I1(\data_in_frame[8]_c [4]), 
            .I2(\data_in_frame[6] [3]), .I3(GND_net), .O(n42784));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_934.LUT_INIT = 16'h9696;
    SB_LUT4 i10638_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[21]), .I3(\data_out_frame[6] [5]), .O(n24052));
    defparam i10638_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_935 (.I0(\data_in_frame[10] [7]), .I1(n23007), 
            .I2(GND_net), .I3(GND_net), .O(n42611));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_935.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_936 (.I0(\data_in_frame[10] [5]), .I1(n42784), 
            .I2(n42474), .I3(\data_in_frame[6][1] ), .O(n22611));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_937 (.I0(\data_in_frame[3] [7]), .I1(n42567), .I2(\data_in_frame[3] [6]), 
            .I3(\data_in_frame[4] [0]), .O(n22538));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_937.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_938 (.I0(\data_in_frame[6] [2]), .I1(n22538), .I2(GND_net), 
            .I3(GND_net), .O(n23049));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_938.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_939 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [1]), 
            .I2(n23309), .I3(GND_net), .O(n23229));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_939.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_in_frame[11] [0]), .I1(n42886), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3231));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_941 (.I0(n23229), .I1(n23049), .I2(\data_in_frame[8]_c [7]), 
            .I3(n6_adj_3231), .O(n23064));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_942 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42867));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_942.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_943 (.I0(n13), .I1(\data_in_frame[11] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n42855));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_944 (.I0(n42675), .I1(n42920), .I2(\data_in_frame[12] [7]), 
            .I3(n23007), .O(n12_adj_3232));   // verilog/coms.v(69[16:27])
    defparam i5_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_945 (.I0(n22594), .I1(n12_adj_3232), .I2(n43029), 
            .I3(n22501), .O(n22993));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i10581_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[14]), .I3(\data_out_frame[13] [6]), .O(n23995));
    defparam i10581_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_4_lut_adj_946 (.I0(\data_in_frame[15] [3]), .I1(n42867), 
            .I2(n23324), .I3(n23064), .O(n12_adj_3233));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i10639_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[20]), .I3(\data_out_frame[6] [4]), .O(n24053));
    defparam i10639_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6_4_lut_adj_947 (.I0(n22993), .I1(n12_adj_3233), .I2(\data_in_frame[19] [5]), 
            .I3(n42575), .O(n42947));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_948 (.I0(\data_in_frame[17] [2]), .I1(n42941), 
            .I2(\data_in_frame[17] [3]), .I3(n42611), .O(n12_adj_3234));   // verilog/coms.v(69[16:27])
    defparam i5_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_949 (.I0(\data_in_frame[14] [6]), .I1(n12_adj_3234), 
            .I2(\data_in_frame[19] [4]), .I3(n42864), .O(n42840));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i10582_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[13]), .I3(\data_out_frame[13] [5]), .O(n23996));
    defparam i10582_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_950 (.I0(n2), .I1(n42614), .I2(GND_net), .I3(GND_net), 
            .O(n42889));
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h6666;
    SB_LUT4 i10536_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[11]), .I3(\data_out_frame[19] [3]), .O(n23950));
    defparam i10536_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42516));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_952 (.I0(n38403), .I1(n42621), .I2(GND_net), 
            .I3(GND_net), .O(n20947));
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i10641_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[18]), .I3(\data_out_frame[6] [2]), .O(n24055));
    defparam i10641_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42858));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i10584_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[11]), .I3(\data_out_frame[13] [3]), .O(n23998));
    defparam i10584_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_954 (.I0(\data_in_frame[1] [6]), .I1(n42708), .I2(\data_in_frame[4] [2]), 
            .I3(GND_net), .O(n22657));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_954.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_955 (.I0(\data_in_frame[8]_c [6]), .I1(\data_in_frame[6] [5]), 
            .I2(n22657), .I3(\data_in_frame[6] [4]), .O(n42572));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_956 (.I0(\data_in_frame[7] [3]), .I1(n43002), .I2(n42892), 
            .I3(\data_in_frame[7] [2]), .O(n44074));
    defparam i3_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_957 (.I0(n15), .I1(n42572), .I2(\data_in_frame[9] [0]), 
            .I3(\data_in_frame[7] [0]), .O(n12_adj_3235));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_958 (.I0(\data_in_frame[9] [1]), .I1(n12_adj_3235), 
            .I2(n42858), .I3(\data_in_frame[6] [6]), .O(n22960));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_959 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3] [0]), 
            .I2(n42562), .I3(GND_net), .O(n8_adj_3236));   // verilog/coms.v(68[16:27])
    defparam i3_3_lut_adj_959.LUT_INIT = 16'h9696;
    SB_LUT4 i10566_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[21]), .I3(\data_out_frame[15] [5]), .O(n23980));
    defparam i10566_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 equal_1011_i16_4_lut (.I0(n23238), .I1(\data_in_frame[4] [7]), 
            .I2(n8_adj_3236), .I3(\data_in_frame[0] [7]), .O(n42614));   // verilog/coms.v(230[9:81])
    defparam equal_1011_i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10469_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n23883));
    defparam i10469_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_960 (.I0(\data_in_frame[5] [0]), .I1(n42562), .I2(n20914), 
            .I3(GND_net), .O(n42852));
    defparam i2_3_lut_adj_960.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_961 (.I0(\data_in_frame[0] [0]), .I1(n42443), .I2(n4_adj_3237), 
            .I3(\data_in_frame[4] [4]), .O(n13));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i10470_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n23884));
    defparam i10470_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_962 (.I0(n22941), .I1(n13), .I2(\data_in_frame[6] [6]), 
            .I3(GND_net), .O(n23309));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_962.LUT_INIT = 16'h9696;
    SB_LUT4 i10642_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[17]), .I3(\data_out_frame[6] [1]), .O(n24056));
    defparam i10642_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_963 (.I0(n22824), .I1(n42852), .I2(GND_net), 
            .I3(GND_net), .O(n1_c));
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_964 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n4_adj_3237));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_964.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_965 (.I0(\data_in_frame[4] [5]), .I1(n5_adj_3238), 
            .I2(n4_adj_3237), .I3(GND_net), .O(n22941));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_adj_965.LUT_INIT = 16'h9696;
    SB_LUT4 i10471_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n23885));
    defparam i10471_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_966 (.I0(\data_in_frame[6] [7]), .I1(n22941), .I2(GND_net), 
            .I3(GND_net), .O(n23178));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h6666;
    SB_LUT4 i10643_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[16]), .I3(\data_out_frame[6] [0]), .O(n24057));
    defparam i10643_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10586_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[9]), .I3(\data_out_frame[13] [1]), .O(n24000));
    defparam i10586_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_967 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42870));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_967.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42736));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_969 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n42708));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_969.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42443));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i10472_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n23886));
    defparam i10472_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_971 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [5]), .I3(GND_net), .O(n23238));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_971.LUT_INIT = 16'h9696;
    SB_LUT4 i10587_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[8]), .I3(\data_out_frame[13] [0]), .O(n24001));
    defparam i10587_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_972 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n5_adj_3238));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_972.LUT_INIT = 16'h9696;
    SB_LUT4 i10645_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(control_mode[6]), .I3(\data_out_frame[5] [6]), .O(n24059));
    defparam i10645_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_973 (.I0(n5_adj_3238), .I1(n23238), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_326));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_973.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_974 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42567));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_974.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_975 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42899));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_975.LUT_INIT = 16'h6666;
    SB_LUT4 i10588_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[23]), .I3(\data_out_frame[12] [7]), .O(n24002));
    defparam i10588_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10646_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(control_mode[5]), .I3(\data_out_frame[5] [5]), .O(n24060));
    defparam i10646_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10473_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n23887));
    defparam i10473_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_976 (.I0(\data_in_frame[0] [6]), .I1(n42567), 
            .I2(\data_in_frame[2] [6]), .I3(n18_adj_3239), .O(n30_adj_3240));   // verilog/coms.v(68[16:27])
    defparam i13_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_977 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_326), 
            .I2(n42787), .I3(n22629), .O(n28_adj_3241));   // verilog/coms.v(68[16:27])
    defparam i11_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_978 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n42708), .I3(\data_in_frame[0] [7]), .O(n29_adj_3242));   // verilog/coms.v(68[16:27])
    defparam i12_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_979 (.I0(n42736), .I1(n42508), .I2(n42870), 
            .I3(n42899), .O(n27_c));   // verilog/coms.v(68[16:27])
    defparam i10_4_lut_adj_979.LUT_INIT = 16'h6996;
    SB_LUT4 i10589_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[22]), .I3(\data_out_frame[12] [6]), .O(n24003));
    defparam i10589_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16_4_lut_adj_980 (.I0(n27_c), .I1(n29_adj_3242), .I2(n28_adj_3241), 
            .I3(n30_adj_3240), .O(n42562));   // verilog/coms.v(68[16:27])
    defparam i16_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_981 (.I0(n42562), .I1(\data_in_frame[5] [1]), .I2(n22837), 
            .I3(GND_net), .O(n2));
    defparam i2_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_982 (.I0(n2), .I1(n42980), .I2(\data_in_frame[7] [2]), 
            .I3(GND_net), .O(n42815));
    defparam i2_3_lut_adj_982.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_983 (.I0(n15), .I1(n42614), .I2(GND_net), .I3(GND_net), 
            .O(n42892));
    defparam i1_2_lut_adj_983.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_984 (.I0(\data_in_frame[11] [5]), .I1(n42892), 
            .I2(n42815), .I3(\data_in_frame[7] [1]), .O(n43008));
    defparam i3_4_lut_adj_984.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_985 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[7] [0]), 
            .I2(n42983), .I3(n42815), .O(n38473));
    defparam i3_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 i10474_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n23888));
    defparam i10474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10647_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(control_mode[4]), .I3(\data_out_frame[5] [4]), .O(n24061));
    defparam i10647_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_986 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[0] [5]), .O(n10_adj_3243));
    defparam i4_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3244));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31360_4_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[2]), 
            .O(n46920));   // verilog/coms.v(104[34:55])
    defparam i31360_4_lut.LUT_INIT = 16'h880a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3245));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_987 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42681));
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h6666;
    SB_LUT4 i28857_4_lut (.I0(n19_adj_3244), .I1(\data_out_frame[22] [0]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n44416));
    defparam i28857_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22629));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h6666;
    SB_LUT4 i10590_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[21]), .I3(\data_out_frame[12] [5]), .O(n24004));
    defparam i10590_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_989 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n20914));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_989.LUT_INIT = 16'h9696;
    SB_LUT4 i28858_3_lut (.I0(n49851), .I1(n44416), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44417));
    defparam i28858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10475_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[1]), 
            .I3(\data_in_frame[6][1] ), .O(n23889));
    defparam i10475_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i28829_4_lut (.I0(n5_adj_3245), .I1(n46920), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n44388));
    defparam i28829_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i28831_4_lut (.I0(n44388), .I1(n44417), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n44390));
    defparam i28831_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i3_4_lut_adj_990 (.I0(\data_in_frame[5] [4]), .I1(n42663), .I2(\data_in_frame[3] [2]), 
            .I3(n20914), .O(n5));
    defparam i3_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i28830_3_lut (.I0(n49953), .I1(n49959), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44389));
    defparam i28830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10591_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[20]), .I3(\data_out_frame[12] [4]), .O(n24005));
    defparam i10591_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_991 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[7] [5]), 
            .I2(n42926), .I3(n5), .O(n42879));
    defparam i3_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_992 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42649));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h6666;
    SB_LUT4 i10592_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[19]), .I3(\data_out_frame[12] [3]), .O(n24006));
    defparam i10592_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10593_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[18]), .I3(\data_out_frame[12] [2]), .O(n24007));
    defparam i10593_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10594_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[17]), .I3(\data_out_frame[12] [1]), .O(n24008));
    defparam i10594_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\data_in_frame[18] [3]), .I1(n39133), 
            .I2(GND_net), .I3(GND_net), .O(n42630));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_994 (.I0(n42649), .I1(n42879), .I2(\data_in_frame[14] [1]), 
            .I3(\data_in_frame[13] [6]), .O(n12_adj_3246));
    defparam i5_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_995 (.I0(n38473), .I1(n12_adj_3246), .I2(n43008), 
            .I3(\data_in_frame[14] [0]), .O(n38982));
    defparam i6_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i10596_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[7]), .I3(\data_out_frame[11] [7]), .O(n24010));
    defparam i10596_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_4_lut_adj_996 (.I0(\data_in_frame[14] [0]), .I1(n22960), 
            .I2(\data_in_frame[16] [0]), .I3(n44074), .O(n12_adj_3247));   // verilog/coms.v(68[16:27])
    defparam i5_4_lut_adj_996.LUT_INIT = 16'h9669;
    SB_LUT4 i10476_3_lut_4_lut (.I0(n8_adj_3124), .I1(n42403), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n23890));
    defparam i10476_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_997 (.I0(n42505), .I1(n12_adj_3247), .I2(n42828), 
            .I3(n22560), .O(n42466));   // verilog/coms.v(68[16:27])
    defparam i6_4_lut_adj_997.LUT_INIT = 16'h6996;
    SB_LUT4 i10597_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[6]), .I3(\data_out_frame[11] [6]), .O(n24011));
    defparam i10597_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i6_4_lut_adj_998 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3248));
    defparam i6_4_lut_adj_998.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_999 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3249));   // verilog/coms.v(232[13:35])
    defparam i6_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1000 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3250));
    defparam i5_4_lut_adj_1000.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1001 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [2]), .O(n13_adj_3251));   // verilog/coms.v(232[13:35])
    defparam i5_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_LUT4 i15020_4_lut (.I0(n13_adj_3251), .I1(n13_adj_3250), .I2(n14_adj_3249), 
            .I3(n14_adj_3248), .O(n28411));
    defparam i15020_4_lut.LUT_INIT = 16'h32fa;
    SB_LUT4 i4_4_lut_adj_1002 (.I0(n42466), .I1(\data_in_frame[16] [2]), 
            .I2(n38982), .I3(n42630), .O(n10_adj_3252));
    defparam i4_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1003 (.I0(\data_in_frame[18] [2]), .I1(n10_adj_3252), 
            .I2(\data_in_frame[20] [4]), .I3(GND_net), .O(n43318));
    defparam i5_3_lut_adj_1003.LUT_INIT = 16'h9696;
    SB_LUT4 i1812_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_3253));
    defparam i1812_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[21] [6]), .I1(n42840), .I2(n42947), 
            .I3(GND_net), .O(n42686));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1004 (.I0(n42591), .I1(n42747), .I2(\data_in_frame[20] [0]), 
            .I3(n39122), .O(n12_adj_3254));
    defparam i5_4_lut_adj_1004.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_1005 (.I0(\data_in_frame[17] [7]), .I1(n39133), 
            .I2(n43047), .I3(GND_net), .O(n8_adj_3255));
    defparam i3_3_lut_adj_1005.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1006 (.I0(Kp_23__N_866), .I1(n12_adj_3254), .I2(n42950), 
            .I3(n22560), .O(n43516));
    defparam i6_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i10598_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[5]), .I3(\data_out_frame[11] [5]), .O(n24012));
    defparam i10598_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_4_lut_adj_1007 (.I0(n39161), .I1(n42524), .I2(\data_in_frame[20] [7]), 
            .I3(n39117), .O(n12_adj_3256));
    defparam i5_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1008 (.I0(\data_in_frame[17] [7]), .I1(n42591), 
            .I2(n39122), .I3(\data_in_frame[20] [1]), .O(n43674));
    defparam i3_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i15182_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n22175), .I3(\FRAME_MATCHER.i [31]), .O(n2857));
    defparam i15182_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 i6_4_lut_adj_1009 (.I0(\data_in_frame[18] [7]), .I1(n12_adj_3256), 
            .I2(n42831), .I3(\data_in_frame[16] [5]), .O(n43338));
    defparam i6_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i10599_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[4]), .I3(\data_out_frame[11] [4]), .O(n24013));
    defparam i10599_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i28758_4_lut (.I0(n43674), .I1(n42460), .I2(n42796), .I3(\data_in_frame[21] [2]), 
            .O(n44317));
    defparam i28758_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i10600_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[3]), .I3(\data_out_frame[11] [3]), .O(n24014));
    defparam i10600_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_1010 (.I0(n42753), .I1(n22723), .I2(\data_in_frame[18] [5]), 
            .I3(n42959), .O(n10_adj_3257));
    defparam i4_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 i10601_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[2]), .I3(\data_out_frame[11] [2]), .O(n24015));
    defparam i10601_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_1011 (.I0(n42947), .I1(n42953), .I2(\data_in_frame[21] [7]), 
            .I3(GND_net), .O(n43536));
    defparam i2_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1012 (.I0(\data_in_frame[18] [4]), .I1(n22464), 
            .I2(\data_in_frame[16] [1]), .I3(n6_adj_3258), .O(n43313));
    defparam i4_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_LUT4 i28754_4_lut (.I0(n42545), .I1(n43318), .I2(n42840), .I3(\data_in_frame[21] [5]), 
            .O(n44313));
    defparam i28754_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i6_4_lut_adj_1013 (.I0(n42545), .I1(n42686), .I2(n42843), 
            .I3(\data_in_frame[21] [4]), .O(n22_adj_3259));
    defparam i6_4_lut_adj_1013.LUT_INIT = 16'h8448;
    SB_LUT4 i28756_4_lut (.I0(\data_in_frame[21] [3]), .I1(n43313), .I2(n42796), 
            .I3(n42843), .O(n44315));
    defparam i28756_4_lut.LUT_INIT = 16'hedde;
    SB_LUT4 i5_4_lut_adj_1014 (.I0(n38377), .I1(n43536), .I2(n10_adj_3257), 
            .I3(\data_in_frame[20] [6]), .O(n21));
    defparam i5_4_lut_adj_1014.LUT_INIT = 16'h8448;
    SB_LUT4 i5_3_lut_adj_1015 (.I0(\data_in_frame[20] [2]), .I1(n39133), 
            .I2(n42950), .I3(GND_net), .O(n14_adj_3260));
    defparam i5_3_lut_adj_1015.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1016 (.I0(n43047), .I1(\data_in_frame[15] [5]), 
            .I2(n42516), .I3(n43044), .O(n15_adj_3261));
    defparam i6_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_adj_3261), .I1(n42717), .I2(n14_adj_3260), 
            .I3(\data_in_frame[16] [0]), .O(n43672));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1017 (.I0(\data_in_frame[20] [3]), .I1(n43516), 
            .I2(n8_adj_3255), .I3(n42956), .O(n18_adj_3262));
    defparam i2_4_lut_adj_1017.LUT_INIT = 16'h2112;
    SB_LUT4 i10_4_lut_adj_1018 (.I0(n44317), .I1(\data_in_frame[21] [1]), 
            .I2(n43338), .I3(n39161), .O(n26_adj_3263));
    defparam i10_4_lut_adj_1018.LUT_INIT = 16'h4010;
    SB_LUT4 i14_4_lut_adj_1019 (.I0(n21), .I1(n44315), .I2(n22_adj_3259), 
            .I3(n44313), .O(n30_adj_3264));
    defparam i14_4_lut_adj_1019.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_1020 (.I0(n39161), .I1(n43672), .I2(n42460), 
            .I3(\data_in_frame[21] [0]), .O(n17_adj_3265));
    defparam i1_4_lut_adj_1020.LUT_INIT = 16'h2112;
    SB_LUT4 i15_4_lut_adj_1021 (.I0(n17_adj_3265), .I1(n30_adj_3264), .I2(n26_adj_3263), 
            .I3(n18_adj_3262), .O(Kp_23__N_152));
    defparam i15_4_lut_adj_1021.LUT_INIT = 16'h8000;
    SB_LUT4 equal_61_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3124));
    defparam equal_61_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i10602_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[1]), .I3(\data_out_frame[11] [1]), .O(n24016));
    defparam i10602_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10603_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[0]), .I3(\data_out_frame[11] [0]), .O(n24017));
    defparam i10603_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10604_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[15]), .I3(\data_out_frame[10] [7]), .O(n24018));
    defparam i10604_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10606_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[13]), .I3(\data_out_frame[10] [5]), .O(n24020));
    defparam i10606_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10605_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[14]), .I3(\data_out_frame[10] [6]), .O(n24019));
    defparam i10605_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10524_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[7]), .I3(\data_out_frame[20] [7]), .O(n23938));
    defparam i10524_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_1022 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(n22289), .I3(GND_net), .O(n63_adj_3266));   // verilog/coms.v(253[5:27])
    defparam i2_3_lut_adj_1022.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1023 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42403), .I3(\FRAME_MATCHER.i [0]), .O(n20471));
    defparam i1_2_lut_3_lut_4_lut_adj_1023.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1024 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42411), .I3(\FRAME_MATCHER.i [0]), .O(n42418));
    defparam i1_2_lut_3_lut_4_lut_adj_1024.LUT_INIT = 16'hf7ff;
    SB_LUT4 i10525_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[6]), .I3(\data_out_frame[20] [6]), .O(n23939));
    defparam i10525_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10532_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[15]), .I3(\data_out_frame[19] [7]), .O(n23946));
    defparam i10532_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15039_2_lut (.I0(Kp_23__N_152), .I1(n28411), .I2(GND_net), 
            .I3(GND_net), .O(n28433));
    defparam i15039_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i10526_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[5]), .I3(\data_out_frame[20] [5]), .O(n23940));
    defparam i10526_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10527_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[4]), .I3(\data_out_frame[20] [4]), .O(n23941));
    defparam i10527_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10529_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[2]), .I3(\data_out_frame[20] [2]), .O(n23943));
    defparam i10529_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10530_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[1]), .I3(\data_out_frame[20] [1]), .O(n23944));
    defparam i10530_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10531_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[0]), .I3(\data_out_frame[20] [0]), .O(n23945));
    defparam i10531_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10533_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[14]), .I3(\data_out_frame[19] [6]), .O(n23947));
    defparam i10533_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10534_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[13]), .I3(\data_out_frame[19] [5]), .O(n23948));
    defparam i10534_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10535_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[12]), .I3(\data_out_frame[19] [4]), .O(n23949));
    defparam i10535_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10537_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[10]), .I3(\data_out_frame[19] [2]), .O(n23951));
    defparam i10537_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10538_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[9]), .I3(\data_out_frame[19] [1]), .O(n23952));
    defparam i10538_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[16] [0]), .O(n3790));
    defparam mux_921_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10539_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[8]), .I3(\data_out_frame[19] [0]), .O(n23953));
    defparam i10539_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10544_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[19]), .I3(\data_out_frame[18] [3]), .O(n23958));
    defparam i10544_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16_2_lut (.I0(n407), .I1(\PID_CONTROLLER.result[13] ), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(32[23:29])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10540_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[23]), .I3(\data_out_frame[18] [7]), .O(n23954));
    defparam i10540_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10541_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[22]), .I3(\data_out_frame[18] [6]), .O(n23955));
    defparam i10541_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10542_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[21]), .I3(\data_out_frame[18] [5]), .O(n23956));
    defparam i10542_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[16] [1]), .O(n3791));
    defparam mux_921_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[16] [2]), .O(n3792));
    defparam mux_921_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34276 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n49830));
    defparam byte_transmit_counter_0__bdd_4_lut_34276.LUT_INIT = 16'he4aa;
    SB_LUT4 i10543_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[20]), .I3(\data_out_frame[18] [4]), .O(n23957));
    defparam i10543_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10545_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[18]), .I3(\data_out_frame[18] [2]), .O(n23959));
    defparam i10545_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10546_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[17]), .I3(\data_out_frame[18] [1]), .O(n23960));
    defparam i10546_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[16] [3]), .O(n3793));
    defparam mux_921_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10547_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[16]), .I3(\data_out_frame[18] [0]), .O(n23961));
    defparam i10547_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10549_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[6]), .I3(\data_out_frame[17] [6]), .O(n23963));
    defparam i10549_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10554_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[1]), .I3(\data_out_frame[17] [1]), .O(n23968));
    defparam i10554_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n49830_bdd_4_lut (.I0(n49830), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n49833));
    defparam n49830_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_921_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[16] [4]), .O(n3794));
    defparam mux_921_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10550_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[5]), .I3(\data_out_frame[17] [5]), .O(n23964));
    defparam i10550_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10551_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[4]), .I3(\data_out_frame[17] [4]), .O(n23965));
    defparam i10551_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2024_2_lut (.I0(n3346), .I1(\FRAME_MATCHER.state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n5017));
    defparam i2024_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i10552_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[3]), .I3(\data_out_frame[17] [3]), .O(n23966));
    defparam i10552_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34271 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n49824));
    defparam byte_transmit_counter_0__bdd_4_lut_34271.LUT_INIT = 16'he4aa;
    SB_LUT4 i10553_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[2]), .I3(\data_out_frame[17] [2]), .O(n23967));
    defparam i10553_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10555_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[0]), .I3(\data_out_frame[17] [0]), .O(n23969));
    defparam i10555_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[16] [5]), .O(n3795));
    defparam mux_921_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[16] [6]), .O(n3796));
    defparam mux_921_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[16] [7]), .O(n3797));
    defparam mux_921_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10557_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[14]), .I3(\data_out_frame[16] [6]), .O(n23971));
    defparam i10557_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10559_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[12]), .I3(\data_out_frame[16] [4]), .O(n23973));
    defparam i10559_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10560_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[11]), .I3(\data_out_frame[16] [3]), .O(n23974));
    defparam i10560_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i23_4_lut_adj_1025 (.I0(n3831), .I1(n30654), .I2(n45), .I3(byte_transmit_counter[7]), 
            .O(n24177));
    defparam i23_4_lut_adj_1025.LUT_INIT = 16'hcac0;
    SB_LUT4 i10561_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[10]), .I3(\data_out_frame[16] [2]), .O(n23975));
    defparam i10561_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10562_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[9]), .I3(\data_out_frame[16] [1]), .O(n23976));
    defparam i10562_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10563_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[8]), .I3(\data_out_frame[16] [0]), .O(n23977));
    defparam i10563_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10564_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[23]), .I3(\data_out_frame[15] [7]), .O(n23978));
    defparam i10564_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[15] [0]), .O(n3798));
    defparam mux_921_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10565_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[22]), .I3(\data_out_frame[15] [6]), .O(n23979));
    defparam i10565_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10567_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[20]), .I3(\data_out_frame[15] [4]), .O(n23981));
    defparam i10567_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10568_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[19]), .I3(\data_out_frame[15] [3]), .O(n23982));
    defparam i10568_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[15] [1]), .O(n3799));
    defparam mux_921_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10569_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[18]), .I3(\data_out_frame[15] [2]), .O(n23983));
    defparam i10569_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10570_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[17]), .I3(\data_out_frame[15] [1]), .O(n23984));
    defparam i10570_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i17311_3_lut (.I0(n23411), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n23582));   // verilog/uart_tx.v(31[16:25])
    defparam i17311_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 mux_921_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[15] [2]), .O(n3800));
    defparam mux_921_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_2_lut_adj_1026 (.I0(deadband[13]), .I1(\PID_CONTROLLER.result[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_3));   // verilog/motorControl.v(32[23:29])
    defparam i17_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i10571_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[16]), .I3(\data_out_frame[15] [0]), .O(n23985));
    defparam i10571_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10572_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[7]), .I3(\data_out_frame[14] [7]), .O(n23986));
    defparam i10572_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10573_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[6]), .I3(\data_out_frame[14] [6]), .O(n23987));
    defparam i10573_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10574_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[5]), .I3(\data_out_frame[14] [5]), .O(n23988));
    defparam i10574_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10575_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[4]), .I3(\data_out_frame[14] [4]), .O(n23989));
    defparam i10575_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[15] [3]), .O(n3801));
    defparam mux_921_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3269));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31521_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n47082));   // verilog/coms.v(104[34:55])
    defparam i31521_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3270));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28827_4_lut (.I0(n19_adj_3269), .I1(\data_out_frame[22] [7]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n44386));
    defparam i28827_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28828_3_lut (.I0(n49839), .I1(n44386), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44387));
    defparam i28828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10576_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[3]), .I3(\data_out_frame[14] [3]), .O(n23990));
    defparam i10576_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i28853_4_lut (.I0(n5_adj_3270), .I1(n47082), .I2(n45253), 
            .I3(byte_transmit_counter[0]), .O(n44412));
    defparam i28853_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i28855_4_lut (.I0(n44412), .I1(n44387), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n44414));
    defparam i28855_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28854_3_lut (.I0(n49887), .I1(n49881), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44413));
    defparam i28854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3271));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31514_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n47075));   // verilog/coms.v(104[34:55])
    defparam i31514_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3272));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28824_4_lut (.I0(n19_adj_3271), .I1(\data_out_frame[22] [6]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n44383));
    defparam i28824_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28825_3_lut (.I0(n49833), .I1(n44383), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44384));
    defparam i28825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_2_lut (.I0(PWMLimit[13]), .I1(\PID_CONTROLLER.result[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4));   // verilog/motorControl.v(32[23:29])
    defparam i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28850_4_lut (.I0(n5_adj_3272), .I1(n47075), .I2(n45253), 
            .I3(byte_transmit_counter[0]), .O(n44409));
    defparam i28850_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i28852_4_lut (.I0(n44409), .I1(n44384), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n44411));
    defparam i28852_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28851_3_lut (.I0(n49899), .I1(n49893), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44410));
    defparam i28851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10618_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[17]), .I3(\data_out_frame[9] [1]), .O(n24032));
    defparam i10618_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10619_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[16]), .I3(\data_out_frame[9] [0]), .O(n24033));
    defparam i10619_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3274));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n47070));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3275));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28821_4_lut (.I0(n19_adj_3274), .I1(\data_out_frame[22] [5]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n44380));
    defparam i28821_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10577_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[2]), .I3(\data_out_frame[14] [2]), .O(n23991));
    defparam i10577_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i28822_3_lut (.I0(n49827), .I1(n44380), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44381));
    defparam i28822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28847_4_lut (.I0(n5_adj_3275), .I1(byte_transmit_counter[0]), 
            .I2(n45253), .I3(n47070), .O(n44406));
    defparam i28847_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i28849_4_lut (.I0(n44406), .I1(n44381), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n44408));
    defparam i28849_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28848_3_lut (.I0(n49911), .I1(n49905), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44407));
    defparam i28848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10578_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[1]), .I3(\data_out_frame[14] [1]), .O(n23992));
    defparam i10578_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10620_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[7]), .I3(\data_out_frame[8] [7]), .O(n24034));
    defparam i10620_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3276));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28818_4_lut (.I0(n19_adj_3276), .I1(\data_out_frame[22] [4]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n44377));
    defparam i28818_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33238_3_lut (.I0(n49869), .I1(n49875), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n48799));
    defparam i33238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28819_3_lut (.I0(n49821), .I1(n44377), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44378));
    defparam i28819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33242_3_lut (.I0(n49965), .I1(n48799), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n48803));   // verilog/coms.v(104[34:55])
    defparam i33242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33243_4_lut (.I0(n48803), .I1(n44378), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam i33243_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10621_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[6]), .I3(\data_out_frame[8] [6]), .O(n24035));
    defparam i10621_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10595_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[16]), .I3(\data_out_frame[12] [0]), .O(n24009));
    defparam i10595_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i31500_2_lut (.I0(\data_out_frame[0][3] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n46666));   // verilog/coms.v(104[34:55])
    defparam i31500_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n46666), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3277));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3278));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28838_3_lut (.I0(n5_adj_3278), .I1(n6_adj_3277), .I2(n45253), 
            .I3(GND_net), .O(n44397));
    defparam i28838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10650_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(control_mode[1]), .I3(\data_out_frame[5] [1]), .O(n24064));
    defparam i10650_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i28840_4_lut (.I0(n44397), .I1(n49971), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n44399));
    defparam i28840_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28839_3_lut (.I0(n49923), .I1(n49917), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44398));
    defparam i28839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10644_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(control_mode[7]), .I3(\data_out_frame[5] [7]), .O(n24058));
    defparam i10644_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i31894_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n46663));   // verilog/coms.v(104[34:55])
    defparam i31894_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3279));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5][2] ), 
            .I1(n46663), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3280));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha00c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3281));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28863_4_lut (.I0(n19_adj_3279), .I1(\data_out_frame[22] [2]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n44422));
    defparam i28863_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28864_3_lut (.I0(n49863), .I1(n44422), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44423));
    defparam i28864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28835_3_lut (.I0(n5_adj_3281), .I1(n6_adj_3280), .I2(n45253), 
            .I3(GND_net), .O(n44394));
    defparam i28835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28837_4_lut (.I0(n44394), .I1(n44423), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n44396));
    defparam i28837_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28836_3_lut (.I0(n49935), .I1(n49929), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44395));
    defparam i28836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10585_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(setpoint[10]), .I3(\data_out_frame[13] [2]), .O(n23999));
    defparam i10585_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10640_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[19]), .I3(\data_out_frame[6] [3]), .O(n24054));
    defparam i10640_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_921_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[15] [4]), .O(n3802));
    defparam mux_921_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10614_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[21]), .I3(\data_out_frame[9] [5]), .O(n24028));
    defparam i10614_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10612_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[23]), .I3(\data_out_frame[9] [7]), .O(n24026));
    defparam i10612_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3282));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31491_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n47051));   // verilog/coms.v(104[34:55])
    defparam i31491_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3283));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28860_4_lut (.I0(n19_adj_3282), .I1(\data_out_frame[22] [1]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n44419));
    defparam i28860_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28861_3_lut (.I0(n49857), .I1(n44419), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44420));
    defparam i28861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28832_4_lut (.I0(n5_adj_3283), .I1(n47051), .I2(n45253), 
            .I3(byte_transmit_counter[0]), .O(n44391));
    defparam i28832_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i28834_4_lut (.I0(n44391), .I1(n44420), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n44393));
    defparam i28834_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i28833_3_lut (.I0(n49947), .I1(n49941), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44392));
    defparam i28833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10611_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[8]), .I3(\data_out_frame[10] [0]), .O(n24025));
    defparam i10611_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10610_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[9]), .I3(\data_out_frame[10] [1]), .O(n24024));
    defparam i10610_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10609_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[10]), .I3(\data_out_frame[10] [2]), .O(n24023));
    defparam i10609_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n49824_bdd_4_lut (.I0(n49824), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n49827));
    defparam n49824_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_921_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[15] [5]), .O(n3803));
    defparam mux_921_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10558_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[13]), .I3(\data_out_frame[16] [5]), .O(n23972));
    defparam i10558_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10608_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[11]), .I3(\data_out_frame[10] [3]), .O(n24022));
    defparam i10608_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15_rep_279_2_lut (.I0(\pwm_23__N_2960[13] ), .I1(\PID_CONTROLLER.result[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n50261));   // verilog/motorControl.v(32[23:29])
    defparam i15_rep_279_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_599_i1_4_lut (.I0(n28433), .I1(n28971), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(\FRAME_MATCHER.state [0]), .O(n28985));   // verilog/coms.v(147[4] 288[11])
    defparam mux_599_i1_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i31210_4_lut (.I0(\FRAME_MATCHER.state_c [3]), .I1(n28985), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n4_adj_3284), .O(n46769));   // verilog/coms.v(147[4] 288[11])
    defparam i31210_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i10607_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[12]), .I3(\data_out_frame[10] [4]), .O(n24021));
    defparam i10607_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_adj_1027 (.I0(n5019), .I1(n43149), .I2(\FRAME_MATCHER.state_31__N_1925 [3]), 
            .I3(n5017), .O(n23444));
    defparam i1_4_lut_adj_1027.LUT_INIT = 16'ha022;
    SB_LUT4 mux_921_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[15] [6]), .O(n3804));
    defparam mux_921_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[15] [7]), .O(n3805));
    defparam mux_921_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[14] [0]), .O(n3806));
    defparam mux_921_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10616_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[19]), .I3(\data_out_frame[9] [3]), .O(n24030));
    defparam i10616_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10556_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[15]), .I3(\data_out_frame[16] [7]), .O(n23970));
    defparam i10556_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10617_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[18]), .I3(\data_out_frame[9] [2]), .O(n24031));
    defparam i10617_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i15202_3_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n63_adj_3143), 
            .I2(n63_c), .I3(GND_net), .O(n123));   // verilog/coms.v(139[4] 142[7])
    defparam i15202_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i3644_2_lut (.I0(n63), .I1(n740), .I2(GND_net), .I3(GND_net), 
            .O(n16810));   // verilog/coms.v(157[6] 159[9])
    defparam i3644_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1028 (.I0(n63), .I1(n2857), .I2(n124), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_1989[1] ));
    defparam i2_3_lut_adj_1028.LUT_INIT = 16'hfdfd;
    SB_LUT4 i10632_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[11]), .I3(\data_out_frame[7] [3]), .O(n24046));
    defparam i10632_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10548_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(pwm[7]), .I3(\data_out_frame[17] [7]), .O(n23962));
    defparam i10548_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i28806_4_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [4]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[2] [5]), .O(n44365));
    defparam i28806_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10631_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[12]), .I3(\data_out_frame[7] [4]), .O(n24045));
    defparam i10631_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10651_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(control_mode[0]), .I3(\data_out_frame[5] [0]), .O(n24065));
    defparam i10651_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10615_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder1_position[20]), .I3(\data_out_frame[9] [4]), .O(n24029));
    defparam i10615_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10622_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(encoder0_position[5]), .I3(\data_out_frame[8] [5]), .O(n24036));
    defparam i10622_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10528_3_lut_4_lut (.I0(\FRAME_MATCHER.state[2] ), .I1(n22277), 
            .I2(displacement[3]), .I3(\data_out_frame[20] [3]), .O(n23942));
    defparam i10528_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14_4_lut_adj_1029 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [4]), .O(n38));
    defparam i14_4_lut_adj_1029.LUT_INIT = 16'h8000;
    SB_LUT4 i15_4_lut_adj_1030 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[2] [6]), .O(n39_adj_3285));
    defparam i15_4_lut_adj_1030.LUT_INIT = 16'h0002;
    SB_LUT4 i13_4_lut_adj_1031 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [3]), .O(n37_adj_3286));
    defparam i13_4_lut_adj_1031.LUT_INIT = 16'h2000;
    SB_LUT4 i28802_4_lut (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [7]), .O(n44361));
    defparam i28802_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1032 (.I0(n37_adj_3286), .I1(n39_adj_3285), .I2(n38), 
            .I3(n44365), .O(n46_adj_3287));
    defparam i22_4_lut_adj_1032.LUT_INIT = 16'h0080;
    SB_LUT4 i28804_4_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[2] [7]), .O(n44363));
    defparam i28804_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_3_lut (.I0(n44363), .I1(n46_adj_3287), .I2(n44361), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_1925 [3]));
    defparam i23_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i2026_3_lut (.I0(n3346), .I1(\FRAME_MATCHER.state[2] ), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n5019));
    defparam i2026_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_adj_1033 (.I0(n5019), .I1(\FRAME_MATCHER.state_31__N_1925 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22277));
    defparam i1_2_lut_adj_1033.LUT_INIT = 16'h8888;
    SB_LUT4 mux_921_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[14] [1]), .O(n3807));
    defparam mux_921_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[14] [2]), .O(n3808));
    defparam mux_921_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[14] [3]), .O(n3809));
    defparam mux_921_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[14] [4]), .O(n3810));
    defparam mux_921_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[14] [5]), .O(n3811));
    defparam mux_921_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[14] [6]), .O(n3812));
    defparam mux_921_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_921_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28413), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[14] [7]), .O(n3813));
    defparam mux_921_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1034 (.I0(\data_in_frame[14] [4]), .I1(n38429), 
            .I2(n42666), .I3(n42910), .O(n43038));
    defparam i1_2_lut_3_lut_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1035 (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[18] [0]), 
            .I2(n23105), .I3(n38473), .O(n42950));
    defparam i1_2_lut_3_lut_4_lut_adj_1035.LUT_INIT = 16'h9669;
    SB_LUT4 i10453_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[7]), 
            .I3(\data_in_frame[8]_c [7]), .O(n23867));
    defparam i10453_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10151_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [0]), 
            .I3(IntegralLimit[0]), .O(n23565));
    defparam i10151_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1036 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(n42691), .I3(n6_adj_3288), .O(n43454));
    defparam i4_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1037 (.I0(n38418), .I1(n42902), .I2(n38867), 
            .I3(n38351), .O(n12_adj_3289));
    defparam i5_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1038 (.I0(\data_out_frame[20] [7]), .I1(n12_adj_3289), 
            .I2(n43017), .I3(n23136), .O(n43845));
    defparam i6_4_lut_adj_1038.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1039 (.I0(\data_out_frame[19] [1]), .I1(n1716), 
            .I2(n42758), .I3(n6_adj_3290), .O(n43560));
    defparam i4_4_lut_adj_1039.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1040 (.I0(n38867), .I1(n42491), .I2(\data_out_frame[19] [1]), 
            .I3(n23295), .O(n43853));
    defparam i3_4_lut_adj_1040.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1041 (.I0(\data_out_frame[17] [1]), .I1(n23136), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n42491));
    defparam i2_3_lut_adj_1041.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1042 (.I0(n39131), .I1(n42550), .I2(n22668), 
            .I3(n42849), .O(n10_adj_3291));
    defparam i4_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1043 (.I0(\data_out_frame[19] [3]), .I1(n38351), 
            .I2(n23295), .I3(GND_net), .O(n44169));
    defparam i2_3_lut_adj_1043.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1044 (.I0(n44169), .I1(n42731), .I2(\data_out_frame[17] [3]), 
            .I3(GND_net), .O(n43972));
    defparam i2_3_lut_adj_1044.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1045 (.I0(n23267), .I1(\data_out_frame[19] [4]), 
            .I2(\data_out_frame[17] [2]), .I3(GND_net), .O(n42731));
    defparam i2_3_lut_adj_1045.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1046 (.I0(n1444), .I1(\data_out_frame[6] [3]), 
            .I2(n42803), .I3(n1695), .O(n12_adj_3292));   // verilog/coms.v(72[16:27])
    defparam i5_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1047 (.I0(\data_out_frame[6] [1]), .I1(n12_adj_3292), 
            .I2(n42477), .I3(\data_out_frame[15] [0]), .O(n23295));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1048 (.I0(n23295), .I1(n42731), .I2(n42723), 
            .I3(\data_out_frame[17] [4]), .O(n43976));
    defparam i3_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1049 (.I0(\data_out_frame[13] [0]), .I1(n1509), 
            .I2(n42598), .I3(n1595), .O(n10_adj_3159));
    defparam i4_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(n38210), .I1(n39131), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3293));
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1051 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[14] [7]), 
            .I2(n38954), .I3(n6_adj_3293), .O(n38418));
    defparam i4_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1052 (.I0(n38418), .I1(\data_out_frame[19] [5]), 
            .I2(n22520), .I3(GND_net), .O(n42723));
    defparam i2_3_lut_adj_1052.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1053 (.I0(n42902), .I1(n42917), .I2(\data_out_frame[20] [0]), 
            .I3(n39149), .O(n12_adj_3294));
    defparam i5_4_lut_adj_1053.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1054 (.I0(n42723), .I1(n12_adj_3294), .I2(n43026), 
            .I3(n42595), .O(n44064));
    defparam i6_4_lut_adj_1054.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(n42533), .I1(n42734), .I2(GND_net), 
            .I3(GND_net), .O(n42735));
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1056 (.I0(\data_in_frame[18] [1]), .I1(n38982), 
            .I2(n42879), .I3(n42998), .O(n43044));
    defparam i1_2_lut_3_lut_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1057 (.I0(n42932), .I1(n42944), .I2(n22779), 
            .I3(\data_out_frame[16] [6]), .O(n12_adj_3295));
    defparam i5_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1058 (.I0(n43500), .I1(n12_adj_3295), .I2(n43041), 
            .I3(n39125), .O(n38867));
    defparam i6_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1059 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42932));
    defparam i1_2_lut_adj_1059.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1060 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[19] [3]), 
            .I2(\data_out_frame[19] [2]), .I3(\data_out_frame[19] [5]), 
            .O(n28_adj_3296));
    defparam i10_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1061 (.I0(n43065), .I1(n42876), .I2(n43020), 
            .I3(\data_out_frame[18] [6]), .O(n31_adj_3297));
    defparam i13_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1062 (.I0(n38811), .I1(n42751), .I2(n43026), 
            .I3(n23251), .O(n30_adj_3298));
    defparam i12_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1063 (.I0(n31_adj_3297), .I1(\data_out_frame[18] [3]), 
            .I2(n28_adj_3296), .I3(\data_out_frame[18] [5]), .O(n34));
    defparam i16_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1064 (.I0(\data_out_frame[19] [4]), .I1(n42932), 
            .I2(n22674), .I3(\data_out_frame[18] [4]), .O(n29_adj_3299));
    defparam i11_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1065 (.I0(n23345), .I1(n29_adj_3299), .I2(n34), 
            .I3(n30_adj_3298), .O(n43017));
    defparam i1_4_lut_adj_1065.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1066 (.I0(\data_out_frame[16] [4]), .I1(n38867), 
            .I2(\data_out_frame[18] [7]), .I3(\data_out_frame[19] [0]), 
            .O(n42758));
    defparam i3_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(n22077), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43041));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1068 (.I0(n38811), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[16] [5]), .I3(GND_net), .O(n42929));
    defparam i2_3_lut_adj_1068.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1069 (.I0(n22019), .I1(n42720), .I2(\data_out_frame[20] [4]), 
            .I3(n42764), .O(n16_adj_3300));
    defparam i6_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1070 (.I0(n42542), .I1(n42761), .I2(\data_out_frame[16] [0]), 
            .I3(n42694), .O(n17_adj_3301));
    defparam i7_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1071 (.I0(n17_adj_3301), .I1(n21999), .I2(n16_adj_3300), 
            .I3(\data_out_frame[20] [7]), .O(n42595));
    defparam i9_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1072 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[12] [5]), 
            .I2(n42929), .I3(GND_net), .O(n14_adj_3302));
    defparam i5_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1073 (.I0(n43041), .I1(\data_out_frame[18] [5]), 
            .I2(n42758), .I3(n43017), .O(n15_adj_3303));
    defparam i6_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1074 (.I0(n15_adj_3303), .I1(n42849), .I2(n14_adj_3302), 
            .I3(n23114), .O(n38353));
    defparam i8_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(n38353), .I1(n22017), .I2(n42595), 
            .I3(n39189), .O(n42734));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1076 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[6] [0]), 
            .I2(Kp_23__N_379), .I3(\data_in_frame[5] [7]), .O(n42910));
    defparam i1_2_lut_3_lut_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1077 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[6] [4]), 
            .I2(n42803), .I3(GND_net), .O(n14_adj_3304));   // verilog/coms.v(73[16:27])
    defparam i5_3_lut_adj_1077.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1078 (.I0(n43050), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[12] [6]), .I3(n42977), .O(n15_adj_3305));   // verilog/coms.v(73[16:27])
    defparam i6_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1079 (.I0(n15_adj_3305), .I1(n42704), .I2(n14_adj_3304), 
            .I3(\data_out_frame[13] [0]), .O(n23267));   // verilog/coms.v(73[16:27])
    defparam i8_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1080 (.I0(\data_out_frame[17] [5]), .I1(n22926), 
            .I2(n22520), .I3(GND_net), .O(n23345));
    defparam i2_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i939_2_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1695));   // verilog/coms.v(69[16:27])
    defparam i939_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10152_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[0] ), .O(n23566));
    defparam i10152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10454_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[6]), 
            .I3(\data_in_frame[8]_c [6]), .O(n23868));
    defparam i10454_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10153_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [0]), 
            .I3(\Ki[0] ), .O(n23567));
    defparam i10153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10154_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [0]), 
            .I3(\Kd[0] ), .O(n23568));
    defparam i10154_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10455_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[5]), 
            .I3(\data_in_frame[8]_c [5]), .O(n23869));
    defparam i10455_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10155_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [0]), 
            .I3(gearBoxRatio[0]), .O(n23569));
    defparam i10155_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(n42480), .I1(n42806), .I2(GND_net), 
            .I3(GND_net), .O(n1444));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1082 (.I0(\data_out_frame[14] [5]), .I1(n42781), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[10] [1]), .O(n10_adj_3208));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1083 (.I0(\data_out_frame[10] [2]), .I1(n42434), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[8] [0]), .O(n10_adj_3160));   // verilog/coms.v(69[16:62])
    defparam i4_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1084 (.I0(n22445), .I1(n42480), .I2(\data_out_frame[14] [4]), 
            .I3(\data_out_frame[5][2] ), .O(n12_adj_3306));
    defparam i5_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1085 (.I0(\data_out_frame[12] [3]), .I1(n12_adj_3306), 
            .I2(n42809), .I3(\data_out_frame[12] [2]), .O(n38811));
    defparam i6_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(n38811), .I1(n39144), .I2(GND_net), 
            .I3(GND_net), .O(n22458));
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1087 (.I0(n1515), .I1(\data_out_frame[12] [5]), 
            .I2(n21999), .I3(n42822), .O(n10_adj_3307));
    defparam i4_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1088 (.I0(\data_out_frame[13] [0]), .I1(n22779), 
            .I2(n42992), .I3(n22458), .O(n20));   // verilog/coms.v(71[16:42])
    defparam i8_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1089 (.I0(\data_out_frame[14] [0]), .I1(n1695), 
            .I2(n42883), .I3(\data_out_frame[13] [2]), .O(n19_adj_3308));   // verilog/coms.v(71[16:42])
    defparam i7_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1090 (.I0(n38954), .I1(\data_out_frame[13] [3]), 
            .I2(n42598), .I3(\data_out_frame[13] [1]), .O(n21_adj_3309));   // verilog/coms.v(71[16:42])
    defparam i9_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut (.I0(n21_adj_3309), .I1(n19_adj_3308), .I2(n20), 
            .I3(GND_net), .O(n44021));   // verilog/coms.v(71[16:42])
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1091 (.I0(n44021), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[15] [0]), .I3(\data_out_frame[13] [5]), 
            .O(n18_adj_3310));
    defparam i7_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1092 (.I0(\data_out_frame[15] [4]), .I1(n18_adj_3310), 
            .I2(\data_out_frame[15] [1]), .I3(n42905), .O(n20_adj_3311));
    defparam i9_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut (.I0(n42846), .I1(\data_out_frame[15] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3312));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1093 (.I0(n15_adj_3312), .I1(n20_adj_3311), .I2(\data_out_frame[15] [2]), 
            .I3(n39144), .O(n39125));
    defparam i10_4_lut_adj_1093.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(n38601), .I1(n43500), .I2(GND_net), 
            .I3(GND_net), .O(n42751));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n22674));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1096 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42694));
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1097 (.I0(n22793), .I1(n42694), .I2(\data_out_frame[16] [4]), 
            .I3(GND_net), .O(n42944));
    defparam i2_3_lut_adj_1097.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22668));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[2]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[3]), 
            .O(n35));   // verilog/coms.v(100[12:33])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'haa80;
    SB_LUT4 i4_4_lut_adj_1099 (.I0(n23251), .I1(n39125), .I2(n23136), 
            .I3(n6_adj_3313), .O(n43500));
    defparam i4_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1100 (.I0(n23247), .I1(n22674), .I2(\data_out_frame[20] [0]), 
            .I3(n42751), .O(n12_adj_3314));
    defparam i5_4_lut_adj_1100.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1101 (.I0(n23345), .I1(n12_adj_3314), .I2(n23267), 
            .I3(n43803), .O(n42533));
    defparam i6_4_lut_adj_1101.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1102 (.I0(\data_out_frame[20] [1]), .I1(n42533), 
            .I2(n39189), .I3(GND_net), .O(n43873));
    defparam i2_3_lut_adj_1102.LUT_INIT = 16'h9696;
    SB_LUT4 i10158_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n23572));
    defparam i10158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1103 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n23004));
    defparam i2_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1104 (.I0(n23004), .I1(n42977), .I2(n42938), 
            .I3(\data_out_frame[8] [5]), .O(n1595));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1105 (.I0(\data_out_frame[15] [3]), .I1(n42669), 
            .I2(n1595), .I3(\data_out_frame[13] [1]), .O(n22520));   // verilog/coms.v(71[16:42])
    defparam i3_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1106 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[17] [5]), .I3(GND_net), .O(n42584));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1106.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(n22520), .I1(n43023), .I2(GND_net), 
            .I3(GND_net), .O(n42876));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42542));
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1109 (.I0(n38601), .I1(n42876), .I2(n42584), 
            .I3(\data_out_frame[19] [7]), .O(n39189));
    defparam i3_4_lut_adj_1109.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1110 (.I0(\data_out_frame[9] [0]), .I1(n42450), 
            .I2(n22937), .I3(GND_net), .O(n1506));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1110.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n22482));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1112 (.I0(n42770), .I1(\data_out_frame[17] [6]), 
            .I2(n22482), .I3(n22843), .O(n18_adj_3315));
    defparam i7_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1113 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3316));
    defparam i5_2_lut_adj_1113.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1114 (.I0(n22926), .I1(n18_adj_3315), .I2(\data_out_frame[18] [0]), 
            .I3(\data_out_frame[13] [5]), .O(n20_adj_3317));
    defparam i9_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1115 (.I0(n42935), .I1(n20_adj_3317), .I2(n16_adj_3316), 
            .I3(n42453), .O(n43023));
    defparam i10_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1116 (.I0(n42917), .I1(n43023), .I2(n42672), 
            .I3(GND_net), .O(n22017));
    defparam i2_3_lut_adj_1116.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1117 (.I0(n22017), .I1(\data_out_frame[20] [2]), 
            .I2(n38668), .I3(GND_net), .O(n43657));
    defparam i2_3_lut_adj_1117.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1118 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(n23274), .I3(n42711), .O(n10_adj_3318));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1119 (.I0(\data_out_frame[11] [1]), .I1(n10_adj_3318), 
            .I2(\data_out_frame[11] [2]), .I3(GND_net), .O(n1509));   // verilog/coms.v(73[16:27])
    defparam i5_3_lut_adj_1119.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42453));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_out_frame[13] [3]), .I1(n1509), 
            .I2(GND_net), .I3(GND_net), .O(n42659));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1122 (.I0(\data_out_frame[15] [5]), .I1(n42659), 
            .I2(n42453), .I3(n38210), .O(n38601));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_out_frame[18] [1]), .I1(n38601), 
            .I2(GND_net), .I3(GND_net), .O(n43065));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1124 (.I0(n42642), .I1(n43065), .I2(\data_out_frame[20] [3]), 
            .I3(GND_net), .O(n42761));
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1125 (.I0(n42761), .I1(n43020), .I2(\data_out_frame[16] [1]), 
            .I3(GND_net), .O(n38668));
    defparam i2_3_lut_adj_1125.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_out_frame[5] [0]), .I1(n42700), 
            .I2(GND_net), .I3(GND_net), .O(n42935));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1127 (.I0(n22853), .I1(n42935), .I2(\data_out_frame[8] [6]), 
            .I3(n23111), .O(n38210));
    defparam i3_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1128 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n43050));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3319));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_LUT4 i10159_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [0]), 
            .I3(PWMLimit[0]), .O(n23573));
    defparam i10159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1130 (.I0(n23194), .I1(\data_out_frame[6] [1]), 
            .I2(n42646), .I3(n6_adj_3319), .O(n42806));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i10171_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [0]), 
            .I3(deadband[0]), .O(n23585));
    defparam i10171_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33576_2_lut_3_lut_4_lut (.I0(n20088), .I1(n22289), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(\FRAME_MATCHER.state [0]), .O(n43084));
    defparam i33576_2_lut_3_lut_4_lut.LUT_INIT = 16'h5557;
    SB_LUT4 i2_3_lut_adj_1131 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n22937));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1131.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42704));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1133 (.I0(\data_out_frame[6] [3]), .I1(n22937), 
            .I2(GND_net), .I3(GND_net), .O(n42711));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1134 (.I0(\data_out_frame[10] [4]), .I1(n42646), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n42471));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_adj_1134.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1135 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[7] [7]), .O(n42434));
    defparam i3_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1136 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n42477));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1137 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[11] [2]), .I3(\data_out_frame[6] [4]), .O(n42700));
    defparam i3_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1138 (.I0(\data_out_frame[10] [2]), .I1(n42434), 
            .I2(\data_out_frame[7] [5]), .I3(\data_out_frame[12] [3]), .O(n42781));   // verilog/coms.v(71[16:34])
    defparam i3_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1139 (.I0(\data_out_frame[6] [6]), .I1(n43050), 
            .I2(\data_out_frame[11] [0]), .I3(\data_out_frame[11] [1]), 
            .O(n42450));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1140 (.I0(n42450), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[12] [5]), .I3(n18_adj_3320), .O(n30_adj_3321));   // verilog/coms.v(73[16:27])
    defparam i13_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1141 (.I0(n42498), .I1(\data_out_frame[11] [3]), 
            .I2(n22445), .I3(n42986), .O(n28_adj_3322));   // verilog/coms.v(73[16:27])
    defparam i11_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1142 (.I0(n42781), .I1(n42539), .I2(n42700), 
            .I3(n42477), .O(n29_adj_3323));   // verilog/coms.v(73[16:27])
    defparam i12_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1143 (.I0(n42938), .I1(n43053), .I2(n42471), 
            .I3(n42711), .O(n27_adj_3324));   // verilog/coms.v(73[16:27])
    defparam i10_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1144 (.I0(n27_adj_3324), .I1(n29_adj_3323), .I2(n28_adj_3322), 
            .I3(n30_adj_3321), .O(n38954));   // verilog/coms.v(73[16:27])
    defparam i16_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1145 (.I0(n22289), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n22296));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_3_lut_adj_1145.LUT_INIT = 16'hefef;
    SB_LUT4 i97_2_lut_3_lut (.I0(n22422), .I1(n3761), .I2(n20088), .I3(GND_net), 
            .O(n53));   // verilog/coms.v(113[11:12])
    defparam i97_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1146 (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n22421), .I3(GND_net), .O(n22422));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_3_lut_adj_1146.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_3_lut_4_lut_adj_1147 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n20088), 
            .I2(n2103), .I3(n53), .O(n41720));
    defparam i1_3_lut_4_lut_adj_1147.LUT_INIT = 16'haa80;
    SB_LUT4 i8_4_lut_adj_1148 (.I0(\data_out_frame[11] [5]), .I1(n42549), 
            .I2(n42992), .I3(\data_out_frame[7] [3]), .O(n20_adj_3325));
    defparam i8_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1149 (.I0(\data_out_frame[18] [2]), .I1(n42846), 
            .I2(\data_out_frame[7] [4]), .I3(\data_out_frame[11] [6]), .O(n19_adj_3326));
    defparam i7_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1150 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [3]), .I3(n42550), .O(n21_adj_3327));
    defparam i9_4_lut_adj_1150.LUT_INIT = 16'h9669;
    SB_LUT4 i11_3_lut_adj_1151 (.I0(n21_adj_3327), .I1(n19_adj_3326), .I2(n20_adj_3325), 
            .I3(GND_net), .O(n42913));
    defparam i11_3_lut_adj_1151.LUT_INIT = 16'h9696;
    SB_LUT4 i10690_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [3]), 
            .I3(gearBoxRatio[19]), .O(n24104));
    defparam i10690_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1152 (.I0(n21986), .I1(n42641), .I2(GND_net), 
            .I3(GND_net), .O(n39149));
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22793));
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1154 (.I0(\data_out_frame[20] [4]), .I1(n42965), 
            .I2(n42672), .I3(n22793), .O(n10_adj_3328));
    defparam i4_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1155 (.I0(n42913), .I1(n10_adj_3328), .I2(\data_out_frame[16] [2]), 
            .I3(GND_net), .O(n42463));
    defparam i5_3_lut_adj_1155.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1156 (.I0(n39102), .I1(n42463), .I2(\data_out_frame[20] [5]), 
            .I3(GND_net), .O(n43836));
    defparam i2_3_lut_adj_1156.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22853));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42539));
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23274));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23111));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1161 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42655));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1161.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1162 (.I0(\data_out_frame[11] [4]), .I1(n42655), 
            .I2(n23111), .I3(n23274), .O(n42905));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i33573_2_lut_3_lut (.I0(n5019), .I1(n3346), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(GND_net), .O(n23438));
    defparam i33573_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_out_frame[13] [7]), .I1(n42971), 
            .I2(GND_net), .I3(GND_net), .O(n38948));
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1164 (.I0(\data_out_frame[18] [4]), .I1(n23271), 
            .I2(n42965), .I3(\data_out_frame[16] [3]), .O(n39102));
    defparam i2_3_lut_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1165 (.I0(n1515), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[15] [7]), .I3(n38948), .O(n42641));
    defparam i3_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_out_frame[14] [0]), .I1(n42641), 
            .I2(GND_net), .I3(GND_net), .O(n42642));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1167 (.I0(n42837), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[11] [5]), .I3(n42989), .O(n10_adj_3329));
    defparam i4_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1168 (.I0(n21999), .I1(n23114), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_3330));
    defparam i2_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1169 (.I0(n7_adj_3330), .I1(\data_out_frame[16] [1]), 
            .I2(n42642), .I3(\data_out_frame[18] [3]), .O(n42965));
    defparam i4_4_lut_adj_1169.LUT_INIT = 16'h9669;
    SB_LUT4 i10456_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[4]), 
            .I3(\data_in_frame[8]_c [4]), .O(n23870));
    defparam i10456_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_out_frame[18] [4]), .I1(n23271), 
            .I2(GND_net), .I3(GND_net), .O(n42764));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1171 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22843));
    defparam i1_2_lut_adj_1171.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42501));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42989));
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42774));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1175 (.I0(n42989), .I1(\data_out_frame[7] [0]), 
            .I2(n42501), .I3(n22843), .O(n14_adj_3331));
    defparam i6_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1176 (.I0(\data_out_frame[11] [6]), .I1(n14_adj_3331), 
            .I2(n10_adj_3332), .I3(\data_out_frame[5][2] ), .O(n42971));
    defparam i7_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1177 (.I0(n23114), .I1(n23251), .I2(n23271), 
            .I3(GND_net), .O(n42883));
    defparam i1_2_lut_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1178 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[10] [0]), .I3(\data_out_frame[9] [7]), .O(n42809));
    defparam i1_2_lut_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i10691_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [2]), 
            .I3(gearBoxRatio[18]), .O(n24105));
    defparam i10691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[5][2] ), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42837));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n42430));
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_out_frame[11] [5]), .I1(n42430), 
            .I2(GND_net), .I3(GND_net), .O(n42968));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i10692_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [1]), 
            .I3(gearBoxRatio[17]), .O(n24106));
    defparam i10692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1182 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[12] [2]), .I3(n6_adj_3333), .O(n42498));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23194));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 i10693_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [0]), 
            .I3(gearBoxRatio[16]), .O(n24107));
    defparam i10693_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1184 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n43053));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1184.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42778));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42825));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42770));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42986));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42605));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i10710_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [6]), 
            .I3(\Kd[6] ), .O(n24124));
    defparam i10710_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1190 (.I0(n42809), .I1(n42825), .I2(\data_out_frame[14] [2]), 
            .I3(n42778), .O(n12_adj_3334));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1191 (.I0(n42605), .I1(n12_adj_3334), .I2(n42986), 
            .I3(n42770), .O(n23271));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1192 (.I0(n23194), .I1(n42498), .I2(\data_out_frame[14] [3]), 
            .I3(\data_out_frame[5] [6]), .O(n12_adj_3335));   // verilog/coms.v(72[16:27])
    defparam i5_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1193 (.I0(\data_out_frame[9] [7]), .I1(n12_adj_3335), 
            .I2(n42822), .I3(\data_out_frame[9] [6]), .O(n23251));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1194 (.I0(n23251), .I1(n23271), .I2(GND_net), 
            .I3(GND_net), .O(n1716));
    defparam i1_2_lut_adj_1194.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1195 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[14] [1]), .O(n18_adj_3336));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1196 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3337));   // verilog/coms.v(71[16:27])
    defparam i5_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i10711_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [5]), 
            .I3(\Kd[5] ), .O(n24125));
    defparam i10711_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1197 (.I0(\data_out_frame[13] [7]), .I1(n18_adj_3336), 
            .I2(\data_out_frame[9] [6]), .I3(n42968), .O(n20_adj_3338));   // verilog/coms.v(71[16:27])
    defparam i9_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1198 (.I0(n42774), .I1(n20_adj_3338), .I2(n16_adj_3337), 
            .I3(\data_out_frame[7] [5]), .O(n23114));   // verilog/coms.v(71[16:27])
    defparam i10_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(n21986), .I1(\data_out_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3339));
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1200 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[18] [4]), .I3(n6_adj_3339), .O(n42691));
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1201 (.I0(n42691), .I1(n42883), .I2(\data_out_frame[18] [5]), 
            .I3(GND_net), .O(n22019));
    defparam i2_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42720));
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1203 (.I0(n39102), .I1(n42720), .I2(n22019), 
            .I3(GND_net), .O(n43887));
    defparam i2_3_lut_adj_1203.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1204 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[12] [1]), .I3(GND_net), .O(n6_adj_3333));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1204.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1205 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[5][2] ), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n42822));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1205.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(n22421), .I1(n42390), .I2(GND_net), 
            .I3(GND_net), .O(n3_adj_3340));
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1207 (.I0(\FRAME_MATCHER.state_c [3]), .I1(n37), 
            .I2(n61), .I3(n3_adj_3340), .O(n11));
    defparam i1_4_lut_adj_1207.LUT_INIT = 16'haaa8;
    SB_LUT4 i10712_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [4]), 
            .I3(\Kd[4] ), .O(n24126));
    defparam i10712_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1208 (.I0(n22297), .I1(n11), .I2(n22421), .I3(\FRAME_MATCHER.state_31__N_1925 [3]), 
            .O(n41950));
    defparam i1_4_lut_adj_1208.LUT_INIT = 16'hcdcc;
    SB_LUT4 i10457_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[3]), 
            .I3(\data_in_frame[8]_c [3]), .O(n23871));
    defparam i10457_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41722));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1210 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42385));
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n7_adj_3342), 
            .I2(GND_net), .I3(GND_net), .O(n41796));
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42389));
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n7_adj_3342), 
            .I2(GND_net), .I3(GND_net), .O(n41794));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42381));
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1215 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n7_adj_3342), 
            .I2(GND_net), .I3(GND_net), .O(n41792));
    defparam i1_2_lut_adj_1215.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42379));
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n10_adj_3332));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15036_2_lut (.I0(\FRAME_MATCHER.state_c [8]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n28428));
    defparam i15036_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_4_lut_adj_1217 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[11] [4]), 
            .I2(n10_adj_3329), .I3(n22853), .O(n21999));
    defparam i5_3_lut_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42374));
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1219 (.I0(n21999), .I1(n21986), .I2(n42641), 
            .I3(GND_net), .O(n42672));
    defparam i1_2_lut_3_lut_adj_1219.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42382));
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41724));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42387));
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\FRAME_MATCHER.state_c [12]), .I1(n7_adj_3342), 
            .I2(GND_net), .I3(GND_net), .O(n41790));
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h8888;
    SB_LUT4 i10458_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[2]), 
            .I3(\data_in_frame[8][2] ), .O(n23872));
    defparam i10458_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10713_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [3]), 
            .I3(\Kd[3] ), .O(n24127));
    defparam i10713_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\FRAME_MATCHER.state_c [12]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42383));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1225 (.I0(n38210), .I1(n22077), .I2(n38954), 
            .I3(\data_out_frame[12] [5]), .O(n42550));
    defparam i1_2_lut_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i15037_2_lut (.I0(\FRAME_MATCHER.state_c [13]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n28430));
    defparam i15037_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1226 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n18_adj_3320));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1226.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1227 (.I0(n32579), .I1(\FRAME_MATCHER.state_c [14]), 
            .I2(GND_net), .I3(GND_net), .O(n28432));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_adj_1227.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1228 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[5] [5]), .O(n22445));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i10714_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [2]), 
            .I3(\Kd[2] ), .O(n24128));
    defparam i10714_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i70_2_lut (.I0(n32579), .I1(\FRAME_MATCHER.state_c [15]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_3158));
    defparam i70_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1229 (.I0(n61), .I1(n1_adj_3128), .I2(n22289), 
            .I3(n42371), .O(n7_adj_3342));
    defparam i2_4_lut_adj_1229.LUT_INIT = 16'hefee;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n7_adj_3342), 
            .I2(GND_net), .I3(GND_net), .O(n41788));
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42386));
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1232 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[10] [7]), .I3(GND_net), .O(n42938));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1233 (.I0(\FRAME_MATCHER.state_c [17]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3157));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_adj_1233.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1234 (.I0(n42761), .I1(n43020), .I2(\data_out_frame[16] [1]), 
            .I3(n42463), .O(n42464));
    defparam i1_2_lut_4_lut_adj_1234.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1235 (.I0(\FRAME_MATCHER.state_c [18]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3156));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h8888;
    SB_LUT4 i10715_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [1]), 
            .I3(\Kd[1] ), .O(n24129));
    defparam i10715_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41730));
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1237 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42378));
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41784));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1239 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42380));
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h8888;
    SB_LUT4 i10716_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [7]), 
            .I3(\Ki[7] ), .O(n24130));
    defparam i10716_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10459_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[1]), 
            .I3(\data_in_frame[8]_c [1]), .O(n23873));
    defparam i10459_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(n21986), .I1(n42641), .I2(n42913), 
            .I3(GND_net), .O(n43020));
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'h6969;
    SB_LUT4 i74_2_lut (.I0(n32579), .I1(\FRAME_MATCHER.state_c [21]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_3155));
    defparam i74_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\FRAME_MATCHER.state_c [22]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41782));
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h8888;
    SB_LUT4 i10717_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [6]), 
            .I3(\Ki[6] ), .O(n24131));
    defparam i10717_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\FRAME_MATCHER.state_c [22]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42388));
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1243 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(n38601), .I3(GND_net), .O(n42917));
    defparam i1_2_lut_3_lut_adj_1243.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3154));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\FRAME_MATCHER.state_c [24]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41728));
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h8888;
    SB_LUT4 i10694_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [7]), 
            .I3(gearBoxRatio[15]), .O(n24108));
    defparam i10694_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10695_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [6]), 
            .I3(gearBoxRatio[14]), .O(n24109));
    defparam i10695_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\FRAME_MATCHER.state_c [24]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42384));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h8888;
    SB_LUT4 i10718_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [5]), 
            .I3(\Ki[5] ), .O(n24132));
    defparam i10718_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\FRAME_MATCHER.state_c [25]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41726));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\FRAME_MATCHER.state_c [25]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42376));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1249 (.I0(\data_out_frame[13] [3]), .I1(n1509), 
            .I2(n42669), .I3(\data_out_frame[15] [4]), .O(n22926));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\FRAME_MATCHER.state_c [26]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3153));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h8888;
    SB_LUT4 i10460_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42411), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n23874));
    defparam i10460_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1251 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(n42450), .I3(n22937), .O(n42669));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\FRAME_MATCHER.state_c [27]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3152));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h8888;
    SB_LUT4 i10319_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [7]), 
            .I3(PWMLimit[23]), .O(n23733));
    defparam i10319_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1253 (.I0(n39189), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(n22017), .O(n43874));
    defparam i2_3_lut_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i10320_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [6]), 
            .I3(PWMLimit[22]), .O(n23734));
    defparam i10320_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\FRAME_MATCHER.state_c [28]), .I1(n32579), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3151));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\FRAME_MATCHER.state_c [29]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41732));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\FRAME_MATCHER.state_c [29]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42375));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1257 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[11] [0]), .I3(\data_out_frame[10] [5]), 
            .O(n42977));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1258 (.I0(\data_out_frame[16] [7]), .I1(n22793), 
            .I2(n42694), .I3(\data_out_frame[16] [4]), .O(n6_adj_3313));
    defparam i1_2_lut_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i14974_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [5]), 
            .I3(PWMLimit[21]), .O(n28366));
    defparam i14974_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1259 (.I0(n22421), .I1(n42390), .I2(n22294), 
            .I3(n20078), .O(n42373));
    defparam i1_4_lut_adj_1259.LUT_INIT = 16'h4544;
    SB_LUT4 i1_2_lut_3_lut_adj_1260 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[17] [2]), .I3(GND_net), .O(n23247));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1260.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1261 (.I0(\data_out_frame[11] [5]), .I1(n42430), 
            .I2(n10_adj_3307), .I3(n42778), .O(n42598));
    defparam i5_3_lut_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1262 (.I0(n1_adj_3128), .I1(n22289), .I2(n7_c), 
            .I3(n42371), .O(n12_adj_3341));
    defparam i1_4_lut_adj_1262.LUT_INIT = 16'hbbba;
    SB_LUT4 i14941_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [4]), 
            .I3(PWMLimit[20]), .O(n28334));
    defparam i14941_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n12_adj_3341), 
            .I2(GND_net), .I3(GND_net), .O(n41780));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n42373), 
            .I2(GND_net), .I3(GND_net), .O(n42377));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1265 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n42480), .I3(n42806), .O(n22779));
    defparam i1_2_lut_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1266 (.I0(\data_out_frame[12] [4]), .I1(n42480), 
            .I2(n42806), .I3(GND_net), .O(n42688));
    defparam i1_2_lut_3_lut_adj_1266.LUT_INIT = 16'h9696;
    SB_LUT4 i15183_4_lut (.I0(n10_adj_3253), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n22342), .O(n3761));   // verilog/coms.v(249[9:58])
    defparam i15183_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(n3761), .I1(n20088), .I2(GND_net), 
            .I3(GND_net), .O(n20078));   // verilog/coms.v(249[6] 251[9])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1268 (.I0(n30621), .I1(n5_adj_3343), .I2(n35), 
            .I3(byte_transmit_counter[7]), .O(n89));   // verilog/coms.v(100[12:33])
    defparam i1_4_lut_adj_1268.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_3_lut_adj_1269 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(n38353), .I3(GND_net), .O(n42902));
    defparam i1_2_lut_3_lut_adj_1269.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1270 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [6]), 
            .I2(n10_adj_3291), .I3(\data_out_frame[15] [1]), .O(n38351));
    defparam i5_3_lut_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1271 (.I0(\data_out_frame[19] [3]), .I1(n38351), 
            .I2(n23295), .I3(n42491), .O(n42492));
    defparam i1_2_lut_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1272 (.I0(\FRAME_MATCHER.state[2] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n22297));   // verilog/coms.v(161[5:29])
    defparam i1_2_lut_adj_1272.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1273 (.I0(\data_out_frame[20] [6]), .I1(n38811), 
            .I2(\data_out_frame[16] [3]), .I3(\data_out_frame[16] [5]), 
            .O(n6_adj_3288));
    defparam i1_2_lut_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1274 (.I0(\FRAME_MATCHER.state_c [1]), .I1(n28987), 
            .I2(\FRAME_MATCHER.state_c [3]), .I3(n22297), .O(n22309));   // verilog/coms.v(195[5:24])
    defparam i3_4_lut_adj_1274.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_1275 (.I0(n22289), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n22299));   // verilog/coms.v(148[5:9])
    defparam i1_2_lut_3_lut_adj_1275.LUT_INIT = 16'hfefe;
    SB_LUT4 i10323_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [3]), 
            .I3(PWMLimit[19]), .O(n23737));
    defparam i10323_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_adj_1276 (.I0(n63_adj_3266), .I1(n28564), .I2(n22424), 
            .I3(GND_net), .O(n8_adj_3344));
    defparam i3_3_lut_adj_1276.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut_adj_1277 (.I0(n22309), .I1(n8_adj_3344), .I2(n22421), 
            .I3(\FRAME_MATCHER.state [0]), .O(n2103));
    defparam i4_4_lut_adj_1277.LUT_INIT = 16'h8880;
    SB_LUT4 i6_4_lut_adj_1278 (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [27]), .I3(\FRAME_MATCHER.i [10]), .O(n14_adj_3345));
    defparam i6_4_lut_adj_1278.LUT_INIT = 16'hfffe;
    SB_LUT4 i10324_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [2]), 
            .I3(PWMLimit[18]), .O(n23738));
    defparam i10324_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1279 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [28]), 
            .I2(\FRAME_MATCHER.i [25]), .I3(\FRAME_MATCHER.i [11]), .O(n13_adj_3346));
    defparam i5_4_lut_adj_1279.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1280 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [13]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3347));
    defparam i2_2_lut_adj_1280.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1281 (.I0(\FRAME_MATCHER.i [18]), .I1(n13_adj_3346), 
            .I2(n14_adj_3345), .I3(GND_net), .O(n19_adj_3348));
    defparam i1_3_lut_adj_1281.LUT_INIT = 16'hfefe;
    SB_LUT4 i14_4_lut_adj_1282 (.I0(\FRAME_MATCHER.i [19]), .I1(n19_adj_3348), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n20_adj_3347), .O(n32_adj_3349));
    defparam i14_4_lut_adj_1282.LUT_INIT = 16'hfffe;
    SB_LUT4 i10325_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [1]), 
            .I3(PWMLimit[17]), .O(n23739));
    defparam i10325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1283 (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [29]), .I3(\FRAME_MATCHER.i [20]), .O(n30_adj_3350));
    defparam i12_4_lut_adj_1283.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1284 (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [16]), .I3(\FRAME_MATCHER.i [23]), .O(n31_adj_3351));
    defparam i13_4_lut_adj_1284.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1285 (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [17]), 
            .I2(\FRAME_MATCHER.i [30]), .I3(\FRAME_MATCHER.i [14]), .O(n29_adj_3352));
    defparam i11_4_lut_adj_1285.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1286 (.I0(n29_adj_3352), .I1(n31_adj_3351), .I2(n30_adj_3350), 
            .I3(n32_adj_3349), .O(n22342));
    defparam i17_4_lut_adj_1286.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1287 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_3353));
    defparam i5_3_lut_adj_1287.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1288 (.I0(\data_in[0] [6]), .I1(n22408), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_3354));
    defparam i6_4_lut_adj_1288.LUT_INIT = 16'hfeff;
    SB_LUT4 i10326_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[5] [0]), 
            .I3(PWMLimit[16]), .O(n23740));
    defparam i10326_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1289 (.I0(n15_adj_3354), .I1(\data_in[2] [2]), 
            .I2(n14_adj_3353), .I3(\data_in[0] [3]), .O(n22195));
    defparam i8_4_lut_adj_1289.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_1290 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_3355));
    defparam i6_4_lut_adj_1290.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1291 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_3356));
    defparam i7_4_lut_adj_1291.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1292 (.I0(n17_adj_3356), .I1(\data_in[1] [6]), 
            .I2(n16_adj_3355), .I3(\data_in[3] [7]), .O(n22280));
    defparam i9_4_lut_adj_1292.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1293 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_3357));
    defparam i4_4_lut_adj_1293.LUT_INIT = 16'hfdff;
    SB_LUT4 i10327_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6] [7]), 
            .I3(PWMLimit[15]), .O(n23741));
    defparam i10327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1294 (.I0(\data_in[2] [7]), .I1(n10_adj_3357), 
            .I2(\data_in[3] [4]), .I3(GND_net), .O(n22408));
    defparam i5_3_lut_adj_1294.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1295 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_3358));
    defparam i6_4_lut_adj_1295.LUT_INIT = 16'hfeff;
    SB_LUT4 i14351_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6] [6]), 
            .I3(PWMLimit[14]), .O(n27746));
    defparam i14351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\data_in[3] [5]), .I1(\data_in[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1297 (.I0(n9), .I1(n14_adj_3358), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [1]), .O(n22316));
    defparam i7_4_lut_adj_1297.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1298 (.I0(\data_in[2] [4]), .I1(n22316), .I2(\data_in[1] [5]), 
            .I3(n22408), .O(n18_adj_3359));
    defparam i7_4_lut_adj_1298.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1299 (.I0(\data_in[0] [6]), .I1(n18_adj_3359), 
            .I2(\data_in[3] [0]), .I3(n22280), .O(n20_adj_3360));
    defparam i9_4_lut_adj_1299.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_1300 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3361));
    defparam i4_2_lut_adj_1300.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1301 (.I0(n15_adj_3361), .I1(n20_adj_3360), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_3143));
    defparam i10_4_lut_adj_1301.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1302 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n22195), .O(n16_adj_3362));
    defparam i6_4_lut_adj_1302.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1303 (.I0(n22280), .I1(\data_in[3] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[2] [3]), .O(n17_adj_3363));
    defparam i7_4_lut_adj_1303.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1304 (.I0(n17_adj_3363), .I1(\data_in[3] [1]), 
            .I2(n16_adj_3362), .I3(\data_in[3] [5]), .O(n63_c));
    defparam i9_4_lut_adj_1304.LUT_INIT = 16'hfbff;
    SB_LUT4 i8_4_lut_adj_1305 (.I0(n22316), .I1(\data_in[1] [3]), .I2(n22195), 
            .I3(\data_in[2] [0]), .O(n20_adj_3364));
    defparam i8_4_lut_adj_1305.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1306 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19_adj_3365));
    defparam i7_4_lut_adj_1306.LUT_INIT = 16'hfeff;
    SB_LUT4 i28808_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [5]), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [2]), .O(n44367));
    defparam i28808_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut_adj_1307 (.I0(n44367), .I1(n19_adj_3365), .I2(n20_adj_3364), 
            .I3(GND_net), .O(n63));
    defparam i11_3_lut_adj_1307.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(n22175), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3366));
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'heeee;
    SB_LUT4 i15177_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3366), .I3(\FRAME_MATCHER.i [1]), .O(n740));   // verilog/coms.v(157[9:60])
    defparam i15177_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1309 (.I0(n20088), .I1(n2103), .I2(GND_net), 
            .I3(GND_net), .O(n1_adj_3128));
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h8888;
    SB_LUT4 i72_2_lut (.I0(n32579), .I1(\FRAME_MATCHER.state_c [31]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_3149));
    defparam i72_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14297_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6] [5]), 
            .I3(PWMLimit[13]), .O(n27693));
    defparam i14297_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10330_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6] [4]), 
            .I3(PWMLimit[12]), .O(n23744));
    defparam i10330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10331_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6] [3]), 
            .I3(PWMLimit[11]), .O(n23745));
    defparam i10331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10332_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6] [2]), 
            .I3(PWMLimit[10]), .O(n23746));
    defparam i10332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10333_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6][1] ), 
            .I3(PWMLimit[9]), .O(n23747));
    defparam i10333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_302_Select_2_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state_31__N_1861[2] ), 
            .I1(n22294), .I2(n22421), .I3(n3761), .O(n7));
    defparam select_302_Select_2_i7_3_lut_4_lut.LUT_INIT = 16'h0302;
    SB_LUT4 i10334_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[6] [0]), 
            .I3(PWMLimit[8]), .O(n23748));
    defparam i10334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1310 (.I0(\FRAME_MATCHER.state[2] ), .I1(n63_adj_3143), 
            .I2(n63_c), .I3(n63), .O(\FRAME_MATCHER.state_31__N_1861[2] ));   // verilog/coms.v(143[7:84])
    defparam i1_2_lut_4_lut_adj_1310.LUT_INIT = 16'hb300;
    SB_LUT4 i1_2_lut_3_lut_adj_1311 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n28987), .I3(GND_net), .O(n4_adj_3284));
    defparam i1_2_lut_3_lut_adj_1311.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(n28404), .I1(n10_adj_3127), .I2(GND_net), 
            .I3(GND_net), .O(n42419));
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'hdddd;
    SB_LUT4 mux_550_i1_3_lut_4_lut (.I0(n31), .I1(n28411), .I2(tx_transmit_N_2648), 
            .I3(\FRAME_MATCHER.state [0]), .O(n28971));   // verilog/coms.v(147[4] 288[11])
    defparam mux_550_i1_3_lut_4_lut.LUT_INIT = 16'h0fee;
    SB_LUT4 i33581_4_lut_4_lut (.I0(n28987), .I1(\FRAME_MATCHER.state_c [3]), 
            .I2(\FRAME_MATCHER.state[2] ), .I3(n43205), .O(n42202));
    defparam i33581_4_lut_4_lut.LUT_INIT = 16'hefea;
    SB_LUT4 i13692_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [7]), 
            .I3(PWMLimit[7]), .O(n23749));
    defparam i13692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10336_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [6]), 
            .I3(PWMLimit[6]), .O(n23750));
    defparam i10336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13439_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [5]), 
            .I3(PWMLimit[5]), .O(n26838));
    defparam i13439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i27648_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [3]), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n43205));
    defparam i27648_2_lut_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i10338_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [4]), 
            .I3(PWMLimit[4]), .O(n23752));
    defparam i10338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10339_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [3]), 
            .I3(PWMLimit[3]), .O(n23753));
    defparam i10339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10340_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [2]), 
            .I3(PWMLimit[2]), .O(n23754));
    defparam i10340_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10341_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[7] [1]), 
            .I3(PWMLimit[1]), .O(n23755));
    defparam i10341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3146));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31511_2_lut (.I0(\data_out_frame[5] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46688));
    defparam i31511_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3145));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10342_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n23756));
    defparam i10342_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10343_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n23757));
    defparam i10343_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1313 (.I0(n38982), .I1(n42879), .I2(n42998), 
            .I3(GND_net), .O(n42753));
    defparam i1_2_lut_3_lut_adj_1313.LUT_INIT = 16'h9696;
    SB_LUT4 i10344_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n23758));
    defparam i10344_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10345_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode[4]), .O(n23759));
    defparam i10345_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1314 (.I0(\data_in_frame[20] [5]), .I1(\data_in_frame[18] [3]), 
            .I2(n39133), .I3(GND_net), .O(n6_adj_3258));
    defparam i1_2_lut_3_lut_adj_1314.LUT_INIT = 16'h9696;
    SB_LUT4 i10346_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n23760));
    defparam i10346_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10347_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n23761));
    defparam i10347_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1315 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[9] [6]), 
            .I2(n22777), .I3(GND_net), .O(n42926));
    defparam i1_2_lut_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1316 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[0] [7]), .O(n42663));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1317 (.I0(\data_in_frame[6] [7]), .I1(n22941), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n42980));
    defparam i1_2_lut_3_lut_adj_1317.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1318 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n42787));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_3_lut_adj_1318.LUT_INIT = 16'h9696;
    SB_LUT4 i10719_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [4]), 
            .I3(\Ki[4] ), .O(n24133));
    defparam i10719_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31871_2_lut (.I0(\data_out_frame[22] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46706));
    defparam i31871_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3130));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1319 (.I0(n22824), .I1(n42852), .I2(n23309), 
            .I3(\data_in_frame[9] [2]), .O(n42983));
    defparam i2_3_lut_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i10348_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n23762));
    defparam i10348_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10705_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [4]), 
            .I3(gearBoxRatio[4]), .O(n24119));
    defparam i10705_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut (.I0(n45), .I1(n3831), .I2(n2236[0]), .I3(byte_transmit_counter[0]), 
            .O(n24234));   // verilog/coms.v(110[11:16])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hec20;
    SB_LUT4 i10706_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [3]), 
            .I3(gearBoxRatio[3]), .O(n24120));
    defparam i10706_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10707_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [2]), 
            .I3(gearBoxRatio[2]), .O(n24121));
    defparam i10707_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29694_2_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n45253));
    defparam i29694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10245_2_lut_3_lut (.I0(n45), .I1(n3831), .I2(n23657), .I3(GND_net), 
            .O(n23659));   // verilog/coms.v(110[11:16])
    defparam i10245_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(r_SM_Main_2__N_2756[0]), .I1(tx_active), 
            .I2(GND_net), .I3(GND_net), .O(n30621));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3343));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'heeee;
    SB_LUT4 i33571_4_lut (.I0(n5_adj_3343), .I1(byte_transmit_counter[7]), 
            .I2(n30621), .I3(n35), .O(tx_transmit_N_2648));
    defparam i33571_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i10720_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [3]), 
            .I3(\Ki[3] ), .O(n24134));
    defparam i10720_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10721_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [2]), 
            .I3(\Ki[2] ), .O(n24135));
    defparam i10721_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10242_2_lut_3_lut (.I0(n45), .I1(n3831), .I2(n23654), .I3(GND_net), 
            .O(n23656));   // verilog/coms.v(110[11:16])
    defparam i10242_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i10722_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[3] [1]), 
            .I3(\Ki[1] ), .O(n24136));
    defparam i10722_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34266 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n49818));
    defparam byte_transmit_counter_0__bdd_4_lut_34266.LUT_INIT = 16'he4aa;
    SB_LUT4 i10723_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[7] ), .O(n24137));
    defparam i10723_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10724_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[6] ), .O(n24138));
    defparam i10724_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10725_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[5] ), .O(n24139));
    defparam i10725_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10726_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[4] ), .O(n24140));
    defparam i10726_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10727_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[3] ), .O(n24141));
    defparam i10727_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10239_2_lut_3_lut (.I0(n45), .I1(n3831), .I2(n23651), .I3(GND_net), 
            .O(n23653));   // verilog/coms.v(110[11:16])
    defparam i10239_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i73_2_lut_3_lut (.I0(n45), .I1(n3831), .I2(n19_adj_3122), 
            .I3(GND_net), .O(n23668));   // verilog/coms.v(110[11:16])
    defparam i73_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i10728_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[2] ), .O(n24142));
    defparam i10728_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10729_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[1] ), .O(n24143));
    defparam i10729_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10251_2_lut_3_lut (.I0(n45), .I1(n3831), .I2(n23663), .I3(GND_net), 
            .O(n23665));   // verilog/coms.v(110[11:16])
    defparam i10251_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i10730_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8]_c [7]), 
            .I3(IntegralLimit[23]), .O(n24144));
    defparam i10730_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10731_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8]_c [6]), 
            .I3(IntegralLimit[22]), .O(n24145));
    defparam i10731_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1322 (.I0(n45), .I1(n3831), .I2(n23660), 
            .I3(GND_net), .O(n23662));   // verilog/coms.v(110[11:16])
    defparam i1_2_lut_3_lut_adj_1322.LUT_INIT = 16'he0e0;
    SB_LUT4 i10732_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8]_c [5]), 
            .I3(IntegralLimit[21]), .O(n24146));
    defparam i10732_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10733_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8]_c [4]), 
            .I3(IntegralLimit[20]), .O(n24147));
    defparam i10733_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_1011_i15_2_lut_3_lut (.I0(n5_adj_3238), .I1(n23238), .I2(\data_in_frame[4] [6]), 
            .I3(GND_net), .O(n15));   // verilog/coms.v(230[9:81])
    defparam equal_1011_i15_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(\data_in_frame[11] [6]), .I1(n38403), 
            .I2(n42621), .I3(GND_net), .O(n42828));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'h9696;
    SB_LUT4 i10734_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8]_c [3]), 
            .I3(IntegralLimit[19]), .O(n24148));
    defparam i10734_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[15] [6]), .I3(GND_net), .O(n22560));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'h9696;
    SB_LUT4 i10735_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8][2] ), 
            .I3(IntegralLimit[18]), .O(n24149));
    defparam i10735_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10736_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8]_c [1]), 
            .I3(IntegralLimit[17]), .O(n24150));
    defparam i10736_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10737_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[8] [0]), 
            .I3(IntegralLimit[16]), .O(n24151));
    defparam i10737_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10696_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [5]), 
            .I3(gearBoxRatio[13]), .O(n24110));
    defparam i10696_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10689_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [4]), 
            .I3(gearBoxRatio[20]), .O(n24103));
    defparam i10689_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10688_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [5]), 
            .I3(gearBoxRatio[21]), .O(n24102));
    defparam i10688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10687_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [6]), 
            .I3(gearBoxRatio[22]), .O(n24101));
    defparam i10687_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1325 (.I0(n13), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[13] [1]), .I3(n42572), .O(n42575));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i10686_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[17] [7]), 
            .I3(gearBoxRatio[23]), .O(n24100));
    defparam i10686_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10868_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [7]), 
            .I3(deadband[23]), .O(n24282));
    defparam i10868_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10867_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [6]), 
            .I3(deadband[22]), .O(n24281));
    defparam i10867_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14973_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [5]), 
            .I3(deadband[21]), .O(n24280));
    defparam i14973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14942_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [4]), 
            .I3(deadband[20]), .O(n24279));
    defparam i14942_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10864_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [3]), 
            .I3(deadband[19]), .O(n24278));
    defparam i10864_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10863_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [2]), 
            .I3(deadband[18]), .O(n24277));
    defparam i10863_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10862_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [1]), 
            .I3(deadband[17]), .O(n24276));
    defparam i10862_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n49818_bdd_4_lut (.I0(n49818), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n49821));
    defparam n49818_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13438_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [5]), 
            .I3(deadband[5]), .O(n24264));
    defparam i13438_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10851_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [6]), 
            .I3(deadband[6]), .O(n24265));
    defparam i10851_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13691_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [7]), 
            .I3(deadband[7]), .O(n24266));
    defparam i13691_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10853_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12] [0]), 
            .I3(deadband[8]), .O(n24267));
    defparam i10853_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10854_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12][1] ), 
            .I3(deadband[9]), .O(n24268));
    defparam i10854_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10855_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12] [2]), 
            .I3(deadband[10]), .O(n24269));
    defparam i10855_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10856_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12] [3]), 
            .I3(deadband[11]), .O(n24270));
    defparam i10856_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10857_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12][4] ), 
            .I3(deadband[12]), .O(n24271));
    defparam i10857_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14299_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12] [5]), 
            .I3(deadband[13]), .O(n24272));
    defparam i14299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14350_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12] [6]), 
            .I3(deadband[14]), .O(n24273));
    defparam i14350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10860_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[12] [7]), 
            .I3(deadband[15]), .O(n24274));
    defparam i10860_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10861_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[11] [0]), 
            .I3(deadband[16]), .O(n24275));
    defparam i10861_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1326 (.I0(n22611), .I1(\data_in_frame[10] [7]), 
            .I2(n23007), .I3(\data_in_frame[12] [7]), .O(n23324));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1327 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[3] [6]), .O(Kp_23__N_379));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1328 (.I0(n22657), .I1(\data_in_frame[6] [2]), 
            .I2(n22538), .I3(GND_net), .O(n42608));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_3_lut_adj_1328.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1329 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[1] [7]), 
            .I2(n42443), .I3(\data_in_frame[4] [3]), .O(n23042));   // verilog/coms.v(230[9:81])
    defparam i2_3_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i10749_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [7]), 
            .I3(IntegralLimit[7]), .O(n24163));
    defparam i10749_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10750_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [6]), 
            .I3(IntegralLimit[6]), .O(n24164));
    defparam i10750_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10751_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [5]), 
            .I3(IntegralLimit[5]), .O(n24165));
    defparam i10751_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1330 (.I0(\data_in_frame[6] [0]), .I1(Kp_23__N_379), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n22908));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1330.LUT_INIT = 16'h9696;
    SB_LUT4 i10752_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [4]), 
            .I3(IntegralLimit[4]), .O(n24166));
    defparam i10752_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10753_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [3]), 
            .I3(IntegralLimit[3]), .O(n24167));
    defparam i10753_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10754_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [2]), 
            .I3(IntegralLimit[2]), .O(n24168));
    defparam i10754_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[13] [0]), .I3(GND_net), .O(n6_adj_3229));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1332 (.I0(Kp_23__N_459), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[7] [7]), .I3(\data_in_frame[8]_c [1]), .O(n43029));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1332.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1333 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[16] [2]), .I3(\data_in_frame[16] [6]), .O(n42457));
    defparam i2_3_lut_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1334 (.I0(n22698), .I1(n22960), .I2(n23105), 
            .I3(n42494), .O(n42819));
    defparam i2_3_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1335 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[14] [2]), .I3(n44074), .O(n42998));   // verilog/coms.v(83[17:70])
    defparam i2_3_lut_4_lut_adj_1335.LUT_INIT = 16'h9669;
    SB_LUT4 i15013_2_lut_2_lut_3_lut (.I0(n28564), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n28404));
    defparam i15013_2_lut_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i10755_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[10] [1]), 
            .I3(IntegralLimit[1]), .O(n24169));
    defparam i10755_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1336 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[15] [6]), .I3(\data_in_frame[15] [4]), .O(n42861));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_adj_1337 (.I0(\FRAME_MATCHER.state_c [3]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state [0]), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n4_c));
    defparam i1_4_lut_4_lut_adj_1337.LUT_INIT = 16'h0504;
    SB_LUT4 i6453_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [3]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n19790));
    defparam i6453_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i10845_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [1]), 
            .I3(deadband[1]), .O(n24259));
    defparam i10845_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1338 (.I0(\data_in_frame[17] [5]), .I1(n22611), 
            .I2(n42611), .I3(\data_in_frame[12] [7]), .O(n42995));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1339 (.I0(\data_in_frame[16] [0]), .I1(n22698), 
            .I2(Kp_23__N_866), .I3(n42494), .O(n23244));
    defparam i1_2_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[14] [4]), 
            .I2(n38879), .I3(GND_net), .O(n42831));
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1341 (.I0(n38429), .I1(n42666), .I2(n42910), 
            .I3(GND_net), .O(n42587));
    defparam i1_2_lut_3_lut_adj_1341.LUT_INIT = 16'h9696;
    SB_LUT4 i10847_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [2]), 
            .I3(deadband[2]), .O(n24261));
    defparam i10847_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1342 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [3]), 
            .I2(Kp_23__N_176), .I3(n38426), .O(n42524));
    defparam i2_3_lut_4_lut_adj_1342.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(\data_in_frame[18] [0]), .I1(n23105), 
            .I2(n38473), .I3(GND_net), .O(n42522));
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1344 (.I0(n12_adj_3216), .I1(n23013), .I2(n43673), 
            .I3(GND_net), .O(n43047));
    defparam i1_2_lut_4_lut_adj_1344.LUT_INIT = 16'h6969;
    SB_LUT4 i10848_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [3]), 
            .I3(deadband[3]), .O(n24262));
    defparam i10848_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10849_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[13] [4]), 
            .I3(deadband[4]), .O(n24263));
    defparam i10849_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10745_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [3]), 
            .I3(IntegralLimit[11]), .O(n24159));
    defparam i10745_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10746_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [2]), 
            .I3(IntegralLimit[10]), .O(n24160));
    defparam i10746_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10747_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [1]), 
            .I3(IntegralLimit[9]), .O(n24161));
    defparam i10747_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10748_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [0]), 
            .I3(IntegralLimit[8]), .O(n24162));
    defparam i10748_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10698_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [3]), 
            .I3(gearBoxRatio[11]), .O(n24112));
    defparam i10698_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10699_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [2]), 
            .I3(gearBoxRatio[10]), .O(n24113));
    defparam i10699_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10700_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [1]), 
            .I3(gearBoxRatio[9]), .O(n24114));
    defparam i10700_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10701_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [0]), 
            .I3(gearBoxRatio[8]), .O(n24115));
    defparam i10701_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1345 (.I0(\data_in_frame[12] [5]), .I1(n42799), 
            .I2(n43059), .I3(GND_net), .O(n6_adj_3212));
    defparam i1_2_lut_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1346 (.I0(\data_in_frame[15] [4]), .I1(n23064), 
            .I2(n22698), .I3(n42747), .O(n42953));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 select_267_Select_30_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_3163));
    defparam select_267_Select_30_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_31_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [31]), .O(n3));
    defparam select_267_Select_31_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_29_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_3165));
    defparam select_267_Select_29_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_28_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_3167));
    defparam select_267_Select_28_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n39117), .I3(GND_net), .O(n42460));
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_LUT4 select_267_Select_27_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_3169));
    defparam select_267_Select_27_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_26_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_3171));
    defparam select_267_Select_26_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i10702_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [7]), 
            .I3(gearBoxRatio[7]), .O(n24116));
    defparam i10702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10703_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [6]), 
            .I3(gearBoxRatio[6]), .O(n24117));
    defparam i10703_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_267_Select_25_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_3173));
    defparam select_267_Select_25_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_24_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_3175));
    defparam select_267_Select_24_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_23_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_3177));
    defparam select_267_Select_23_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i10704_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [5]), 
            .I3(gearBoxRatio[5]), .O(n24118));
    defparam i10704_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_267_Select_22_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_3179));
    defparam select_267_Select_22_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_21_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_3181));
    defparam select_267_Select_21_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i10741_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [7]), 
            .I3(IntegralLimit[15]), .O(n24155));
    defparam i10741_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_267_Select_20_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_3183));
    defparam select_267_Select_20_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_19_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_3185));
    defparam select_267_Select_19_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i10742_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [6]), 
            .I3(IntegralLimit[14]), .O(n24156));
    defparam i10742_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_267_Select_18_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_3187));
    defparam select_267_Select_18_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_17_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_3188));
    defparam select_267_Select_17_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i10743_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [5]), 
            .I3(IntegralLimit[13]), .O(n24157));
    defparam i10743_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10744_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[9] [4]), 
            .I3(IntegralLimit[12]), .O(n24158));
    defparam i10744_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10697_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[18] [4]), 
            .I3(gearBoxRatio[12]), .O(n24111));
    defparam i10697_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10708_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[19] [1]), 
            .I3(gearBoxRatio[1]), .O(n24122));
    defparam i10708_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10709_3_lut_4_lut (.I0(n28433), .I1(n63_adj_3266), .I2(\data_in_frame[4] [7]), 
            .I3(\Kd[7] ), .O(n24123));
    defparam i10709_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n44414), .I3(n44413), .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n44411), .I3(n44410), .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 select_267_Select_16_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_3189));
    defparam select_267_Select_16_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_15_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_3190));
    defparam select_267_Select_15_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_14_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_3191));
    defparam select_267_Select_14_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n44408), .I3(n44407), .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 select_267_Select_13_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_3192));
    defparam select_267_Select_13_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_12_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_3193));
    defparam select_267_Select_12_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n44399), .I3(n44398), .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 select_267_Select_11_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_3194));
    defparam select_267_Select_11_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_10_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_3195));
    defparam select_267_Select_10_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n44390), .I3(n44389), .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 select_267_Select_9_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_3196));
    defparam select_267_Select_9_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_8_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_3198));
    defparam select_267_Select_8_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n44393), .I3(n44392), .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 select_267_Select_7_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_3200));
    defparam select_267_Select_7_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_6_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_3202));
    defparam select_267_Select_6_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_5_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_3203));
    defparam select_267_Select_5_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n44396), .I3(n44395), .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 select_267_Select_4_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_3204));
    defparam select_267_Select_4_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_3_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_3205));
    defparam select_267_Select_3_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [2]), 
            .I2(n22824), .I3(GND_net), .O(n22777));
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'h9696;
    SB_LUT4 select_267_Select_2_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_3206));
    defparam select_267_Select_2_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_1_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_3207));
    defparam select_267_Select_1_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_267_Select_0_i3_2_lut_3_lut_4_lut (.I0(n28564), .I1(n22289), 
            .I2(n22297), .I3(\FRAME_MATCHER.i [0]), .O(n3_adj_3220));
    defparam select_267_Select_0_i3_2_lut_3_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1349 (.I0(\data_out_frame[16] [6]), .I1(n38811), 
            .I2(n39144), .I3(\data_out_frame[17] [0]), .O(n23136));
    defparam i1_2_lut_3_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1350 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [2]), 
            .I2(\data_in_frame[9] [4]), .I3(n42852), .O(n43002));
    defparam i2_3_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1351 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [0]), 
            .I2(n20914), .I3(n42899), .O(n22837));
    defparam i2_3_lut_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1352 (.I0(\data_out_frame[16] [6]), .I1(n38811), 
            .I2(n39144), .I3(\data_out_frame[18] [6]), .O(n6_adj_3290));
    defparam i1_2_lut_3_lut_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1353 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [0]), 
            .I2(n10_adj_3243), .I3(\data_in_frame[0] [4]), .O(n22824));
    defparam i5_3_lut_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n18_adj_3239));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1355 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[5] [3]), .I3(n22837), .O(n38403));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1356 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[3] [5]), .O(Kp_23__N_459));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1357 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[17] [3]), 
            .I2(n22668), .I3(n21999), .O(n43026));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1358 (.I0(n42430), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(n42905), .O(n1515));
    defparam i1_2_lut_3_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [4]), 
            .I2(n42971), .I3(GND_net), .O(n42992));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1359 (.I0(n740), .I1(n20088), .I2(n22289), 
            .I3(n22294), .O(n37));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_3_lut_4_lut_adj_1359.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1360 (.I0(n740), .I1(n20088), .I2(\FRAME_MATCHER.state[2] ), 
            .I3(\FRAME_MATCHER.state [0]), .O(n42371));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_3_lut_4_lut_adj_1360.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(n42663), .I3(GND_net), .O(n42508));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[9] [5]), 
            .I2(n43005), .I3(n42828), .O(n8_adj_3215));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n42505));
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(n22554), .I1(\data_in_frame[8]_c [5]), 
            .I2(\data_in_frame[10] [6]), .I3(GND_net), .O(n6_adj_3230));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(n22554), .I1(\data_in_frame[8]_c [5]), 
            .I2(n23042), .I3(n22954), .O(n23007));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i10157_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n23571));
    defparam i10157_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10517_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n23931));
    defparam i10517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10518_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n23932));
    defparam i10518_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10519_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n23933));
    defparam i10519_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10520_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n23934));
    defparam i10520_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10521_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n23935));
    defparam i10521_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10522_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n23936));
    defparam i10522_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10523_3_lut_4_lut (.I0(n8_adj_3126), .I1(n42403), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n23937));
    defparam i10523_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_2_lut_3_lut (.I0(n22538), .I1(Kp_23__N_459), .I2(\data_in_frame[5] [6]), 
            .I3(GND_net), .O(n18));   // verilog/coms.v(230[9:81])
    defparam i6_2_lut_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1365 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n42399), .I3(\FRAME_MATCHER.i [3]), .O(n42400));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1365.LUT_INIT = 16'hfeff;
    SB_LUT4 i27650_4_lut_4_lut (.I0(\FRAME_MATCHER.state_c [3]), .I1(\FRAME_MATCHER.state[2] ), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(\FRAME_MATCHER.state [0]), 
            .O(n43207));
    defparam i27650_4_lut_4_lut.LUT_INIT = 16'h4046;
    SB_LUT4 equal_67_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10));   // verilog/coms.v(154[7:23])
    defparam equal_67_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1366 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n28404), .I3(\FRAME_MATCHER.i [3]), .O(n42411));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1366.LUT_INIT = 16'hefff;
    SB_LUT4 equal_59_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3126));   // verilog/coms.v(154[7:23])
    defparam equal_59_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1367 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42419), .I3(\FRAME_MATCHER.i [0]), .O(n42424));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1367.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1368 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42403), .I3(\FRAME_MATCHER.i [0]), .O(n42405));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1368.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1369 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42411), .I3(\FRAME_MATCHER.i [0]), .O(n42413));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1369.LUT_INIT = 16'hfeff;
    uart_tx tx (.n23609(n23609), .r_Clock_Count({\r_Clock_Count[8] , \r_Clock_Count[7] , 
            \r_Clock_Count[6] , \r_Clock_Count[5] , \r_Clock_Count[4] , 
            \r_Clock_Count[3] , \r_Clock_Count[2] , \r_Clock_Count[1] , 
            Open_38}), .clk32MHz(clk32MHz), .n23612(n23612), .n23615(n23615), 
            .n23618(n23618), .n23621(n23621), .n23624(n23624), .n23627(n23627), 
            .n23630(n23630), .n23634(n23634), .r_Bit_Index({r_Bit_Index}), 
            .n23637(n23637), .n24235(n24235), .r_SM_Main({r_SM_Main}), 
            .n23680(n23680), .tx_data({tx_data}), .n313(n313), .GND_net(GND_net), 
            .n314(n314), .n315(n315), .n316(n316), .n317(n317), .n318(n318), 
            .\r_SM_Main_2__N_2753[1] (\r_SM_Main_2__N_2753[1] ), .n319(n319), 
            .n320(n320), .VCC_net(VCC_net), .n23629(n23629), .n23463(n23463), 
            .n23547(n23547), .n4032(n4032), .o_Tx_Serial_N_2784(o_Tx_Serial_N_2784), 
            .n49982(n49982), .n23583(n23583), .n23582(n23582), .tx_active(tx_active), 
            .n23581(n23581), .tx_o(tx_o), .\r_SM_Main_2__N_2756[0] (r_SM_Main_2__N_2756[0]), 
            .n23411(n23411), .n49(n49), .tx_enable(tx_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.VCC_net(VCC_net), .rx_data_ready(rx_data_ready), .clk32MHz(clk32MHz), 
            .n23640(n23640), .r_Bit_Index({r_Bit_Index_adj_12}), .n23643(n23643), 
            .n28961(n28961), .r_SM_Main({Open_39, \r_SM_Main[1]_adj_8 , 
            Open_40}), .n23683(n23683), .n24171(n24171), .rx_data({rx_data}), 
            .r_Rx_Data(r_Rx_Data), .PIN_13_N_26(PIN_13_N_26), .n46671(n46671), 
            .GND_net(GND_net), .n46670(n46670), .\r_SM_Main[2] (\r_SM_Main[2]_adj_9 ), 
            .n23457(n23457), .n23545(n23545), .n4010(n4010), .n23650(n23650), 
            .n23649(n23649), .n23648(n23648), .n23647(n23647), .n23646(n23646), 
            .n23645(n23645), .n23644(n23644), .n23579(n23579), .n22411(n22411), 
            .n4(n4), .n28925(n28925), .n1(n1), .n28462(n28462), .n4_adj_1(n4_adj_10), 
            .n4_adj_2(n4_adj_11), .n22416(n22416)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n23609, r_Clock_Count, clk32MHz, n23612, n23615, n23618, 
            n23621, n23624, n23627, n23630, n23634, r_Bit_Index, 
            n23637, n24235, r_SM_Main, n23680, tx_data, n313, GND_net, 
            n314, n315, n316, n317, n318, \r_SM_Main_2__N_2753[1] , 
            n319, n320, VCC_net, n23629, n23463, n23547, n4032, 
            o_Tx_Serial_N_2784, n49982, n23583, n23582, tx_active, 
            n23581, tx_o, \r_SM_Main_2__N_2756[0] , n23411, n49, tx_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n23609;
    output [8:0]r_Clock_Count;
    input clk32MHz;
    input n23612;
    input n23615;
    input n23618;
    input n23621;
    input n23624;
    input n23627;
    input n23630;
    input n23634;
    output [2:0]r_Bit_Index;
    input n23637;
    input n24235;
    output [2:0]r_SM_Main;
    input n23680;
    input [7:0]tx_data;
    output n313;
    input GND_net;
    output n314;
    output n315;
    output n316;
    output n317;
    output n318;
    output \r_SM_Main_2__N_2753[1] ;
    output n319;
    output n320;
    input VCC_net;
    output n23629;
    output n23463;
    output n23547;
    output n4032;
    output o_Tx_Serial_N_2784;
    input n49982;
    input n23583;
    input n23582;
    output tx_active;
    input n23581;
    output tx_o;
    input \r_SM_Main_2__N_2756[0] ;
    output n23411;
    output n49;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n42116;
    wire [8:0]r_Clock_Count_c;   // verilog/uart_tx.v(32[16:29])
    
    wire n19916;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n35939, n35938, n35937, n35936, n35935, n35934, n1, n35933, 
        n35932, n46705, n28884, n127, n10, n8, n44351, n44469, 
        n44470, n49842, n44401, n44400, n16844;
    
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n23609));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23612));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23615));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n23618));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23621));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23624));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n23627));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n23630));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23634));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23637));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n24235));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count_c[0]), .C(clk32MHz), .D(n42116));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n23680));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n35939), .O(n313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n35938), .O(n314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_9 (.CI(n35938), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n35939));
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n35937), .O(n315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n35937), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n35938));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n35936), .O(n316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n35936), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n35937));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n35935), .O(n317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n35935), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n35936));
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n35934), .O(n318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n35934), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n35935));
    SB_LUT4 i15197_2_lut (.I0(\r_SM_Main_2__N_2753[1] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i15197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n35933), .O(n319)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_4 (.CI(n35933), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n35934));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n35932), .O(n320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n35932), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n35933));
    SB_LUT4 add_59_2_lut (.I0(n23629), .I1(r_Clock_Count_c[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n46705)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count_c[0]), .I1(GND_net), 
            .CO(n35932));
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n28884));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[8]), .I1(n127), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[4]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[7]), .I1(n10), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_2753[1] ));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i10133_3_lut (.I0(n23463), .I1(r_SM_Main[1]), .I2(n28884), 
            .I3(GND_net), .O(n23547));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10133_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1092_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4032));   // verilog/uart_tx.v(98[36:51])
    defparam i1092_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count_c[0]), .I2(r_Clock_Count[2]), 
            .I3(r_Clock_Count[1]), .O(n127));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[4]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n8));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i28792_4_lut (.I0(r_Clock_Count[8]), .I1(n127), .I2(r_Clock_Count[7]), 
            .I3(r_Clock_Count[6]), .O(n44351));
    defparam i28792_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15011_4_lut (.I0(r_SM_Main[2]), .I1(r_Clock_Count[5]), .I2(n44351), 
            .I3(n8), .O(n23629));
    defparam i15011_4_lut.LUT_INIT = 16'habaa;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n44469), 
            .I2(n44470), .I3(r_Bit_Index[2]), .O(n49842));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n49842_bdd_4_lut (.I0(n49842), .I1(n44401), .I2(n44400), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_2784));
    defparam n49842_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n19916), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n49982));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n23583));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n23582));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n23581));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_2756[0] ), 
            .I3(r_SM_Main[1]), .O(n19916));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2753[1] ), .O(n23463));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i21_3_lut (.I0(r_Clock_Count_c[0]), .I1(n46705), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n42116));
    defparam i21_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2756[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n16844));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n16844), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n1), .O(n23411));
    defparam i2_4_lut.LUT_INIT = 16'h3202;
    SB_LUT4 i47_4_lut (.I0(\r_SM_Main_2__N_2756[0] ), .I1(n28884), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_2753[1] ), .O(n49));   // verilog/uart_tx.v(31[16:25])
    defparam i47_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i28841_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44400));
    defparam i28841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28842_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44401));
    defparam i28842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28911_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44470));
    defparam i28911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28910_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n44469));
    defparam i28910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12370_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(tx_enable));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12370_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (VCC_net, rx_data_ready, clk32MHz, n23640, r_Bit_Index, 
            n23643, n28961, r_SM_Main, n23683, n24171, rx_data, 
            r_Rx_Data, PIN_13_N_26, n46671, GND_net, n46670, \r_SM_Main[2] , 
            n23457, n23545, n4010, n23650, n23649, n23648, n23647, 
            n23646, n23645, n23644, n23579, n22411, n4, n28925, 
            n1, n28462, n4_adj_1, n4_adj_2, n22416) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input VCC_net;
    output rx_data_ready;
    input clk32MHz;
    input n23640;
    output [2:0]r_Bit_Index;
    input n23643;
    input n28961;
    output [2:0]r_SM_Main;
    input n23683;
    input n24171;
    output [7:0]rx_data;
    output r_Rx_Data;
    input PIN_13_N_26;
    output n46671;
    input GND_net;
    output n46670;
    output \r_SM_Main[2] ;
    output n23457;
    output n23545;
    output n4010;
    input n23650;
    input n23649;
    input n23648;
    input n23647;
    input n23646;
    input n23645;
    input n23644;
    input n23579;
    output n22411;
    output n4;
    output n28925;
    output n1;
    output n28462;
    output n4_adj_1;
    output n4_adj_2;
    output n22416;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n41862, n23588;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n23591, n23594, n23597, n23600, n23603, n41854, n23674, 
        r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_2682;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    wire [2:0]r_SM_Main_2__N_2688;
    
    wire n46647, n35931, n138, n46645, n35930, n46644, n35929, 
        n46648, n35928, n46646, n35927, n46650, n35926, n46693, 
        n35925, n46649, n42358, n28858, n43082, n42363, n8, n158, 
        n46699, n46700, n28, n28824, n44041, n22163, n23398;
    
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n41862));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23588));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23591));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n23594));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23597));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23600));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n23603));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n41854));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23640));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23643));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n28961));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n23674));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n23683));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n24171));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_26));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i31811_2_lut (.I0(r_SM_Main_2__N_2682[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46671));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i31811_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31519_3_lut (.I0(r_SM_Main_c[0]), .I1(r_SM_Main_2__N_2688[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n46670));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i31519_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 add_62_9_lut (.I0(n138), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n35931), .O(n46647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n138), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n35930), .O(n46645)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_8 (.CI(n35930), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n35931));
    SB_LUT4 add_62_7_lut (.I0(n138), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n35929), .O(n46644)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n35929), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n35930));
    SB_LUT4 add_62_6_lut (.I0(n138), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n35928), .O(n46648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n35928), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n35929));
    SB_LUT4 add_62_5_lut (.I0(n138), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n35927), .O(n46646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n35927), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n35928));
    SB_LUT4 add_62_4_lut (.I0(n138), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n35926), .O(n46650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_4 (.CI(n35926), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n35927));
    SB_LUT4 add_62_3_lut (.I0(n138), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n35925), .O(n46693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n35925), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n35926));
    SB_LUT4 add_62_2_lut (.I0(n138), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n46649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n35925));
    SB_DFFSR r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk32MHz), .D(r_SM_Main_2__N_2682[2]), 
            .R(n42358));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n28858));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(\r_SM_Main[2] ), .I1(r_SM_Main_2__N_2682[2]), 
            .I2(r_SM_Main_c[0]), .I3(r_SM_Main[1]), .O(n23457));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i10131_3_lut (.I0(n23457), .I1(n28858), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n23545));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10131_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1070_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4010));   // verilog/uart_rx.v(102[36:51])
    defparam i1070_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i11_3_lut (.I0(r_Clock_Count[1]), .I1(n46693), .I2(n43082), 
            .I3(GND_net), .O(n41854));
    defparam i11_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17002_3_lut (.I0(r_Clock_Count[2]), .I1(n46650), .I2(n43082), 
            .I3(GND_net), .O(n23603));
    defparam i17002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16976_3_lut (.I0(r_Clock_Count[3]), .I1(n46646), .I2(n43082), 
            .I3(GND_net), .O(n23600));
    defparam i16976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16990_3_lut (.I0(r_Clock_Count[4]), .I1(n46648), .I2(n43082), 
            .I3(GND_net), .O(n23597));
    defparam i16990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16964_3_lut (.I0(r_Clock_Count[5]), .I1(n46644), .I2(n43082), 
            .I3(GND_net), .O(n23594));
    defparam i16964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16970_3_lut (.I0(r_Clock_Count[6]), .I1(n46645), .I2(n43082), 
            .I3(GND_net), .O(n23591));
    defparam i16970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_3_lut (.I0(r_Clock_Count[3]), .I1(n42363), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i31870_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main_c[0]), .I2(n8), 
            .I3(n158), .O(n46699));
    defparam i31870_4_lut.LUT_INIT = 16'h3373;
    SB_LUT4 i1_4_lut (.I0(\r_SM_Main[2] ), .I1(n46699), .I2(n46700), .I3(r_SM_Main[1]), 
            .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_3_lut_adj_824 (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[2]), .I3(GND_net), .O(n28824));
    defparam i2_3_lut_adj_824.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_2__N_2688[0]), .I2(r_Rx_Data), 
            .I3(r_SM_Main_c[0]), .O(n44041));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i27532_3_lut (.I0(\r_SM_Main[2] ), .I1(n28), .I2(n44041), 
            .I3(GND_net), .O(n43082));
    defparam i27532_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i16984_3_lut (.I0(r_Clock_Count[7]), .I1(n46647), .I2(n43082), 
            .I3(GND_net), .O(n23588));
    defparam i16984_3_lut.LUT_INIT = 16'hacac;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n23650));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n23649));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n23648));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n23647));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n23646));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n23645));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n23644));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n23579));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_3_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n158));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_825 (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), 
            .I2(r_Clock_Count[1]), .I3(GND_net), .O(n42363));
    defparam i2_3_lut_adj_825.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut_adj_826 (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(\r_SM_Main[2] ), 
            .I3(r_SM_Main_2__N_2682[2]), .O(n22163));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut_adj_826.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(r_Bit_Index[0]), .I1(n22163), .I2(GND_net), 
            .I3(GND_net), .O(n22411));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_75_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_75_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16996_3_lut (.I0(r_Clock_Count[0]), .I1(n46649), .I2(n43082), 
            .I3(GND_net), .O(n23674));
    defparam i16996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n28858), .I1(r_SM_Main_2__N_2682[2]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n28925));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_2688[0]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i15068_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n28462));
    defparam i15068_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_71_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_71_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_73_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_73_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_827 (.I0(n22163), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n22416));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_827.LUT_INIT = 16'hbbbb;
    SB_LUT4 i34249_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n42358));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34249_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), .I2(r_SM_Main_2__N_2682[2]), 
            .I3(r_SM_Main_c[0]), .O(n23398));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), .I2(n23398), 
            .I3(rx_data_ready), .O(n41862));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i31868_3_lut_4_lut (.I0(n158), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[3]), 
            .I3(n28824), .O(n46700));
    defparam i31868_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_3_lut_4_lut (.I0(n158), .I1(r_Clock_Count[7]), .I2(n28824), 
            .I3(r_Clock_Count[3]), .O(r_SM_Main_2__N_2688[0]));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i15473_3_lut_4_lut (.I0(n158), .I1(r_Clock_Count[7]), .I2(n42363), 
            .I3(r_Clock_Count[3]), .O(r_SM_Main_2__N_2682[2]));
    defparam i15473_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i29_1_lut_4_lut (.I0(\r_SM_Main[2] ), .I1(n46699), .I2(n46700), 
            .I3(r_SM_Main[1]), .O(n138));
    defparam i29_1_lut_4_lut.LUT_INIT = 16'hafbb;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n2276, encoder0_position, GND_net, 
            data_o, clk32MHz, n23706, n23705, n23704, n23703, n23702, 
            n23701, n23700, n23699, n23698, n23697, n23696, n23695, 
            n23694, n23693, n23692, n23691, n23690, n23689, n23688, 
            n23687, n23686, n23685, n23684, n23576, count_enable, 
            n24227, reg_B, n44196, PIN_23_c_1, PIN_24_c_0, n23578) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n2276;
    output [23:0]encoder0_position;
    input GND_net;
    output [1:0]data_o;
    input clk32MHz;
    input n23706;
    input n23705;
    input n23704;
    input n23703;
    input n23702;
    input n23701;
    input n23700;
    input n23699;
    input n23698;
    input n23697;
    input n23696;
    input n23695;
    input n23694;
    input n23693;
    input n23692;
    input n23691;
    input n23690;
    input n23689;
    input n23688;
    input n23687;
    input n23686;
    input n23685;
    input n23684;
    input n23576;
    output count_enable;
    input n24227;
    output [1:0]reg_B;
    output n44196;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n23578;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n2272, n35957, n35958, n35956, n35955, n35954, n35953, 
        n35952, n35951, n35950, n35949, n35948, n35947, n35946, 
        B_delayed, A_delayed, n35945, n35944, n35943, n35942, n35941, 
        count_direction, n35940, n35963, n35962, n35961, n35960, 
        n35959;
    
    SB_LUT4 add_533_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2272), 
            .I3(n35957), .O(n2276[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_19 (.CI(n35957), .I0(encoder0_position[17]), .I1(n2272), 
            .CO(n35958));
    SB_LUT4 add_533_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2272), 
            .I3(n35956), .O(n2276[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_18 (.CI(n35956), .I0(encoder0_position[16]), .I1(n2272), 
            .CO(n35957));
    SB_LUT4 add_533_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2272), 
            .I3(n35955), .O(n2276[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_17 (.CI(n35955), .I0(encoder0_position[15]), .I1(n2272), 
            .CO(n35956));
    SB_LUT4 add_533_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2272), 
            .I3(n35954), .O(n2276[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_16 (.CI(n35954), .I0(encoder0_position[14]), .I1(n2272), 
            .CO(n35955));
    SB_LUT4 add_533_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2272), 
            .I3(n35953), .O(n2276[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_15 (.CI(n35953), .I0(encoder0_position[13]), .I1(n2272), 
            .CO(n35954));
    SB_LUT4 add_533_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2272), 
            .I3(n35952), .O(n2276[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_14 (.CI(n35952), .I0(encoder0_position[12]), .I1(n2272), 
            .CO(n35953));
    SB_LUT4 add_533_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2272), 
            .I3(n35951), .O(n2276[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_13 (.CI(n35951), .I0(encoder0_position[11]), .I1(n2272), 
            .CO(n35952));
    SB_LUT4 add_533_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2272), 
            .I3(n35950), .O(n2276[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_12 (.CI(n35950), .I0(encoder0_position[10]), .I1(n2272), 
            .CO(n35951));
    SB_LUT4 add_533_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2272), 
            .I3(n35949), .O(n2276[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_11 (.CI(n35949), .I0(encoder0_position[9]), .I1(n2272), 
            .CO(n35950));
    SB_LUT4 add_533_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2272), 
            .I3(n35948), .O(n2276[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_10 (.CI(n35948), .I0(encoder0_position[8]), .I1(n2272), 
            .CO(n35949));
    SB_LUT4 add_533_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2272), 
            .I3(n35947), .O(n2276[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_9 (.CI(n35947), .I0(encoder0_position[7]), .I1(n2272), 
            .CO(n35948));
    SB_LUT4 add_533_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2272), 
            .I3(n35946), .O(n2276[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_533_8 (.CI(n35946), .I0(encoder0_position[6]), .I1(n2272), 
            .CO(n35947));
    SB_LUT4 add_533_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2272), 
            .I3(n35945), .O(n2276[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_7 (.CI(n35945), .I0(encoder0_position[5]), .I1(n2272), 
            .CO(n35946));
    SB_LUT4 add_533_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2272), 
            .I3(n35944), .O(n2276[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_6 (.CI(n35944), .I0(encoder0_position[4]), .I1(n2272), 
            .CO(n35945));
    SB_LUT4 add_533_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2272), 
            .I3(n35943), .O(n2276[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_5 (.CI(n35943), .I0(encoder0_position[3]), .I1(n2272), 
            .CO(n35944));
    SB_LUT4 add_533_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2272), 
            .I3(n35942), .O(n2276[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_4 (.CI(n35942), .I0(encoder0_position[2]), .I1(n2272), 
            .CO(n35943));
    SB_LUT4 add_533_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2272), 
            .I3(n35941), .O(n2276[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_3 (.CI(n35941), .I0(encoder0_position[1]), .I1(n2272), 
            .CO(n35942));
    SB_LUT4 add_533_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n35940), .O(n2276[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_2 (.CI(n35940), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n35941));
    SB_CARRY add_533_1 (.CI(GND_net), .I0(n2272), .I1(n2272), .CO(n35940));
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n23706));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n23705));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n23704));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n23703));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n23702));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n23701));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n23700));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n23699));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n23698));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n23697));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n23696));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n23695));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n23694));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n23693));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n23692));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n23691));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n23690));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n23689));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n23688));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n23687));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n23686));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n23685));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n23684));   // quad.v(35[10] 41[6])
    SB_LUT4 add_533_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2272), 
            .I3(n35963), .O(n2276[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_533_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2272), 
            .I3(n35962), .O(n2276[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_24 (.CI(n35962), .I0(encoder0_position[22]), .I1(n2272), 
            .CO(n35963));
    SB_LUT4 add_533_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2272), 
            .I3(n35961), .O(n2276[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_23 (.CI(n35961), .I0(encoder0_position[21]), .I1(n2272), 
            .CO(n35962));
    SB_LUT4 add_533_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2272), 
            .I3(n35960), .O(n2276[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_22 (.CI(n35960), .I0(encoder0_position[20]), .I1(n2272), 
            .CO(n35961));
    SB_LUT4 add_533_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2272), 
            .I3(n35959), .O(n2276[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_21 (.CI(n35959), .I0(encoder0_position[19]), .I1(n2272), 
            .CO(n35960));
    SB_LUT4 add_533_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2272), 
            .I3(n35958), .O(n2276[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_533_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_533_20 (.CI(n35958), .I0(encoder0_position[18]), .I1(n2272), 
            .CO(n35959));
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n23576));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i755_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // quad.v(37[5] 40[8])
    defparam i755_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n24227(n24227), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .n44196(n44196), .GND_net(GND_net), 
            .PIN_23_c_1(PIN_23_c_1), .PIN_24_c_0(PIN_24_c_0), .n23578(n23578)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n24227, data_o, clk32MHz, reg_B, n44196, 
            GND_net, PIN_23_c_1, PIN_24_c_0, n23578) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24227;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    output n44196;
    input GND_net;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n23578;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n1, cnt_next_2__N_3113;
    wire [2:0]n17;
    
    wire n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24227));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[2]), 
            .I3(GND_net), .O(n44196));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_23_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1016__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n1), .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_24_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23578));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1016__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1016__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22267_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22267_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22260_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22260_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n44196), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3113));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i1244_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(170[42:59])
    defparam i1244_1_lut.LUT_INIT = 16'h5555;
    
endmodule
