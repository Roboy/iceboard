-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Jan 29 2020 19:19:01

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n2553_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal n2554 : std_logic;
signal n26 : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal n25 : std_logic;
signal n2294 : std_logic;
signal n24 : std_logic;
signal n2295 : std_logic;
signal n23 : std_logic;
signal n2296 : std_logic;
signal n22 : std_logic;
signal n2297 : std_logic;
signal n21 : std_logic;
signal n2298 : std_logic;
signal n20 : std_logic;
signal n2299 : std_logic;
signal n19 : std_logic;
signal n2300 : std_logic;
signal n2301 : std_logic;
signal n18 : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal n17 : std_logic;
signal n2302 : std_logic;
signal n16 : std_logic;
signal n2303 : std_logic;
signal n15 : std_logic;
signal n2304 : std_logic;
signal n14 : std_logic;
signal n2305 : std_logic;
signal n13 : std_logic;
signal n2306 : std_logic;
signal n12 : std_logic;
signal n2307 : std_logic;
signal n11 : std_logic;
signal n2308 : std_logic;
signal n2309 : std_logic;
signal n10 : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal n9 : std_logic;
signal n2310 : std_logic;
signal n8_adj_409 : std_logic;
signal n2311 : std_logic;
signal n7 : std_logic;
signal n2312 : std_logic;
signal n6_adj_410 : std_logic;
signal n2313 : std_logic;
signal blink_counter_21 : std_logic;
signal n2314 : std_logic;
signal blink_counter_22 : std_logic;
signal n2315 : std_logic;
signal blink_counter_23 : std_logic;
signal n2316 : std_logic;
signal n2317 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal n2318 : std_logic;
signal blink_counter_25 : std_logic;
signal \n693_cascade_\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal n2263 : std_logic;
signal n2264 : std_logic;
signal n2265 : std_logic;
signal n2266 : std_logic;
signal n2267 : std_logic;
signal n2268 : std_logic;
signal n2269 : std_logic;
signal n2270 : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal n2271 : std_logic;
signal n2272 : std_logic;
signal n2273 : std_logic;
signal n2274 : std_logic;
signal n2275 : std_logic;
signal n2276 : std_logic;
signal n2277 : std_logic;
signal n2278 : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal n2279 : std_logic;
signal n2280 : std_logic;
signal n2281 : std_logic;
signal n2282 : std_logic;
signal n2283 : std_logic;
signal n2284 : std_logic;
signal n2285 : std_logic;
signal n2286 : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal n2287 : std_logic;
signal n2288 : std_logic;
signal n2289 : std_logic;
signal n2290 : std_logic;
signal n2291 : std_logic;
signal n2292 : std_logic;
signal n2293 : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \eeprom.n2241\ : std_logic;
signal \eeprom.delay_counter_2\ : std_logic;
signal \eeprom.delay_counter_15_N_171_2\ : std_logic;
signal \eeprom.n2242\ : std_logic;
signal \eeprom.n2243\ : std_logic;
signal \eeprom.n2244\ : std_logic;
signal \eeprom.n2245\ : std_logic;
signal \eeprom.delay_counter_6\ : std_logic;
signal \eeprom.delay_counter_15_N_171_6\ : std_logic;
signal \eeprom.n2246\ : std_logic;
signal \eeprom.n2247\ : std_logic;
signal \eeprom.n2248\ : std_logic;
signal \eeprom.delay_counter_8\ : std_logic;
signal \eeprom.delay_counter_15_N_171_8\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \eeprom.n2249\ : std_logic;
signal \eeprom.n2250\ : std_logic;
signal \eeprom.n2251\ : std_logic;
signal \eeprom.delay_counter_12\ : std_logic;
signal \eeprom.delay_counter_15_N_171_12\ : std_logic;
signal \eeprom.n2252\ : std_logic;
signal \eeprom.n2253\ : std_logic;
signal \eeprom.n2254\ : std_logic;
signal \eeprom.n642\ : std_logic;
signal \eeprom.n2255\ : std_logic;
signal \eeprom.n14\ : std_logic;
signal \eeprom.n13_cascade_\ : std_logic;
signal \eeprom.n7_cascade_\ : std_logic;
signal \eeprom.delay_counter_15_N_171_1\ : std_logic;
signal \eeprom.delay_counter_1\ : std_logic;
signal \eeprom.delay_counter_15_N_171_0\ : std_logic;
signal \eeprom.delay_counter_0\ : std_logic;
signal \eeprom.delay_counter_15_N_171_5\ : std_logic;
signal \eeprom.delay_counter_5\ : std_logic;
signal \eeprom.delay_counter_15_N_171_10\ : std_logic;
signal \eeprom.delay_counter_10\ : std_logic;
signal \eeprom.delay_counter_15_N_171_4\ : std_logic;
signal \eeprom.delay_counter_4\ : std_logic;
signal n324 : std_logic;
signal \eeprom.n1500\ : std_logic;
signal \n6_adj_405_cascade_\ : std_logic;
signal n41 : std_logic;
signal \eeprom.n1018\ : std_logic;
signal \n2483_cascade_\ : std_logic;
signal \eeprom.n2453\ : std_logic;
signal \n1568_cascade_\ : std_logic;
signal state_1 : std_logic;
signal n1568 : std_logic;
signal delay_counter_7 : std_logic;
signal delay_counter_8 : std_logic;
signal delay_counter_1 : std_logic;
signal delay_counter_4 : std_logic;
signal delay_counter_10 : std_logic;
signal delay_counter_12 : std_logic;
signal delay_counter_11 : std_logic;
signal delay_counter_13 : std_logic;
signal \n2512_cascade_\ : std_logic;
signal delay_counter_16 : std_logic;
signal delay_counter_18 : std_logic;
signal \n2495_cascade_\ : std_logic;
signal delay_counter_19 : std_logic;
signal delay_counter_9 : std_logic;
signal delay_counter_6 : std_logic;
signal delay_counter_3 : std_logic;
signal delay_counter_0 : std_logic;
signal delay_counter_17 : std_logic;
signal delay_counter_15 : std_logic;
signal delay_counter_14 : std_logic;
signal n8 : std_logic;
signal delay_counter_21 : std_logic;
signal delay_counter_23 : std_logic;
signal n6_adj_413 : std_logic;
signal delay_counter_5 : std_logic;
signal n16_adj_407 : std_logic;
signal delay_counter_2 : std_logic;
signal n17_adj_406 : std_logic;
signal n2536 : std_logic;
signal \read_N\ : std_logic;
signal delay_counter_22 : std_logic;
signal delay_counter_25 : std_logic;
signal delay_counter_20 : std_logic;
signal n8_adj_412 : std_logic;
signal n9_adj_404 : std_logic;
signal delay_counter_31 : std_logic;
signal \n9_adj_404_cascade_\ : std_logic;
signal \addr_10__N_70\ : std_logic;
signal delay_counter_29 : std_logic;
signal delay_counter_28 : std_logic;
signal n10_adj_403 : std_logic;
signal delay_counter_26 : std_logic;
signal delay_counter_30 : std_logic;
signal delay_counter_27 : std_logic;
signal delay_counter_24 : std_logic;
signal n14_adj_401 : std_logic;
signal \eeprom.delay_counter_15_N_171_7\ : std_logic;
signal \eeprom.delay_counter_15_N_171_3\ : std_logic;
signal \eeprom.delay_counter_3\ : std_logic;
signal \eeprom.delay_counter_15_N_171_11\ : std_logic;
signal \eeprom.delay_counter_15_N_171_9\ : std_logic;
signal \eeprom.delay_counter_11\ : std_logic;
signal \eeprom.delay_counter_7\ : std_logic;
signal \eeprom.n6_cascade_\ : std_logic;
signal \eeprom.delay_counter_9\ : std_logic;
signal \eeprom.n8\ : std_logic;
signal \eeprom.delay_counter_15_N_171_15\ : std_logic;
signal \eeprom.delay_counter_15\ : std_logic;
signal \eeprom.delay_counter_15_N_171_14\ : std_logic;
signal \eeprom.delay_counter_14\ : std_logic;
signal state_0 : std_logic;
signal \eeprom.n1601\ : std_logic;
signal \eeprom.delay_counter_15_N_171_13\ : std_logic;
signal \eeprom.delay_counter_13\ : std_logic;
signal \INVeeprom.i2c.write_enable_132C_net\ : std_logic;
signal \n11_adj_399_cascade_\ : std_logic;
signal \eeprom.i2c.n1669\ : std_logic;
signal \eeprom.i2c.n37_cascade_\ : std_logic;
signal \eeprom.i2c.n33\ : std_logic;
signal \eeprom.i2c.n39_cascade_\ : std_logic;
signal \eeprom.i2c.n1027\ : std_logic;
signal \eeprom.i2c.n11_adj_379\ : std_logic;
signal \INVeeprom.i2c.sda_out_133C_net\ : std_logic;
signal \eeprom.i2c.n6_cascade_\ : std_logic;
signal \eeprom.i2c.counter2_7__N_256_cascade_\ : std_logic;
signal \eeprom.i2c.n1580\ : std_logic;
signal rw : std_logic;
signal \n1835_cascade_\ : std_logic;
signal n2569 : std_logic;
signal \n949_cascade_\ : std_logic;
signal n949 : std_logic;
signal \n2547_cascade_\ : std_logic;
signal \eeprom.i2c.n2574_cascade_\ : std_logic;
signal \eeprom.i2c.n2557\ : std_logic;
signal \eeprom.enable\ : std_logic;
signal \n2538_cascade_\ : std_logic;
signal \n4_adj_411_cascade_\ : std_logic;
signal n1835 : std_logic;
signal \n2507_cascade_\ : std_logic;
signal n10_adj_394 : std_logic;
signal saved_addr_0 : std_logic;
signal n11_adj_399 : std_logic;
signal n2566 : std_logic;
signal \eeprom.i2c.n39\ : std_logic;
signal \eeprom.i2c.n2406\ : std_logic;
signal \eeprom.i2c.n37\ : std_logic;
signal \eeprom.i2c.n1051_cascade_\ : std_logic;
signal \eeprom.i2c.n13\ : std_logic;
signal sda_out : std_logic;
signal sda_enable : std_logic;
signal \state_7_N_285_3_cascade_\ : std_logic;
signal \eeprom.i2c.n2475\ : std_logic;
signal \eeprom.i2c.n2475_cascade_\ : std_logic;
signal \eeprom.i2c.n9\ : std_logic;
signal \eeprom.i2c.counter2_0\ : std_logic;
signal \bfn_21_18_0_\ : std_logic;
signal \eeprom.i2c.counter2_1\ : std_logic;
signal \eeprom.i2c.n2319\ : std_logic;
signal \eeprom.i2c.counter2_2\ : std_logic;
signal \eeprom.i2c.n2320\ : std_logic;
signal \eeprom.i2c.counter2_3\ : std_logic;
signal \eeprom.i2c.n2321\ : std_logic;
signal \eeprom.i2c.n2322\ : std_logic;
signal \eeprom.i2c.counter2_4\ : std_logic;
signal \CLK_N\ : std_logic;
signal \eeprom.i2c.counter2_7__N_256\ : std_logic;
signal n306 : std_logic;
signal \n10_adj_398_cascade_\ : std_logic;
signal \state_7_N_269_0\ : std_logic;
signal \n2460_cascade_\ : std_logic;
signal n2560 : std_logic;
signal n308 : std_logic;
signal n320 : std_logic;
signal n318 : std_logic;
signal n1817 : std_logic;
signal \eeprom.i2c.n12_cascade_\ : std_logic;
signal n4_adj_408 : std_logic;
signal \eeprom.i2c.n942\ : std_logic;
signal n10_adj_398 : std_logic;
signal n11_adj_400 : std_logic;
signal \eeprom.i2c.n942_cascade_\ : std_logic;
signal n1532 : std_logic;
signal \eeprom.i2c.counter_0\ : std_logic;
signal \bfn_21_22_0_\ : std_logic;
signal \eeprom.i2c.n2256\ : std_logic;
signal \eeprom.i2c.n2257\ : std_logic;
signal \eeprom.i2c.counter_3\ : std_logic;
signal \eeprom.i2c.n2258\ : std_logic;
signal \eeprom.i2c.counter_4\ : std_logic;
signal \eeprom.i2c.n2259\ : std_logic;
signal \eeprom.i2c.counter_5\ : std_logic;
signal \eeprom.i2c.n2260\ : std_logic;
signal \eeprom.i2c.counter_6\ : std_logic;
signal \eeprom.i2c.n2261\ : std_logic;
signal \eeprom.i2c.n2262\ : std_logic;
signal \eeprom.i2c.counter_7\ : std_logic;
signal \eeprom.i2c.n1548\ : std_logic;
signal \eeprom.i2c.n1655\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n15_adj_393 : std_logic;
signal \eeprom.i2c.n10_cascade_\ : std_logic;
signal \INVeeprom.i2c.i2c_scl_enable_124C_net\ : std_logic;
signal state_2 : std_logic;
signal state_0_adj_397 : std_logic;
signal state_1_adj_396 : std_logic;
signal state_3 : std_logic;
signal n1826 : std_logic;
signal n314 : std_logic;
signal n1518 : std_logic;
signal \n4_adj_395_cascade_\ : std_logic;
signal n310 : std_logic;
signal n4_adj_395 : std_logic;
signal n312 : std_logic;
signal \eeprom.i2c.counter_1\ : std_logic;
signal \eeprom.i2c.counter_2\ : std_logic;
signal n4 : std_logic;
signal n1523 : std_logic;
signal \n4_cascade_\ : std_logic;
signal \state_7_N_285_3\ : std_logic;
signal n316 : std_logic;
signal scl_enable : std_logic;
signal \eeprom.i2c.i2c_clk\ : std_logic;
signal scl_c : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6589\,
            DIN => \N__6588\,
            DOUT => \N__6587\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6589\,
            PADOUT => \N__6588\,
            PADIN => \N__6587\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6580\,
            DIN => \N__6579\,
            DOUT => \N__6578\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6580\,
            PADOUT => \N__6579\,
            PADIN => \N__6578\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6571\,
            DIN => \N__6570\,
            DOUT => \N__6569\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6571\,
            PADOUT => \N__6570\,
            PADIN => \N__6569\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6562\,
            DIN => \N__6561\,
            DOUT => \N__6560\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6562\,
            PADOUT => \N__6561\,
            PADIN => \N__6560\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6553\,
            DIN => \N__6552\,
            DOUT => \N__6551\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6553\,
            PADOUT => \N__6552\,
            PADIN => \N__6551\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6544\,
            DIN => \N__6543\,
            DOUT => \N__6542\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6544\,
            PADOUT => \N__6543\,
            PADIN => \N__6542\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6535\,
            DIN => \N__6534\,
            DOUT => \N__6533\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6535\,
            PADOUT => \N__6534\,
            PADIN => \N__6533\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6526\,
            DIN => \N__6525\,
            DOUT => \N__6524\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6526\,
            PADOUT => \N__6525\,
            PADIN => \N__6524\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6517\,
            DIN => \N__6516\,
            DOUT => \N__6515\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6517\,
            PADOUT => \N__6516\,
            PADIN => \N__6515\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6508\,
            DIN => \N__6507\,
            DOUT => \N__6506\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6508\,
            PADOUT => \N__6507\,
            PADIN => \N__6506\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2838\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6499\,
            DIN => \N__6498\,
            DOUT => \N__6497\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6499\,
            PADOUT => \N__6498\,
            PADIN => \N__6497\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6490\,
            DIN => \N__6489\,
            DOUT => \N__6488\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6490\,
            PADOUT => \N__6489\,
            PADIN => \N__6488\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6481\,
            DIN => \N__6480\,
            DOUT => \N__6479\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6481\,
            PADOUT => \N__6480\,
            PADIN => \N__6479\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \scl_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__6472\,
            DIN => \N__6471\,
            DOUT => \N__6470\,
            PACKAGEPIN => SCL
        );

    \scl_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6472\,
            PADOUT => \N__6471\,
            PADIN => \N__6470\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6063\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__6207\
        );

    \sda_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__6463\,
            DIN => \N__6462\,
            DOUT => \N__6461\,
            PACKAGEPIN => SDA
        );

    \sda_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6463\,
            PADOUT => \N__6462\,
            PADIN => \N__6461\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__6282\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__4941\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6454\,
            DIN => \N__6453\,
            DOUT => \N__6452\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6454\,
            PADOUT => \N__6453\,
            PADIN => \N__6452\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1455\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6428\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6434\,
            I => \N__6428\
        );

    \I__1453\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6425\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6428\,
            I => \N__6421\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__6425\,
            I => \N__6418\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6415\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__6421\,
            I => n1518
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__6418\,
            I => n1518
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6415\,
            I => n1518
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__6408\,
            I => \n4_adj_395_cascade_\
        );

    \I__1445\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6402\,
            I => n310
        );

    \I__1443\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6396\,
            I => n4_adj_395
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6387\,
            I => n312
        );

    \I__1438\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6374\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6374\
        );

    \I__1436\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6371\
        );

    \I__1435\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6366\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6380\,
            I => \N__6366\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6379\,
            I => \N__6363\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6374\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6371\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6366\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6363\,
            I => \eeprom.i2c.counter_1\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__6354\,
            I => \N__6349\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6341\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6341\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6338\
        );

    \I__1424\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6335\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6332\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6329\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6341\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6338\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__6335\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6332\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6329\,
            I => \eeprom.i2c.counter_2\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6315\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6315\,
            I => n4
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__6312\,
            I => \N__6307\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6301\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6301\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6296\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6296\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6301\,
            I => \N__6293\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6290\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__6293\,
            I => n1523
        );

    \I__1406\ : Odrv4
    port map (
            O => \N__6290\,
            I => n1523
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__6285\,
            I => \n4_cascade_\
        );

    \I__1404\ : IoInMux
    port map (
            O => \N__6282\,
            I => \N__6279\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6279\,
            I => \N__6276\
        );

    \I__1402\ : Span4Mux_s0_h
    port map (
            O => \N__6276\,
            I => \N__6273\
        );

    \I__1401\ : Sp12to4
    port map (
            O => \N__6273\,
            I => \N__6270\
        );

    \I__1400\ : Span12Mux_v
    port map (
            O => \N__6270\,
            I => \N__6262\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6259\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6247\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6247\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6247\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6247\
        );

    \I__1394\ : Span12Mux_h
    port map (
            O => \N__6262\,
            I => \N__6242\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6259\,
            I => \N__6239\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6232\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6257\,
            I => \N__6232\
        );

    \I__1390\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6232\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6247\,
            I => \N__6229\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6224\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6224\
        );

    \I__1386\ : Odrv12
    port map (
            O => \N__6242\,
            I => \state_7_N_285_3\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__6239\,
            I => \state_7_N_285_3\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__6232\,
            I => \state_7_N_285_3\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__6229\,
            I => \state_7_N_285_3\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__6224\,
            I => \state_7_N_285_3\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6210\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6210\,
            I => n316
        );

    \I__1379\ : IoInMux
    port map (
            O => \N__6207\,
            I => \N__6204\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6204\,
            I => \N__6201\
        );

    \I__1377\ : IoSpan4Mux
    port map (
            O => \N__6201\,
            I => \N__6198\
        );

    \I__1376\ : Span4Mux_s2_h
    port map (
            O => \N__6198\,
            I => \N__6195\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__6195\,
            I => \N__6191\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6188\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__6191\,
            I => scl_enable
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6188\,
            I => scl_enable
        );

    \I__1371\ : ClkMux
    port map (
            O => \N__6183\,
            I => \N__6177\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6174\
        );

    \I__1369\ : ClkMux
    port map (
            O => \N__6181\,
            I => \N__6171\
        );

    \I__1368\ : ClkMux
    port map (
            O => \N__6180\,
            I => \N__6166\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__6177\,
            I => \N__6162\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6157\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6157\
        );

    \I__1364\ : ClkMux
    port map (
            O => \N__6170\,
            I => \N__6154\
        );

    \I__1363\ : ClkMux
    port map (
            O => \N__6169\,
            I => \N__6150\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6166\,
            I => \N__6147\
        );

    \I__1361\ : ClkMux
    port map (
            O => \N__6165\,
            I => \N__6144\
        );

    \I__1360\ : Span4Mux_v
    port map (
            O => \N__6162\,
            I => \N__6137\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__6157\,
            I => \N__6137\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6154\,
            I => \N__6137\
        );

    \I__1357\ : ClkMux
    port map (
            O => \N__6153\,
            I => \N__6134\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6131\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__6147\,
            I => \N__6126\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6144\,
            I => \N__6123\
        );

    \I__1353\ : Span4Mux_h
    port map (
            O => \N__6137\,
            I => \N__6118\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6134\,
            I => \N__6118\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__6131\,
            I => \N__6114\
        );

    \I__1350\ : ClkMux
    port map (
            O => \N__6130\,
            I => \N__6111\
        );

    \I__1349\ : ClkMux
    port map (
            O => \N__6129\,
            I => \N__6107\
        );

    \I__1348\ : Span4Mux_h
    port map (
            O => \N__6126\,
            I => \N__6103\
        );

    \I__1347\ : Span4Mux_h
    port map (
            O => \N__6123\,
            I => \N__6100\
        );

    \I__1346\ : Sp12to4
    port map (
            O => \N__6118\,
            I => \N__6097\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6094\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__6114\,
            I => \N__6089\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6089\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6086\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6107\,
            I => \N__6083\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6080\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__6103\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__6100\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1337\ : Odrv12
    port map (
            O => \N__6097\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6094\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__6089\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6086\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__6083\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6080\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1331\ : IoInMux
    port map (
            O => \N__6063\,
            I => \N__6060\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6060\,
            I => \N__6057\
        );

    \I__1329\ : Sp12to4
    port map (
            O => \N__6057\,
            I => \N__6054\
        );

    \I__1328\ : Odrv12
    port map (
            O => \N__6054\,
            I => scl_c
        );

    \I__1327\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6047\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6044\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6047\,
            I => \eeprom.i2c.counter_5\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6044\,
            I => \eeprom.i2c.counter_5\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6039\,
            I => \eeprom.i2c.n2260\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__6036\,
            I => \N__6033\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6029\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6026\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6029\,
            I => \eeprom.i2c.counter_6\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6026\,
            I => \eeprom.i2c.counter_6\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6021\,
            I => \eeprom.i2c.n2261\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6018\,
            I => \eeprom.i2c.n2262\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6011\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6008\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6011\,
            I => \eeprom.i2c.counter_7\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6008\,
            I => \eeprom.i2c.counter_7\
        );

    \I__1311\ : CEMux
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6000\,
            I => \eeprom.i2c.n1548\
        );

    \I__1309\ : SRMux
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__5991\,
            I => \eeprom.i2c.n1655\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__5988\,
            I => \N__5981\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__5987\,
            I => \N__5977\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__5986\,
            I => \N__5973\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5958\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5958\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5958\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5958\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5958\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5958\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5958\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__5955\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__5952\,
            I => \N__5948\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5939\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5939\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5936\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__5946\,
            I => \N__5933\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__5945\,
            I => \N__5930\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__5944\,
            I => \N__5926\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5923\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5936\,
            I => \N__5920\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5933\,
            I => \N__5917\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5910\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5910\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5910\
        );

    \I__1281\ : Span4Mux_h
    port map (
            O => \N__5923\,
            I => \N__5905\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__5920\,
            I => \N__5902\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5917\,
            I => \N__5897\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5910\,
            I => \N__5897\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5894\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5891\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__5905\,
            I => n15_adj_393
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__5902\,
            I => n15_adj_393
        );

    \I__1273\ : Odrv12
    port map (
            O => \N__5897\,
            I => n15_adj_393
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5894\,
            I => n15_adj_393
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5891\,
            I => n15_adj_393
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__5880\,
            I => \eeprom.i2c.n10_cascade_\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5867\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5862\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5862\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5854\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5845\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5845\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5845\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5845\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5834\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5862\,
            I => \N__5831\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5828\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5825\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5818\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5818\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5818\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5854\,
            I => \N__5813\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__5845\,
            I => \N__5813\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5804\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5843\,
            I => \N__5804\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5804\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5804\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5795\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5795\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5795\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5795\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__5834\,
            I => state_2
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__5831\,
            I => state_2
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5828\,
            I => state_2
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5825\,
            I => state_2
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5818\,
            I => state_2
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__5813\,
            I => state_2
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5804\,
            I => state_2
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5795\,
            I => state_2
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__5778\,
            I => \N__5773\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5762\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5776\,
            I => \N__5751\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5751\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5751\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5746\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5746\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5738\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5735\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5728\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5728\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5728\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5762\,
            I => \N__5721\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5718\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5715\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5710\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5710\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5751\,
            I => \N__5705\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5705\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5694\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5694\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5694\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5694\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5694\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5687\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5735\,
            I => \N__5687\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5728\,
            I => \N__5687\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5678\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5678\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5678\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5678\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__5721\,
            I => state_0_adj_397
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5718\,
            I => state_0_adj_397
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5715\,
            I => state_0_adj_397
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5710\,
            I => state_0_adj_397
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__5705\,
            I => state_0_adj_397
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5694\,
            I => state_0_adj_397
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__5687\,
            I => state_0_adj_397
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5678\,
            I => state_0_adj_397
        );

    \I__1197\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5657\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__5660\,
            I => \N__5654\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5657\,
            I => \N__5645\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5640\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5640\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5632\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5632\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__5650\,
            I => \N__5626\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__5649\,
            I => \N__5620\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__5648\,
            I => \N__5612\
        );

    \I__1187\ : Span4Mux_h
    port map (
            O => \N__5645\,
            I => \N__5607\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5640\,
            I => \N__5607\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5600\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5600\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5600\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5632\,
            I => \N__5597\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5588\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5588\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5588\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5588\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5581\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5581\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5581\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5578\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5565\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5565\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5565\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5565\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5565\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5565\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__5607\,
            I => state_1_adj_396
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5600\,
            I => state_1_adj_396
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__5597\,
            I => state_1_adj_396
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5588\,
            I => state_1_adj_396
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5581\,
            I => state_1_adj_396
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5578\,
            I => state_1_adj_396
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5565\,
            I => state_1_adj_396
        );

    \I__1160\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5545\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5540\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5540\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5545\,
            I => \N__5529\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5540\,
            I => \N__5526\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__5539\,
            I => \N__5518\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5510\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5510\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5505\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5505\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5498\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5498\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5498\
        );

    \I__1147\ : Span4Mux_h
    port map (
            O => \N__5529\,
            I => \N__5493\
        );

    \I__1146\ : Span4Mux_h
    port map (
            O => \N__5526\,
            I => \N__5493\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5490\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5481\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5481\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5481\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5481\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5472\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5472\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5472\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5472\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5510\,
            I => state_3
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5505\,
            I => state_3
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5498\,
            I => state_3
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__5493\,
            I => state_3
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5490\,
            I => state_3
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5481\,
            I => state_3
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5472\,
            I => state_3
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__5457\,
            I => \N__5453\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5450\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5447\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5450\,
            I => \N__5442\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5442\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__5442\,
            I => n1826
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5439\,
            I => \N__5436\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5433\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5433\,
            I => n314
        );

    \I__1120\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5426\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5423\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5426\,
            I => n1817
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5423\,
            I => n1817
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__5418\,
            I => \eeprom.i2c.n12_cascade_\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5406\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5406\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5406\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5406\,
            I => n4_adj_408
        );

    \I__1111\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5400\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5400\,
            I => \eeprom.i2c.n942\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5397\,
            I => \N__5393\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5389\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5386\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5383\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5389\,
            I => \N__5380\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5386\,
            I => n10_adj_398
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5383\,
            I => n10_adj_398
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__5380\,
            I => n10_adj_398
        );

    \I__1101\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5369\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5366\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5363\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5366\,
            I => n11_adj_400
        );

    \I__1097\ : Odrv4
    port map (
            O => \N__5363\,
            I => n11_adj_400
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__5358\,
            I => \eeprom.i2c.n942_cascade_\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5351\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5348\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5351\,
            I => n1532
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__5348\,
            I => n1532
        );

    \I__1091\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5337\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5337\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5331\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5328\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5325\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5322\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__5331\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5328\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5325\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5322\,
            I => \eeprom.i2c.counter_0\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5313\,
            I => \bfn_21_22_0_\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5310\,
            I => \eeprom.i2c.n2256\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5307\,
            I => \eeprom.i2c.n2257\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5300\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5300\,
            I => \eeprom.i2c.counter_3\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5297\,
            I => \eeprom.i2c.counter_3\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5292\,
            I => \eeprom.i2c.n2258\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__5289\,
            I => \N__5285\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__5288\,
            I => \N__5282\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5279\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5276\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5279\,
            I => \eeprom.i2c.counter_4\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5276\,
            I => \eeprom.i2c.counter_4\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5271\,
            I => \eeprom.i2c.n2259\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__5268\,
            I => \n10_adj_398_cascade_\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5261\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5258\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5261\,
            I => \state_7_N_269_0\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5258\,
            I => \state_7_N_269_0\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__5253\,
            I => \n2460_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__5244\,
            I => n2560
        );

    \I__1057\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5238\,
            I => n308
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5229\,
            I => n320
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5220\,
            I => n318
        );

    \I__1049\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5214\,
            I => \eeprom.i2c.n9\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5207\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5204\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5207\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5204\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5199\,
            I => \bfn_21_18_0_\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5192\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5189\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5192\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5189\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5184\,
            I => \eeprom.i2c.n2319\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5177\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5174\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5177\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5174\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5169\,
            I => \eeprom.i2c.n2320\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5162\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5159\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5162\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5159\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5154\,
            I => \eeprom.i2c.n2321\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5151\,
            I => \eeprom.i2c.n2322\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5144\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5141\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5144\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5141\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__1022\ : ClkMux
    port map (
            O => \N__5136\,
            I => \N__5076\
        );

    \I__1021\ : ClkMux
    port map (
            O => \N__5135\,
            I => \N__5076\
        );

    \I__1020\ : ClkMux
    port map (
            O => \N__5134\,
            I => \N__5076\
        );

    \I__1019\ : ClkMux
    port map (
            O => \N__5133\,
            I => \N__5076\
        );

    \I__1018\ : ClkMux
    port map (
            O => \N__5132\,
            I => \N__5076\
        );

    \I__1017\ : ClkMux
    port map (
            O => \N__5131\,
            I => \N__5076\
        );

    \I__1016\ : ClkMux
    port map (
            O => \N__5130\,
            I => \N__5076\
        );

    \I__1015\ : ClkMux
    port map (
            O => \N__5129\,
            I => \N__5076\
        );

    \I__1014\ : ClkMux
    port map (
            O => \N__5128\,
            I => \N__5076\
        );

    \I__1013\ : ClkMux
    port map (
            O => \N__5127\,
            I => \N__5076\
        );

    \I__1012\ : ClkMux
    port map (
            O => \N__5126\,
            I => \N__5076\
        );

    \I__1011\ : ClkMux
    port map (
            O => \N__5125\,
            I => \N__5076\
        );

    \I__1010\ : ClkMux
    port map (
            O => \N__5124\,
            I => \N__5076\
        );

    \I__1009\ : ClkMux
    port map (
            O => \N__5123\,
            I => \N__5076\
        );

    \I__1008\ : ClkMux
    port map (
            O => \N__5122\,
            I => \N__5076\
        );

    \I__1007\ : ClkMux
    port map (
            O => \N__5121\,
            I => \N__5076\
        );

    \I__1006\ : ClkMux
    port map (
            O => \N__5120\,
            I => \N__5076\
        );

    \I__1005\ : ClkMux
    port map (
            O => \N__5119\,
            I => \N__5076\
        );

    \I__1004\ : ClkMux
    port map (
            O => \N__5118\,
            I => \N__5076\
        );

    \I__1003\ : ClkMux
    port map (
            O => \N__5117\,
            I => \N__5076\
        );

    \I__1002\ : GlobalMux
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__1001\ : gio2CtrlBuf
    port map (
            O => \N__5073\,
            I => \CLK_N\
        );

    \I__1000\ : SRMux
    port map (
            O => \N__5070\,
            I => \N__5067\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5062\
        );

    \I__998\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5059\
        );

    \I__997\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5056\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__5062\,
            I => \eeprom.i2c.counter2_7__N_256\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5059\,
            I => \eeprom.i2c.counter2_7__N_256\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5056\,
            I => \eeprom.i2c.counter2_7__N_256\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__992\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5043\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5043\,
            I => n306
        );

    \I__990\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5035\
        );

    \I__989\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5030\
        );

    \I__988\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5030\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5035\,
            I => saved_addr_0
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5030\,
            I => saved_addr_0
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__984\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5018\
        );

    \I__983\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5015\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5018\,
            I => n11_adj_399
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5015\,
            I => n11_adj_399
        );

    \I__980\ : InMux
    port map (
            O => \N__5010\,
            I => \N__5007\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5007\,
            I => n2566
        );

    \I__978\ : InMux
    port map (
            O => \N__5004\,
            I => \N__5001\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5001\,
            I => \eeprom.i2c.n39\
        );

    \I__976\ : CEMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__974\ : Span4Mux_v
    port map (
            O => \N__4992\,
            I => \N__4989\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__4989\,
            I => \eeprom.i2c.n2406\
        );

    \I__972\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4982\
        );

    \I__971\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4979\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4979\,
            I => \eeprom.i2c.n37\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__4976\,
            I => \eeprom.i2c.n37\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__4971\,
            I => \eeprom.i2c.n1051_cascade_\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__965\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4962\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4962\,
            I => \eeprom.i2c.n13\
        );

    \I__963\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4954\
        );

    \I__962\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4951\
        );

    \I__961\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4948\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4954\,
            I => sda_out
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4951\,
            I => sda_out
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4948\,
            I => sda_out
        );

    \I__957\ : IoInMux
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__955\ : Span4Mux_s1_h
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__954\ : Sp12to4
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__953\ : Span12Mux_v
    port map (
            O => \N__4929\,
            I => \N__4925\
        );

    \I__952\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4920\
        );

    \I__951\ : Span12Mux_h
    port map (
            O => \N__4925\,
            I => \N__4917\
        );

    \I__950\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4914\
        );

    \I__949\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4911\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4908\
        );

    \I__947\ : Odrv12
    port map (
            O => \N__4917\,
            I => sda_enable
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4914\,
            I => sda_enable
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4911\,
            I => sda_enable
        );

    \I__944\ : Odrv4
    port map (
            O => \N__4908\,
            I => sda_enable
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__4899\,
            I => \state_7_N_285_3_cascade_\
        );

    \I__942\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4893\,
            I => \eeprom.i2c.n2475\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__4890\,
            I => \eeprom.i2c.n2475_cascade_\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__4887\,
            I => \n949_cascade_\
        );

    \I__938\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4880\
        );

    \I__937\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4877\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4880\,
            I => n949
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4877\,
            I => n949
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__4872\,
            I => \n2547_cascade_\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__4869\,
            I => \eeprom.i2c.n2574_cascade_\
        );

    \I__932\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4863\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4863\,
            I => \eeprom.i2c.n2557\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__4860\,
            I => \N__4857\
        );

    \I__929\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4853\
        );

    \I__928\ : SRMux
    port map (
            O => \N__4856\,
            I => \N__4850\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4853\,
            I => \N__4846\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4850\,
            I => \N__4843\
        );

    \I__925\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4840\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__4846\,
            I => \N__4837\
        );

    \I__923\ : Span4Mux_h
    port map (
            O => \N__4843\,
            I => \N__4834\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4840\,
            I => \N__4831\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__4837\,
            I => \eeprom.enable\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__4834\,
            I => \eeprom.enable\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__4831\,
            I => \eeprom.enable\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__4824\,
            I => \n2538_cascade_\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__4821\,
            I => \n4_adj_411_cascade_\
        );

    \I__916\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4815\,
            I => n1835
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__4812\,
            I => \n2507_cascade_\
        );

    \I__913\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4806\,
            I => n10_adj_394
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__4803\,
            I => \N__4800\
        );

    \I__910\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4795\
        );

    \I__909\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4792\
        );

    \I__908\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4789\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4795\,
            I => \eeprom.i2c.n11_adj_379\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4792\,
            I => \eeprom.i2c.n11_adj_379\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4789\,
            I => \eeprom.i2c.n11_adj_379\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__4782\,
            I => \eeprom.i2c.n6_cascade_\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__4779\,
            I => \eeprom.i2c.counter2_7__N_256_cascade_\
        );

    \I__902\ : CEMux
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4773\,
            I => \eeprom.i2c.n1580\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__899\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4764\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4764\,
            I => \N__4760\
        );

    \I__897\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4757\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__4760\,
            I => rw
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4757\,
            I => rw
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__4752\,
            I => \n1835_cascade_\
        );

    \I__893\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4746\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4746\,
            I => n2569
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__4743\,
            I => \n11_adj_399_cascade_\
        );

    \I__890\ : SRMux
    port map (
            O => \N__4740\,
            I => \N__4737\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4737\,
            I => \eeprom.i2c.n1669\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__4734\,
            I => \eeprom.i2c.n37_cascade_\
        );

    \I__887\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4725\
        );

    \I__886\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4725\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4725\,
            I => \eeprom.i2c.n33\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__4722\,
            I => \eeprom.i2c.n39_cascade_\
        );

    \I__883\ : CEMux
    port map (
            O => \N__4719\,
            I => \N__4716\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__4713\,
            I => \eeprom.i2c.n1027\
        );

    \I__880\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4707\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4707\,
            I => \eeprom.delay_counter_15_N_171_3\
        );

    \I__878\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4701\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4701\,
            I => \N__4696\
        );

    \I__876\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4693\
        );

    \I__875\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4690\
        );

    \I__874\ : Span4Mux_v
    port map (
            O => \N__4696\,
            I => \N__4687\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4693\,
            I => \eeprom.delay_counter_3\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4690\,
            I => \eeprom.delay_counter_3\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__4687\,
            I => \eeprom.delay_counter_3\
        );

    \I__870\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4677\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4677\,
            I => \eeprom.delay_counter_15_N_171_11\
        );

    \I__868\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4671\,
            I => \eeprom.delay_counter_15_N_171_9\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__865\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4660\
        );

    \I__864\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4655\
        );

    \I__863\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4655\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4660\,
            I => \eeprom.delay_counter_11\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4655\,
            I => \eeprom.delay_counter_11\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__4650\,
            I => \N__4646\
        );

    \I__859\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4643\
        );

    \I__858\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4639\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4643\,
            I => \N__4636\
        );

    \I__856\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4633\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4639\,
            I => \eeprom.delay_counter_7\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__4636\,
            I => \eeprom.delay_counter_7\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4633\,
            I => \eeprom.delay_counter_7\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__4626\,
            I => \eeprom.n6_cascade_\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \N__4619\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__4622\,
            I => \N__4616\
        );

    \I__849\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4613\
        );

    \I__848\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4610\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4613\,
            I => \N__4604\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4604\
        );

    \I__845\ : InMux
    port map (
            O => \N__4609\,
            I => \N__4601\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__4604\,
            I => \eeprom.delay_counter_9\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4601\,
            I => \eeprom.delay_counter_9\
        );

    \I__842\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4593\,
            I => \eeprom.n8\
        );

    \I__840\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4587\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4587\,
            I => \eeprom.delay_counter_15_N_171_15\
        );

    \I__838\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4579\
        );

    \I__837\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4574\
        );

    \I__836\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4574\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4579\,
            I => \eeprom.delay_counter_15\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4574\,
            I => \eeprom.delay_counter_15\
        );

    \I__833\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4566\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4566\,
            I => \eeprom.delay_counter_15_N_171_14\
        );

    \I__831\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4558\
        );

    \I__830\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4553\
        );

    \I__829\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4553\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4558\,
            I => \eeprom.delay_counter_14\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4553\,
            I => \eeprom.delay_counter_14\
        );

    \I__826\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4535\
        );

    \I__825\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4532\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4546\,
            I => \N__4525\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__4545\,
            I => \N__4522\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4544\,
            I => \N__4519\
        );

    \I__821\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4507\
        );

    \I__820\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4507\
        );

    \I__819\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4507\
        );

    \I__818\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4507\
        );

    \I__817\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4504\
        );

    \I__816\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4501\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4535\,
            I => \N__4496\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4496\
        );

    \I__813\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4491\
        );

    \I__812\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4491\
        );

    \I__811\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4486\
        );

    \I__810\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4486\
        );

    \I__809\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4475\
        );

    \I__808\ : InMux
    port map (
            O => \N__4522\,
            I => \N__4475\
        );

    \I__807\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4475\
        );

    \I__806\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4475\
        );

    \I__805\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4475\
        );

    \I__804\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4464\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4507\,
            I => \N__4461\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4458\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4501\,
            I => \N__4451\
        );

    \I__800\ : Span4Mux_h
    port map (
            O => \N__4496\,
            I => \N__4451\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4491\,
            I => \N__4451\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4486\,
            I => \N__4446\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4475\,
            I => \N__4446\
        );

    \I__796\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4439\
        );

    \I__795\ : InMux
    port map (
            O => \N__4473\,
            I => \N__4439\
        );

    \I__794\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4439\
        );

    \I__793\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4428\
        );

    \I__792\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4428\
        );

    \I__791\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4428\
        );

    \I__790\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4428\
        );

    \I__789\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4428\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4464\,
            I => state_0
        );

    \I__787\ : Odrv4
    port map (
            O => \N__4461\,
            I => state_0
        );

    \I__786\ : Odrv4
    port map (
            O => \N__4458\,
            I => state_0
        );

    \I__785\ : Odrv4
    port map (
            O => \N__4451\,
            I => state_0
        );

    \I__784\ : Odrv4
    port map (
            O => \N__4446\,
            I => state_0
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4439\,
            I => state_0
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4428\,
            I => state_0
        );

    \I__781\ : CascadeMux
    port map (
            O => \N__4413\,
            I => \N__4405\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__4412\,
            I => \N__4401\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__4411\,
            I => \N__4398\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__4410\,
            I => \N__4395\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__4409\,
            I => \N__4392\
        );

    \I__776\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4387\
        );

    \I__775\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4387\
        );

    \I__774\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4384\
        );

    \I__773\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4377\
        );

    \I__772\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4377\
        );

    \I__771\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4377\
        );

    \I__770\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4374\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4387\,
            I => \N__4367\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4384\,
            I => \N__4362\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4377\,
            I => \N__4362\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4374\,
            I => \N__4359\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__4373\,
            I => \N__4353\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__4372\,
            I => \N__4350\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__4371\,
            I => \N__4346\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__4370\,
            I => \N__4343\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__4367\,
            I => \N__4339\
        );

    \I__760\ : Span4Mux_h
    port map (
            O => \N__4362\,
            I => \N__4336\
        );

    \I__759\ : Span4Mux_h
    port map (
            O => \N__4359\,
            I => \N__4333\
        );

    \I__758\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4322\
        );

    \I__757\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4322\
        );

    \I__756\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4322\
        );

    \I__755\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4322\
        );

    \I__754\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4322\
        );

    \I__753\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4319\
        );

    \I__752\ : InMux
    port map (
            O => \N__4346\,
            I => \N__4312\
        );

    \I__751\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4312\
        );

    \I__750\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4312\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__4339\,
            I => \eeprom.n1601\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__4336\,
            I => \eeprom.n1601\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__4333\,
            I => \eeprom.n1601\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4322\,
            I => \eeprom.n1601\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4319\,
            I => \eeprom.n1601\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4312\,
            I => \eeprom.n1601\
        );

    \I__743\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4296\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4296\,
            I => \eeprom.delay_counter_15_N_171_13\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__4293\,
            I => \N__4289\
        );

    \I__740\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4285\
        );

    \I__739\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4282\
        );

    \I__738\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4279\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4285\,
            I => \eeprom.delay_counter_13\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4282\,
            I => \eeprom.delay_counter_13\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4279\,
            I => \eeprom.delay_counter_13\
        );

    \I__734\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4268\
        );

    \I__733\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4265\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4268\,
            I => \N__4262\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4265\,
            I => delay_counter_5
        );

    \I__730\ : Odrv4
    port map (
            O => \N__4262\,
            I => delay_counter_5
        );

    \I__729\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4254\,
            I => n16_adj_407
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__4251\,
            I => \N__4248\
        );

    \I__726\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4244\
        );

    \I__725\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4241\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4244\,
            I => \N__4238\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4241\,
            I => delay_counter_2
        );

    \I__722\ : Odrv4
    port map (
            O => \N__4238\,
            I => delay_counter_2
        );

    \I__721\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4230\,
            I => n17_adj_406
        );

    \I__719\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4224\,
            I => n2536
        );

    \I__717\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4215\
        );

    \I__716\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4210\
        );

    \I__715\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4210\
        );

    \I__714\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4207\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4215\,
            I => \N__4204\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4201\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4198\
        );

    \I__710\ : Span4Mux_v
    port map (
            O => \N__4204\,
            I => \N__4193\
        );

    \I__709\ : Span4Mux_h
    port map (
            O => \N__4201\,
            I => \N__4193\
        );

    \I__708\ : Odrv4
    port map (
            O => \N__4198\,
            I => \read_N\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__4193\,
            I => \read_N\
        );

    \I__706\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4184\
        );

    \I__705\ : InMux
    port map (
            O => \N__4187\,
            I => \N__4181\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__4184\,
            I => delay_counter_22
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4181\,
            I => delay_counter_22
        );

    \I__702\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4172\
        );

    \I__701\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4169\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4172\,
            I => delay_counter_25
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4169\,
            I => delay_counter_25
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__4164\,
            I => \N__4160\
        );

    \I__697\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4157\
        );

    \I__696\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4154\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4157\,
            I => delay_counter_20
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4154\,
            I => delay_counter_20
        );

    \I__693\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4146\,
            I => n8_adj_412
        );

    \I__691\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4140\,
            I => n9_adj_404
        );

    \I__689\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4130\
        );

    \I__688\ : InMux
    port map (
            O => \N__4136\,
            I => \N__4130\
        );

    \I__687\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4127\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4130\,
            I => \N__4124\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4127\,
            I => delay_counter_31
        );

    \I__684\ : Odrv4
    port map (
            O => \N__4124\,
            I => delay_counter_31
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__4119\,
            I => \n9_adj_404_cascade_\
        );

    \I__682\ : SRMux
    port map (
            O => \N__4116\,
            I => \N__4113\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4113\,
            I => \N__4108\
        );

    \I__680\ : SRMux
    port map (
            O => \N__4112\,
            I => \N__4105\
        );

    \I__679\ : SRMux
    port map (
            O => \N__4111\,
            I => \N__4102\
        );

    \I__678\ : Span4Mux_v
    port map (
            O => \N__4108\,
            I => \N__4096\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4105\,
            I => \N__4096\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4102\,
            I => \N__4093\
        );

    \I__675\ : SRMux
    port map (
            O => \N__4101\,
            I => \N__4090\
        );

    \I__674\ : Span4Mux_h
    port map (
            O => \N__4096\,
            I => \N__4087\
        );

    \I__673\ : Span4Mux_h
    port map (
            O => \N__4093\,
            I => \N__4084\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4090\,
            I => \N__4081\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__4087\,
            I => \addr_10__N_70\
        );

    \I__670\ : Odrv4
    port map (
            O => \N__4084\,
            I => \addr_10__N_70\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__4081\,
            I => \addr_10__N_70\
        );

    \I__668\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4070\
        );

    \I__667\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4067\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4070\,
            I => delay_counter_29
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4067\,
            I => delay_counter_29
        );

    \I__664\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4058\
        );

    \I__663\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4055\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4058\,
            I => delay_counter_28
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4055\,
            I => delay_counter_28
        );

    \I__660\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4044\
        );

    \I__659\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4044\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__4041\,
            I => n10_adj_403
        );

    \I__656\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4034\
        );

    \I__655\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4031\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4034\,
            I => delay_counter_26
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4031\,
            I => delay_counter_26
        );

    \I__652\ : InMux
    port map (
            O => \N__4026\,
            I => \N__4022\
        );

    \I__651\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4019\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4022\,
            I => delay_counter_30
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4019\,
            I => delay_counter_30
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__4014\,
            I => \N__4010\
        );

    \I__647\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4007\
        );

    \I__646\ : InMux
    port map (
            O => \N__4010\,
            I => \N__4004\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4007\,
            I => delay_counter_27
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4004\,
            I => delay_counter_27
        );

    \I__643\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3995\
        );

    \I__642\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3992\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3995\,
            I => delay_counter_24
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3992\,
            I => delay_counter_24
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__638\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3980\
        );

    \I__637\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3977\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3974\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3977\,
            I => \N__3971\
        );

    \I__634\ : Odrv4
    port map (
            O => \N__3974\,
            I => n14_adj_401
        );

    \I__633\ : Odrv4
    port map (
            O => \N__3971\,
            I => n14_adj_401
        );

    \I__632\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3963\,
            I => \eeprom.delay_counter_15_N_171_7\
        );

    \I__630\ : SRMux
    port map (
            O => \N__3960\,
            I => \N__3957\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__628\ : Span4Mux_h
    port map (
            O => \N__3954\,
            I => \N__3944\
        );

    \I__627\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3941\
        );

    \I__626\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3936\
        );

    \I__625\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3936\
        );

    \I__624\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3927\
        );

    \I__623\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3927\
        );

    \I__622\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3927\
        );

    \I__621\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3927\
        );

    \I__620\ : Odrv4
    port map (
            O => \N__3944\,
            I => state_1
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3941\,
            I => state_1
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3936\,
            I => state_1
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3927\,
            I => state_1
        );

    \I__616\ : CEMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__614\ : Odrv12
    port map (
            O => \N__3912\,
            I => n1568
        );

    \I__613\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3905\
        );

    \I__612\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3902\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3905\,
            I => delay_counter_7
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3902\,
            I => delay_counter_7
        );

    \I__609\ : InMux
    port map (
            O => \N__3897\,
            I => \N__3893\
        );

    \I__608\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3890\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3893\,
            I => delay_counter_8
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3890\,
            I => delay_counter_8
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__3885\,
            I => \N__3881\
        );

    \I__604\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3878\
        );

    \I__603\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3875\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3878\,
            I => delay_counter_1
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3875\,
            I => delay_counter_1
        );

    \I__600\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3866\
        );

    \I__599\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3863\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3866\,
            I => delay_counter_4
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3863\,
            I => delay_counter_4
        );

    \I__596\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3854\
        );

    \I__595\ : InMux
    port map (
            O => \N__3857\,
            I => \N__3851\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3854\,
            I => delay_counter_10
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3851\,
            I => delay_counter_10
        );

    \I__592\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3842\
        );

    \I__591\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3839\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3842\,
            I => delay_counter_12
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3839\,
            I => delay_counter_12
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3834\,
            I => \N__3830\
        );

    \I__587\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3827\
        );

    \I__586\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3824\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3827\,
            I => delay_counter_11
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3824\,
            I => delay_counter_11
        );

    \I__583\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3815\
        );

    \I__582\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3812\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3815\,
            I => delay_counter_13
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3812\,
            I => delay_counter_13
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__3807\,
            I => \n2512_cascade_\
        );

    \I__578\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3800\
        );

    \I__577\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3797\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3800\,
            I => delay_counter_16
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3797\,
            I => delay_counter_16
        );

    \I__574\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3788\
        );

    \I__573\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3785\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3788\,
            I => delay_counter_18
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3785\,
            I => delay_counter_18
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__3780\,
            I => \n2495_cascade_\
        );

    \I__569\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3773\
        );

    \I__568\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3770\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3773\,
            I => delay_counter_19
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3770\,
            I => delay_counter_19
        );

    \I__565\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3761\
        );

    \I__564\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3758\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3761\,
            I => delay_counter_9
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3758\,
            I => delay_counter_9
        );

    \I__561\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3749\
        );

    \I__560\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3746\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3749\,
            I => delay_counter_6
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3746\,
            I => delay_counter_6
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__3741\,
            I => \N__3737\
        );

    \I__556\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3734\
        );

    \I__555\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3731\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3734\,
            I => delay_counter_3
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3731\,
            I => delay_counter_3
        );

    \I__552\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3722\
        );

    \I__551\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3719\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3722\,
            I => delay_counter_0
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3719\,
            I => delay_counter_0
        );

    \I__548\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3710\
        );

    \I__547\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3707\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3710\,
            I => delay_counter_17
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3707\,
            I => delay_counter_17
        );

    \I__544\ : InMux
    port map (
            O => \N__3702\,
            I => \N__3698\
        );

    \I__543\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3695\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3698\,
            I => delay_counter_15
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3695\,
            I => delay_counter_15
        );

    \I__540\ : InMux
    port map (
            O => \N__3690\,
            I => \N__3686\
        );

    \I__539\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3683\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3686\,
            I => delay_counter_14
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3683\,
            I => delay_counter_14
        );

    \I__536\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3675\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3675\,
            I => n8
        );

    \I__534\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3668\
        );

    \I__533\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3665\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3668\,
            I => delay_counter_21
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3665\,
            I => delay_counter_21
        );

    \I__530\ : InMux
    port map (
            O => \N__3660\,
            I => \N__3656\
        );

    \I__529\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3653\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3656\,
            I => delay_counter_23
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3653\,
            I => delay_counter_23
        );

    \I__526\ : InMux
    port map (
            O => \N__3648\,
            I => \N__3645\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3645\,
            I => n6_adj_413
        );

    \I__524\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3639\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3639\,
            I => \N__3636\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__3636\,
            I => \eeprom.delay_counter_15_N_171_4\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__3633\,
            I => \N__3630\
        );

    \I__520\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3627\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3627\,
            I => \N__3622\
        );

    \I__518\ : InMux
    port map (
            O => \N__3626\,
            I => \N__3617\
        );

    \I__517\ : InMux
    port map (
            O => \N__3625\,
            I => \N__3617\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__3622\,
            I => \eeprom.delay_counter_4\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3617\,
            I => \eeprom.delay_counter_4\
        );

    \I__514\ : InMux
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3609\,
            I => n324
        );

    \I__512\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3600\
        );

    \I__511\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3597\
        );

    \I__510\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3592\
        );

    \I__509\ : InMux
    port map (
            O => \N__3603\,
            I => \N__3592\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3600\,
            I => \eeprom.n1500\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3597\,
            I => \eeprom.n1500\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3592\,
            I => \eeprom.n1500\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__3585\,
            I => \n6_adj_405_cascade_\
        );

    \I__504\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3579\,
            I => n41
        );

    \I__502\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3573\,
            I => \eeprom.n1018\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__3570\,
            I => \n2483_cascade_\
        );

    \I__499\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3564\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3564\,
            I => \eeprom.n2453\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3561\,
            I => \n1568_cascade_\
        );

    \I__496\ : InMux
    port map (
            O => \N__3558\,
            I => \eeprom.n2254\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__3555\,
            I => \N__3544\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__3554\,
            I => \N__3540\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__3553\,
            I => \N__3536\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__3552\,
            I => \N__3532\
        );

    \I__491\ : CascadeMux
    port map (
            O => \N__3551\,
            I => \N__3529\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3550\,
            I => \N__3525\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__3549\,
            I => \N__3521\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3548\,
            I => \N__3517\
        );

    \I__487\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3499\
        );

    \I__486\ : InMux
    port map (
            O => \N__3544\,
            I => \N__3499\
        );

    \I__485\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3499\
        );

    \I__484\ : InMux
    port map (
            O => \N__3540\,
            I => \N__3499\
        );

    \I__483\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3499\
        );

    \I__482\ : InMux
    port map (
            O => \N__3536\,
            I => \N__3499\
        );

    \I__481\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3499\
        );

    \I__480\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3499\
        );

    \I__479\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3482\
        );

    \I__478\ : InMux
    port map (
            O => \N__3528\,
            I => \N__3482\
        );

    \I__477\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3482\
        );

    \I__476\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3482\
        );

    \I__475\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3482\
        );

    \I__474\ : InMux
    port map (
            O => \N__3520\,
            I => \N__3482\
        );

    \I__473\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3482\
        );

    \I__472\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3482\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3499\,
            I => \eeprom.n642\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3482\,
            I => \eeprom.n642\
        );

    \I__469\ : InMux
    port map (
            O => \N__3477\,
            I => \eeprom.n2255\
        );

    \I__468\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3471\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3471\,
            I => \eeprom.n14\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__3468\,
            I => \eeprom.n13_cascade_\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__3465\,
            I => \eeprom.n7_cascade_\
        );

    \I__464\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3459\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3459\,
            I => \N__3456\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__3456\,
            I => \eeprom.delay_counter_15_N_171_1\
        );

    \I__461\ : InMux
    port map (
            O => \N__3453\,
            I => \N__3450\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3450\,
            I => \N__3445\
        );

    \I__459\ : InMux
    port map (
            O => \N__3449\,
            I => \N__3440\
        );

    \I__458\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3440\
        );

    \I__457\ : Odrv4
    port map (
            O => \N__3445\,
            I => \eeprom.delay_counter_1\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3440\,
            I => \eeprom.delay_counter_1\
        );

    \I__455\ : InMux
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3432\,
            I => \N__3429\
        );

    \I__453\ : Odrv4
    port map (
            O => \N__3429\,
            I => \eeprom.delay_counter_15_N_171_0\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__3426\,
            I => \N__3423\
        );

    \I__451\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3420\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3415\
        );

    \I__449\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3410\
        );

    \I__448\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3410\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__3415\,
            I => \eeprom.delay_counter_0\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3410\,
            I => \eeprom.delay_counter_0\
        );

    \I__445\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3402\,
            I => \N__3399\
        );

    \I__443\ : Odrv4
    port map (
            O => \N__3399\,
            I => \eeprom.delay_counter_15_N_171_5\
        );

    \I__442\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3393\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3393\,
            I => \N__3388\
        );

    \I__440\ : InMux
    port map (
            O => \N__3392\,
            I => \N__3383\
        );

    \I__439\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3383\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__3388\,
            I => \eeprom.delay_counter_5\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3383\,
            I => \eeprom.delay_counter_5\
        );

    \I__436\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3375\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3375\,
            I => \eeprom.delay_counter_15_N_171_10\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__3372\,
            I => \N__3367\
        );

    \I__433\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3364\
        );

    \I__432\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3359\
        );

    \I__431\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3359\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3364\,
            I => \eeprom.delay_counter_10\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3359\,
            I => \eeprom.delay_counter_10\
        );

    \I__428\ : InMux
    port map (
            O => \N__3354\,
            I => \eeprom.n2245\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__3351\,
            I => \N__3348\
        );

    \I__426\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3344\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3347\,
            I => \N__3340\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3344\,
            I => \N__3337\
        );

    \I__423\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3332\
        );

    \I__422\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3332\
        );

    \I__421\ : Odrv4
    port map (
            O => \N__3337\,
            I => \eeprom.delay_counter_6\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3332\,
            I => \eeprom.delay_counter_6\
        );

    \I__419\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__3321\,
            I => \eeprom.delay_counter_15_N_171_6\
        );

    \I__416\ : InMux
    port map (
            O => \N__3318\,
            I => \eeprom.n2246\
        );

    \I__415\ : InMux
    port map (
            O => \N__3315\,
            I => \eeprom.n2247\
        );

    \I__414\ : InMux
    port map (
            O => \N__3312\,
            I => \N__3307\
        );

    \I__413\ : InMux
    port map (
            O => \N__3311\,
            I => \N__3302\
        );

    \I__412\ : InMux
    port map (
            O => \N__3310\,
            I => \N__3302\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3307\,
            I => \eeprom.delay_counter_8\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3302\,
            I => \eeprom.delay_counter_8\
        );

    \I__409\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3294\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3294\,
            I => \eeprom.delay_counter_15_N_171_8\
        );

    \I__407\ : InMux
    port map (
            O => \N__3291\,
            I => \bfn_18_18_0_\
        );

    \I__406\ : InMux
    port map (
            O => \N__3288\,
            I => \eeprom.n2249\
        );

    \I__405\ : InMux
    port map (
            O => \N__3285\,
            I => \eeprom.n2250\
        );

    \I__404\ : InMux
    port map (
            O => \N__3282\,
            I => \eeprom.n2251\
        );

    \I__403\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3274\
        );

    \I__402\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3269\
        );

    \I__401\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3269\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3274\,
            I => \eeprom.delay_counter_12\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3269\,
            I => \eeprom.delay_counter_12\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__3264\,
            I => \N__3261\
        );

    \I__397\ : InMux
    port map (
            O => \N__3261\,
            I => \N__3258\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3258\,
            I => \eeprom.delay_counter_15_N_171_12\
        );

    \I__395\ : InMux
    port map (
            O => \N__3255\,
            I => \eeprom.n2252\
        );

    \I__394\ : InMux
    port map (
            O => \N__3252\,
            I => \eeprom.n2253\
        );

    \I__393\ : InMux
    port map (
            O => \N__3249\,
            I => n2290
        );

    \I__392\ : InMux
    port map (
            O => \N__3246\,
            I => n2291
        );

    \I__391\ : InMux
    port map (
            O => \N__3243\,
            I => n2292
        );

    \I__390\ : InMux
    port map (
            O => \N__3240\,
            I => n2293
        );

    \I__389\ : InMux
    port map (
            O => \N__3237\,
            I => \eeprom.n2241\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__3234\,
            I => \N__3231\
        );

    \I__387\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3228\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3228\,
            I => \N__3223\
        );

    \I__385\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3218\
        );

    \I__384\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3218\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__3223\,
            I => \eeprom.delay_counter_2\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3218\,
            I => \eeprom.delay_counter_2\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__3213\,
            I => \N__3210\
        );

    \I__380\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3207\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3207\,
            I => \N__3204\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__3204\,
            I => \eeprom.delay_counter_15_N_171_2\
        );

    \I__377\ : InMux
    port map (
            O => \N__3201\,
            I => \eeprom.n2242\
        );

    \I__376\ : InMux
    port map (
            O => \N__3198\,
            I => \eeprom.n2243\
        );

    \I__375\ : InMux
    port map (
            O => \N__3195\,
            I => \eeprom.n2244\
        );

    \I__374\ : InMux
    port map (
            O => \N__3192\,
            I => n2281
        );

    \I__373\ : InMux
    port map (
            O => \N__3189\,
            I => n2282
        );

    \I__372\ : InMux
    port map (
            O => \N__3186\,
            I => n2283
        );

    \I__371\ : InMux
    port map (
            O => \N__3183\,
            I => n2284
        );

    \I__370\ : InMux
    port map (
            O => \N__3180\,
            I => n2285
        );

    \I__369\ : InMux
    port map (
            O => \N__3177\,
            I => \bfn_17_24_0_\
        );

    \I__368\ : InMux
    port map (
            O => \N__3174\,
            I => n2287
        );

    \I__367\ : InMux
    port map (
            O => \N__3171\,
            I => n2288
        );

    \I__366\ : InMux
    port map (
            O => \N__3168\,
            I => n2289
        );

    \I__365\ : InMux
    port map (
            O => \N__3165\,
            I => n2272
        );

    \I__364\ : InMux
    port map (
            O => \N__3162\,
            I => n2273
        );

    \I__363\ : InMux
    port map (
            O => \N__3159\,
            I => n2274
        );

    \I__362\ : InMux
    port map (
            O => \N__3156\,
            I => n2275
        );

    \I__361\ : InMux
    port map (
            O => \N__3153\,
            I => n2276
        );

    \I__360\ : InMux
    port map (
            O => \N__3150\,
            I => n2277
        );

    \I__359\ : InMux
    port map (
            O => \N__3147\,
            I => \bfn_17_23_0_\
        );

    \I__358\ : InMux
    port map (
            O => \N__3144\,
            I => n2279
        );

    \I__357\ : InMux
    port map (
            O => \N__3141\,
            I => n2280
        );

    \I__356\ : InMux
    port map (
            O => \N__3138\,
            I => n2263
        );

    \I__355\ : InMux
    port map (
            O => \N__3135\,
            I => n2264
        );

    \I__354\ : InMux
    port map (
            O => \N__3132\,
            I => n2265
        );

    \I__353\ : InMux
    port map (
            O => \N__3129\,
            I => n2266
        );

    \I__352\ : InMux
    port map (
            O => \N__3126\,
            I => n2267
        );

    \I__351\ : InMux
    port map (
            O => \N__3123\,
            I => n2268
        );

    \I__350\ : InMux
    port map (
            O => \N__3120\,
            I => n2269
        );

    \I__349\ : InMux
    port map (
            O => \N__3117\,
            I => \bfn_17_22_0_\
        );

    \I__348\ : InMux
    port map (
            O => \N__3114\,
            I => n2271
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__3111\,
            I => \n693_cascade_\
        );

    \I__346\ : InMux
    port map (
            O => \N__3108\,
            I => \bfn_17_21_0_\
        );

    \I__345\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3102\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3102\,
            I => n7
        );

    \I__343\ : InMux
    port map (
            O => \N__3099\,
            I => n2312
        );

    \I__342\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3093\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3093\,
            I => n6_adj_410
        );

    \I__340\ : InMux
    port map (
            O => \N__3090\,
            I => n2313
        );

    \I__339\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3080\
        );

    \I__338\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3080\
        );

    \I__337\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3077\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3080\,
            I => blink_counter_21
        );

    \I__335\ : LocalMux
    port map (
            O => \N__3077\,
            I => blink_counter_21
        );

    \I__334\ : InMux
    port map (
            O => \N__3072\,
            I => n2314
        );

    \I__333\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3062\
        );

    \I__332\ : InMux
    port map (
            O => \N__3068\,
            I => \N__3062\
        );

    \I__331\ : InMux
    port map (
            O => \N__3067\,
            I => \N__3059\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3062\,
            I => blink_counter_22
        );

    \I__329\ : LocalMux
    port map (
            O => \N__3059\,
            I => blink_counter_22
        );

    \I__328\ : InMux
    port map (
            O => \N__3054\,
            I => n2315
        );

    \I__327\ : CascadeMux
    port map (
            O => \N__3051\,
            I => \N__3047\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__3050\,
            I => \N__3044\
        );

    \I__325\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3038\
        );

    \I__324\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3038\
        );

    \I__323\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3035\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3038\,
            I => blink_counter_23
        );

    \I__321\ : LocalMux
    port map (
            O => \N__3035\,
            I => blink_counter_23
        );

    \I__320\ : InMux
    port map (
            O => \N__3030\,
            I => n2316
        );

    \I__319\ : InMux
    port map (
            O => \N__3027\,
            I => \N__3020\
        );

    \I__318\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3020\
        );

    \I__317\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3017\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3020\,
            I => blink_counter_24
        );

    \I__315\ : LocalMux
    port map (
            O => \N__3017\,
            I => blink_counter_24
        );

    \I__314\ : InMux
    port map (
            O => \N__3012\,
            I => \bfn_14_24_0_\
        );

    \I__313\ : InMux
    port map (
            O => \N__3009\,
            I => n2318
        );

    \I__312\ : InMux
    port map (
            O => \N__3006\,
            I => \N__3002\
        );

    \I__311\ : InMux
    port map (
            O => \N__3005\,
            I => \N__2999\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__3002\,
            I => blink_counter_25
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2999\,
            I => blink_counter_25
        );

    \I__308\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2991\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2991\,
            I => n16
        );

    \I__306\ : InMux
    port map (
            O => \N__2988\,
            I => n2303
        );

    \I__305\ : InMux
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2982\,
            I => n15
        );

    \I__303\ : InMux
    port map (
            O => \N__2979\,
            I => n2304
        );

    \I__302\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2973\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2973\,
            I => n14
        );

    \I__300\ : InMux
    port map (
            O => \N__2970\,
            I => n2305
        );

    \I__299\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2964\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2964\,
            I => n13
        );

    \I__297\ : InMux
    port map (
            O => \N__2961\,
            I => n2306
        );

    \I__296\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2955\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2955\,
            I => n12
        );

    \I__294\ : InMux
    port map (
            O => \N__2952\,
            I => n2307
        );

    \I__293\ : InMux
    port map (
            O => \N__2949\,
            I => \N__2946\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2946\,
            I => n11
        );

    \I__291\ : InMux
    port map (
            O => \N__2943\,
            I => n2308
        );

    \I__290\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2937\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2937\,
            I => n10
        );

    \I__288\ : InMux
    port map (
            O => \N__2934\,
            I => \bfn_14_23_0_\
        );

    \I__287\ : InMux
    port map (
            O => \N__2931\,
            I => \N__2928\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2928\,
            I => n9
        );

    \I__285\ : InMux
    port map (
            O => \N__2925\,
            I => n2310
        );

    \I__284\ : InMux
    port map (
            O => \N__2922\,
            I => \N__2919\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2919\,
            I => n8_adj_409
        );

    \I__282\ : InMux
    port map (
            O => \N__2916\,
            I => n2311
        );

    \I__281\ : InMux
    port map (
            O => \N__2913\,
            I => \N__2910\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2910\,
            I => n24
        );

    \I__279\ : InMux
    port map (
            O => \N__2907\,
            I => n2295
        );

    \I__278\ : InMux
    port map (
            O => \N__2904\,
            I => \N__2901\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2901\,
            I => n23
        );

    \I__276\ : InMux
    port map (
            O => \N__2898\,
            I => n2296
        );

    \I__275\ : InMux
    port map (
            O => \N__2895\,
            I => \N__2892\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2892\,
            I => n22
        );

    \I__273\ : InMux
    port map (
            O => \N__2889\,
            I => n2297
        );

    \I__272\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2883\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2883\,
            I => n21
        );

    \I__270\ : InMux
    port map (
            O => \N__2880\,
            I => n2298
        );

    \I__269\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2874\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2874\,
            I => n20
        );

    \I__267\ : InMux
    port map (
            O => \N__2871\,
            I => n2299
        );

    \I__266\ : InMux
    port map (
            O => \N__2868\,
            I => \N__2865\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2865\,
            I => n19
        );

    \I__264\ : InMux
    port map (
            O => \N__2862\,
            I => n2300
        );

    \I__263\ : InMux
    port map (
            O => \N__2859\,
            I => \N__2856\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2856\,
            I => n18
        );

    \I__261\ : InMux
    port map (
            O => \N__2853\,
            I => \bfn_14_22_0_\
        );

    \I__260\ : InMux
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2847\,
            I => n17
        );

    \I__258\ : InMux
    port map (
            O => \N__2844\,
            I => n2302
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__2841\,
            I => \n2553_cascade_\
        );

    \I__256\ : IoInMux
    port map (
            O => \N__2838\,
            I => \N__2835\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2835\,
            I => \N__2832\
        );

    \I__254\ : Span12Mux_s9_v
    port map (
            O => \N__2832\,
            I => \N__2829\
        );

    \I__253\ : Odrv12
    port map (
            O => \N__2829\,
            I => \LED_c\
        );

    \I__252\ : InMux
    port map (
            O => \N__2826\,
            I => \N__2823\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2823\,
            I => n2554
        );

    \I__250\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2817\,
            I => n26
        );

    \I__248\ : InMux
    port map (
            O => \N__2814\,
            I => \bfn_14_21_0_\
        );

    \I__247\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2808\,
            I => n25
        );

    \I__245\ : InMux
    port map (
            O => \N__2805\,
            I => n2294
        );

    \I__244\ : IoInMux
    port map (
            O => \N__2802\,
            I => \N__2799\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2799\,
            I => \N__2796\
        );

    \I__242\ : IoSpan4Mux
    port map (
            O => \N__2796\,
            I => \N__2793\
        );

    \I__241\ : IoSpan4Mux
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__240\ : IoSpan4Mux
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__239\ : Odrv4
    port map (
            O => \N__2787\,
            I => \CLK_pad_gb_input\
        );

    \INVeeprom.i2c.i2c_scl_enable_124C\ : INV
    port map (
            O => \INVeeprom.i2c.i2c_scl_enable_124C_net\,
            I => \N__6181\
        );

    \INVeeprom.i2c.sda_out_133C\ : INV
    port map (
            O => \INVeeprom.i2c.sda_out_133C_net\,
            I => \N__6153\
        );

    \INVeeprom.i2c.write_enable_132C\ : INV
    port map (
            O => \INVeeprom.i2c.write_enable_132C_net\,
            I => \N__6129\
        );

    \IN_MUX_bfv_21_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_22_0_\
        );

    \IN_MUX_bfv_21_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_18_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n2248\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2270,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2278,
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2286,
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2301,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2309,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2317,
            carryinitout => \bfn_14_24_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2802\,
            GLOBALBUFFEROUTPUT => \CLK_N\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i1635_4_lut_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000000"
        )
    port map (
            in0 => \N__3026\,
            in1 => \N__3068\,
            in2 => \N__3050\,
            in3 => \N__3086\,
            lcout => OPEN,
            ltout => \n2553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1637_3_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__2826\,
            in1 => \_gnd_net_\,
            in2 => \N__2841\,
            in3 => \N__3006\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1636_4_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010110000"
        )
    port map (
            in0 => \N__3027\,
            in1 => \N__3069\,
            in2 => \N__3051\,
            in3 => \N__3087\,
            lcout => n2554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i0_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2820\,
            in2 => \_gnd_net_\,
            in3 => \N__2814\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => n2294,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i1_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2811\,
            in2 => \_gnd_net_\,
            in3 => \N__2805\,
            lcout => n25,
            ltout => OPEN,
            carryin => n2294,
            carryout => n2295,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i2_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2913\,
            in2 => \_gnd_net_\,
            in3 => \N__2907\,
            lcout => n24,
            ltout => OPEN,
            carryin => n2295,
            carryout => n2296,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i3_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2904\,
            in2 => \_gnd_net_\,
            in3 => \N__2898\,
            lcout => n23,
            ltout => OPEN,
            carryin => n2296,
            carryout => n2297,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i4_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2895\,
            in2 => \_gnd_net_\,
            in3 => \N__2889\,
            lcout => n22,
            ltout => OPEN,
            carryin => n2297,
            carryout => n2298,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i5_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2886\,
            in2 => \_gnd_net_\,
            in3 => \N__2880\,
            lcout => n21,
            ltout => OPEN,
            carryin => n2298,
            carryout => n2299,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i6_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2877\,
            in2 => \_gnd_net_\,
            in3 => \N__2871\,
            lcout => n20,
            ltout => OPEN,
            carryin => n2299,
            carryout => n2300,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i7_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2868\,
            in2 => \_gnd_net_\,
            in3 => \N__2862\,
            lcout => n19,
            ltout => OPEN,
            carryin => n2300,
            carryout => n2301,
            clk => \N__5117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i8_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2859\,
            in2 => \_gnd_net_\,
            in3 => \N__2853\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => n2302,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i9_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2850\,
            in2 => \_gnd_net_\,
            in3 => \N__2844\,
            lcout => n17,
            ltout => OPEN,
            carryin => n2302,
            carryout => n2303,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i10_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2994\,
            in2 => \_gnd_net_\,
            in3 => \N__2988\,
            lcout => n16,
            ltout => OPEN,
            carryin => n2303,
            carryout => n2304,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i11_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2985\,
            in2 => \_gnd_net_\,
            in3 => \N__2979\,
            lcout => n15,
            ltout => OPEN,
            carryin => n2304,
            carryout => n2305,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i12_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2976\,
            in2 => \_gnd_net_\,
            in3 => \N__2970\,
            lcout => n14,
            ltout => OPEN,
            carryin => n2305,
            carryout => n2306,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i13_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2967\,
            in2 => \_gnd_net_\,
            in3 => \N__2961\,
            lcout => n13,
            ltout => OPEN,
            carryin => n2306,
            carryout => n2307,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i14_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2958\,
            in2 => \_gnd_net_\,
            in3 => \N__2952\,
            lcout => n12,
            ltout => OPEN,
            carryin => n2307,
            carryout => n2308,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i15_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2949\,
            in2 => \_gnd_net_\,
            in3 => \N__2943\,
            lcout => n11,
            ltout => OPEN,
            carryin => n2308,
            carryout => n2309,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i16_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2940\,
            in2 => \_gnd_net_\,
            in3 => \N__2934\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => n2310,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i17_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2931\,
            in2 => \_gnd_net_\,
            in3 => \N__2925\,
            lcout => n9,
            ltout => OPEN,
            carryin => n2310,
            carryout => n2311,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i18_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2922\,
            in2 => \_gnd_net_\,
            in3 => \N__2916\,
            lcout => n8_adj_409,
            ltout => OPEN,
            carryin => n2311,
            carryout => n2312,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i19_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3105\,
            in2 => \_gnd_net_\,
            in3 => \N__3099\,
            lcout => n7,
            ltout => OPEN,
            carryin => n2312,
            carryout => n2313,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i20_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3096\,
            in2 => \_gnd_net_\,
            in3 => \N__3090\,
            lcout => n6_adj_410,
            ltout => OPEN,
            carryin => n2313,
            carryout => n2314,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i21_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3085\,
            in2 => \_gnd_net_\,
            in3 => \N__3072\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n2314,
            carryout => n2315,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i22_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3067\,
            in2 => \_gnd_net_\,
            in3 => \N__3054\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n2315,
            carryout => n2316,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i23_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3043\,
            in2 => \_gnd_net_\,
            in3 => \N__3030\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n2316,
            carryout => n2317,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i24_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3025\,
            in2 => \_gnd_net_\,
            in3 => \N__3012\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => n2318,
            clk => \N__5126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_363__i25_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3005\,
            in2 => \_gnd_net_\,
            in3 => \N__3009\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.enable_39_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000100"
        )
    port map (
            in0 => \N__3604\,
            in1 => \N__4538\,
            in2 => \N__5952\,
            in3 => \N__4221\,
            lcout => \eeprom.enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5118\,
            ce => 'H',
            sr => \N__3960\
        );

    \eeprom.i1696_2_lut_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5951\,
            in2 => \_gnd_net_\,
            in3 => \N__3603\,
            lcout => \eeprom.n642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_4_lut_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3226\,
            in1 => \N__3277\,
            in2 => \N__3347\,
            in3 => \N__3310\,
            lcout => \eeprom.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i12_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__3278\,
            in1 => \N__4530\,
            in2 => \N__3264\,
            in3 => \N__4342\,
            lcout => \eeprom.delay_counter_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i8_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111010000"
        )
    port map (
            in0 => \N__4531\,
            in1 => \N__3297\,
            in2 => \N__4371\,
            in3 => \N__3311\,
            lcout => \eeprom.delay_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i6_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__3343\,
            in1 => \N__4529\,
            in2 => \N__4370\,
            in3 => \N__3327\,
            lcout => \eeprom.delay_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i2_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__3227\,
            in1 => \N__4349\,
            in2 => \N__3213\,
            in3 => \N__4528\,
            lcout => \eeprom.delay_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.mux_182_Mux_0_i1_4_lut_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__4473\,
            in1 => \N__4220\,
            in2 => \N__5946\,
            in3 => \N__3606\,
            lcout => OPEN,
            ltout => \n693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rw_43_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__4763\,
            in1 => \N__3952\,
            in2 => \N__3111\,
            in3 => \N__4474\,
            lcout => rw,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_13_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4219\,
            in1 => \N__3951\,
            in2 => \_gnd_net_\,
            in3 => \N__4472\,
            lcout => \eeprom.n1601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_counter_362__i0_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3726\,
            in2 => \_gnd_net_\,
            in3 => \N__3108\,
            lcout => delay_counter_0,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => n2263,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i1_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3884\,
            in2 => \_gnd_net_\,
            in3 => \N__3138\,
            lcout => delay_counter_1,
            ltout => OPEN,
            carryin => n2263,
            carryout => n2264,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i2_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4247\,
            in2 => \_gnd_net_\,
            in3 => \N__3135\,
            lcout => delay_counter_2,
            ltout => OPEN,
            carryin => n2264,
            carryout => n2265,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i3_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3740\,
            in2 => \_gnd_net_\,
            in3 => \N__3132\,
            lcout => delay_counter_3,
            ltout => OPEN,
            carryin => n2265,
            carryout => n2266,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i4_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3870\,
            in2 => \_gnd_net_\,
            in3 => \N__3129\,
            lcout => delay_counter_4,
            ltout => OPEN,
            carryin => n2266,
            carryout => n2267,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i5_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4271\,
            in2 => \_gnd_net_\,
            in3 => \N__3126\,
            lcout => delay_counter_5,
            ltout => OPEN,
            carryin => n2267,
            carryout => n2268,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i6_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3753\,
            in2 => \_gnd_net_\,
            in3 => \N__3123\,
            lcout => delay_counter_6,
            ltout => OPEN,
            carryin => n2268,
            carryout => n2269,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i7_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3909\,
            in2 => \_gnd_net_\,
            in3 => \N__3120\,
            lcout => delay_counter_7,
            ltout => OPEN,
            carryin => n2269,
            carryout => n2270,
            clk => \N__5127\,
            ce => 'H',
            sr => \N__4116\
        );

    \delay_counter_362__i8_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3897\,
            in2 => \_gnd_net_\,
            in3 => \N__3117\,
            lcout => delay_counter_8,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => n2271,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i9_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3765\,
            in2 => \_gnd_net_\,
            in3 => \N__3114\,
            lcout => delay_counter_9,
            ltout => OPEN,
            carryin => n2271,
            carryout => n2272,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i10_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3858\,
            in2 => \_gnd_net_\,
            in3 => \N__3165\,
            lcout => delay_counter_10,
            ltout => OPEN,
            carryin => n2272,
            carryout => n2273,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i11_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3833\,
            in2 => \_gnd_net_\,
            in3 => \N__3162\,
            lcout => delay_counter_11,
            ltout => OPEN,
            carryin => n2273,
            carryout => n2274,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i12_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3846\,
            in2 => \_gnd_net_\,
            in3 => \N__3159\,
            lcout => delay_counter_12,
            ltout => OPEN,
            carryin => n2274,
            carryout => n2275,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i13_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3819\,
            in2 => \_gnd_net_\,
            in3 => \N__3156\,
            lcout => delay_counter_13,
            ltout => OPEN,
            carryin => n2275,
            carryout => n2276,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i14_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3690\,
            in2 => \_gnd_net_\,
            in3 => \N__3153\,
            lcout => delay_counter_14,
            ltout => OPEN,
            carryin => n2276,
            carryout => n2277,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i15_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3702\,
            in2 => \_gnd_net_\,
            in3 => \N__3150\,
            lcout => delay_counter_15,
            ltout => OPEN,
            carryin => n2277,
            carryout => n2278,
            clk => \N__5130\,
            ce => 'H',
            sr => \N__4111\
        );

    \delay_counter_362__i16_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3804\,
            in2 => \_gnd_net_\,
            in3 => \N__3147\,
            lcout => delay_counter_16,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => n2279,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i17_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3714\,
            in2 => \_gnd_net_\,
            in3 => \N__3144\,
            lcout => delay_counter_17,
            ltout => OPEN,
            carryin => n2279,
            carryout => n2280,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i18_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3792\,
            in2 => \_gnd_net_\,
            in3 => \N__3141\,
            lcout => delay_counter_18,
            ltout => OPEN,
            carryin => n2280,
            carryout => n2281,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i19_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3777\,
            in2 => \_gnd_net_\,
            in3 => \N__3192\,
            lcout => delay_counter_19,
            ltout => OPEN,
            carryin => n2281,
            carryout => n2282,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i20_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4163\,
            in2 => \_gnd_net_\,
            in3 => \N__3189\,
            lcout => delay_counter_20,
            ltout => OPEN,
            carryin => n2282,
            carryout => n2283,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i21_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3672\,
            in2 => \_gnd_net_\,
            in3 => \N__3186\,
            lcout => delay_counter_21,
            ltout => OPEN,
            carryin => n2283,
            carryout => n2284,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i22_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4188\,
            in2 => \_gnd_net_\,
            in3 => \N__3183\,
            lcout => delay_counter_22,
            ltout => OPEN,
            carryin => n2284,
            carryout => n2285,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i23_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3660\,
            in2 => \_gnd_net_\,
            in3 => \N__3180\,
            lcout => delay_counter_23,
            ltout => OPEN,
            carryin => n2285,
            carryout => n2286,
            clk => \N__5134\,
            ce => 'H',
            sr => \N__4101\
        );

    \delay_counter_362__i24_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3999\,
            in2 => \_gnd_net_\,
            in3 => \N__3177\,
            lcout => delay_counter_24,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => n2287,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \delay_counter_362__i25_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4176\,
            in2 => \_gnd_net_\,
            in3 => \N__3174\,
            lcout => delay_counter_25,
            ltout => OPEN,
            carryin => n2287,
            carryout => n2288,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \delay_counter_362__i26_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4038\,
            in2 => \_gnd_net_\,
            in3 => \N__3171\,
            lcout => delay_counter_26,
            ltout => OPEN,
            carryin => n2288,
            carryout => n2289,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \delay_counter_362__i27_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4013\,
            in2 => \_gnd_net_\,
            in3 => \N__3168\,
            lcout => delay_counter_27,
            ltout => OPEN,
            carryin => n2289,
            carryout => n2290,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \delay_counter_362__i28_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4062\,
            in2 => \_gnd_net_\,
            in3 => \N__3249\,
            lcout => delay_counter_28,
            ltout => OPEN,
            carryin => n2290,
            carryout => n2291,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \delay_counter_362__i29_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4074\,
            in2 => \_gnd_net_\,
            in3 => \N__3246\,
            lcout => delay_counter_29,
            ltout => OPEN,
            carryin => n2291,
            carryout => n2292,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \delay_counter_362__i30_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4026\,
            in2 => \_gnd_net_\,
            in3 => \N__3243\,
            lcout => delay_counter_30,
            ltout => OPEN,
            carryin => n2292,
            carryout => n2293,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \delay_counter_362__i31_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4135\,
            in2 => \_gnd_net_\,
            in3 => \N__3240\,
            lcout => delay_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5135\,
            ce => 'H',
            sr => \N__4112\
        );

    \eeprom.add_158_2_lut_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3516\,
            in2 => \N__3426\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.delay_counter_15_N_171_0\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \eeprom.n2241\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_3_lut_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3453\,
            in2 => \N__3548\,
            in3 => \N__3237\,
            lcout => \eeprom.delay_counter_15_N_171_1\,
            ltout => OPEN,
            carryin => \eeprom.n2241\,
            carryout => \eeprom.n2242\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_4_lut_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3520\,
            in2 => \N__3234\,
            in3 => \N__3201\,
            lcout => \eeprom.delay_counter_15_N_171_2\,
            ltout => OPEN,
            carryin => \eeprom.n2242\,
            carryout => \eeprom.n2243\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_5_lut_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4699\,
            in2 => \N__3549\,
            in3 => \N__3198\,
            lcout => \eeprom.delay_counter_15_N_171_3\,
            ltout => OPEN,
            carryin => \eeprom.n2243\,
            carryout => \eeprom.n2244\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_6_lut_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3524\,
            in2 => \N__3633\,
            in3 => \N__3195\,
            lcout => \eeprom.delay_counter_15_N_171_4\,
            ltout => OPEN,
            carryin => \eeprom.n2244\,
            carryout => \eeprom.n2245\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_7_lut_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3396\,
            in2 => \N__3550\,
            in3 => \N__3354\,
            lcout => \eeprom.delay_counter_15_N_171_5\,
            ltout => OPEN,
            carryin => \eeprom.n2245\,
            carryout => \eeprom.n2246\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_8_lut_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3528\,
            in2 => \N__3351\,
            in3 => \N__3318\,
            lcout => \eeprom.delay_counter_15_N_171_6\,
            ltout => OPEN,
            carryin => \eeprom.n2246\,
            carryout => \eeprom.n2247\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_9_lut_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4649\,
            in2 => \N__3551\,
            in3 => \N__3315\,
            lcout => \eeprom.delay_counter_15_N_171_7\,
            ltout => OPEN,
            carryin => \eeprom.n2247\,
            carryout => \eeprom.n2248\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_10_lut_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3312\,
            in2 => \N__3552\,
            in3 => \N__3291\,
            lcout => \eeprom.delay_counter_15_N_171_8\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \eeprom.n2249\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_11_lut_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3535\,
            in2 => \N__4622\,
            in3 => \N__3288\,
            lcout => \eeprom.delay_counter_15_N_171_9\,
            ltout => OPEN,
            carryin => \eeprom.n2249\,
            carryout => \eeprom.n2250\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_12_lut_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3371\,
            in2 => \N__3553\,
            in3 => \N__3285\,
            lcout => \eeprom.delay_counter_15_N_171_10\,
            ltout => OPEN,
            carryin => \eeprom.n2250\,
            carryout => \eeprom.n2251\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_13_lut_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3539\,
            in2 => \N__4668\,
            in3 => \N__3282\,
            lcout => \eeprom.delay_counter_15_N_171_11\,
            ltout => OPEN,
            carryin => \eeprom.n2251\,
            carryout => \eeprom.n2252\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_14_lut_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3279\,
            in2 => \N__3554\,
            in3 => \N__3255\,
            lcout => \eeprom.delay_counter_15_N_171_12\,
            ltout => OPEN,
            carryin => \eeprom.n2252\,
            carryout => \eeprom.n2253\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_15_lut_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3543\,
            in2 => \N__4293\,
            in3 => \N__3252\,
            lcout => \eeprom.delay_counter_15_N_171_13\,
            ltout => OPEN,
            carryin => \eeprom.n2253\,
            carryout => \eeprom.n2254\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_16_lut_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4563\,
            in2 => \N__3555\,
            in3 => \N__3558\,
            lcout => \eeprom.delay_counter_15_N_171_14\,
            ltout => OPEN,
            carryin => \eeprom.n2254\,
            carryout => \eeprom.n2255\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_158_17_lut_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__4584\,
            in1 => \N__3547\,
            in2 => \_gnd_net_\,
            in3 => \N__3477\,
            lcout => \eeprom.delay_counter_15_N_171_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_15_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3418\,
            in1 => \N__3391\,
            in2 => \N__3372\,
            in3 => \N__3625\,
            lcout => OPEN,
            ltout => \eeprom.n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3474\,
            in2 => \N__3468\,
            in3 => \N__4288\,
            lcout => OPEN,
            ltout => \eeprom.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3448\,
            in1 => \N__4704\,
            in2 => \N__3465\,
            in3 => \N__4596\,
            lcout => \eeprom.n1500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i1_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__3462\,
            in1 => \N__4356\,
            in2 => \N__4544\,
            in3 => \N__3449\,
            lcout => \eeprom.delay_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i0_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__3419\,
            in1 => \N__4517\,
            in2 => \N__4372\,
            in3 => \N__3435\,
            lcout => \eeprom.delay_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i5_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__3392\,
            in1 => \N__4358\,
            in2 => \N__4546\,
            in3 => \N__3405\,
            lcout => \eeprom.delay_counter_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i10_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__3370\,
            in1 => \N__4518\,
            in2 => \N__4373\,
            in3 => \N__3378\,
            lcout => \eeprom.delay_counter_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i4_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000101110"
        )
    port map (
            in0 => \N__3626\,
            in1 => \N__4357\,
            in2 => \N__4545\,
            in3 => \N__3642\,
            lcout => \eeprom.delay_counter_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1682_2_lut_3_lut_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__4469\,
            in1 => \N__5929\,
            in2 => \_gnd_net_\,
            in3 => \N__3947\,
            lcout => \eeprom.n2453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.data_ready_42_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000010"
        )
    port map (
            in0 => \N__3949\,
            in1 => \N__4471\,
            in2 => \N__5944\,
            in3 => \N__3612\,
            lcout => n324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_10_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5661\,
            lcout => n41,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i525_3_lut_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101000"
        )
    port map (
            in0 => \N__3948\,
            in1 => \N__4468\,
            in2 => \N__5945\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n1018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2_2_lut_adj_14_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3605\,
            in2 => \_gnd_net_\,
            in3 => \N__5550\,
            lcout => OPEN,
            ltout => \n6_adj_405_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1566_4_lut_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__5777\,
            in1 => \N__4467\,
            in2 => \N__3585\,
            in3 => \N__3582\,
            lcout => OPEN,
            ltout => \n2483_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2_4_lut_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__4218\,
            in1 => \N__3576\,
            in2 => \N__3570\,
            in3 => \N__3567\,
            lcout => n1568,
            ltout => \n1568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i1_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__3950\,
            in1 => \N__4470\,
            in2 => \N__3561\,
            in3 => \_gnd_net_\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i0_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__5947\,
            in1 => \N__3953\,
            in2 => \_gnd_net_\,
            in3 => \N__4516\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5131\,
            ce => \N__3918\,
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3908\,
            in1 => \N__3896\,
            in2 => \N__3885\,
            in3 => \N__3869\,
            lcout => n17_adj_406,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__3857\,
            in1 => \N__3845\,
            in2 => \N__3834\,
            in3 => \N__4227\,
            lcout => OPEN,
            ltout => \n2512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__3818\,
            in1 => \N__3678\,
            in2 => \N__3807\,
            in3 => \N__3803\,
            lcout => OPEN,
            ltout => \n2495_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__3791\,
            in1 => \N__3648\,
            in2 => \N__3780\,
            in3 => \N__3776\,
            lcout => n8_adj_412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3764\,
            in1 => \N__3752\,
            in2 => \N__3741\,
            in3 => \N__3725\,
            lcout => n16_adj_407,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_3_lut_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3713\,
            in1 => \N__3701\,
            in2 => \_gnd_net_\,
            in3 => \N__3689\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3671\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3659\,
            lcout => n6_adj_413,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4272\,
            in1 => \N__4257\,
            in2 => \N__4251\,
            in3 => \N__4233\,
            lcout => n2536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \read_15_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__4137\,
            in1 => \N__4050\,
            in2 => \N__3987\,
            in3 => \N__4143\,
            lcout => \read_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5136\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_19_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__4187\,
            in1 => \N__4175\,
            in2 => \N__4164\,
            in3 => \N__4149\,
            lcout => n9_adj_404,
            ltout => \n9_adj_404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1011_4_lut_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__4136\,
            in1 => \N__4049\,
            in2 => \N__4119\,
            in3 => \N__3983\,
            lcout => \addr_10__N_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4073\,
            in2 => \_gnd_net_\,
            in3 => \N__4061\,
            lcout => n10_adj_403,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_18_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4037\,
            in1 => \N__4025\,
            in2 => \N__4014\,
            in3 => \N__3998\,
            lcout => n14_adj_401,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i7_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__4548\,
            in1 => \N__4408\,
            in2 => \N__4650\,
            in3 => \N__3966\,
            lcout => \eeprom.delay_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i3_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__4547\,
            in1 => \N__4700\,
            in2 => \N__4413\,
            in3 => \N__4710\,
            lcout => \eeprom.delay_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i11_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__4540\,
            in1 => \N__4664\,
            in2 => \N__4410\,
            in3 => \N__4680\,
            lcout => \eeprom.delay_counter_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i9_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__4404\,
            in1 => \N__4543\,
            in2 => \N__4623\,
            in3 => \N__4674\,
            lcout => \eeprom.delay_counter_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2_2_lut_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4561\,
            in2 => \_gnd_net_\,
            in3 => \N__4582\,
            lcout => OPEN,
            ltout => \eeprom.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2_4_lut_adj_16_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4663\,
            in1 => \N__4642\,
            in2 => \N__4626\,
            in3 => \N__4609\,
            lcout => \eeprom.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i15_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__4542\,
            in1 => \N__4583\,
            in2 => \N__4412\,
            in3 => \N__4590\,
            lcout => \eeprom.delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i14_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__4541\,
            in1 => \N__4569\,
            in2 => \N__4411\,
            in3 => \N__4562\,
            lcout => \eeprom.delay_counter_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_clk_122_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5066\,
            lcout => \eeprom.i2c.i2c_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i13_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__4539\,
            in1 => \N__4292\,
            in2 => \N__4409\,
            in3 => \N__4299\,
            lcout => \eeprom.delay_counter_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.write_enable_132_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4799\,
            in1 => \N__5761\,
            in2 => \_gnd_net_\,
            in3 => \N__5861\,
            lcout => sda_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.write_enable_132C_net\,
            ce => \N__4719\,
            sr => \N__4740\
        );

    \eeprom.i2c.i22_3_lut_3_lut_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__5517\,
            in1 => \N__5616\,
            in2 => \_gnd_net_\,
            in3 => \N__5726\,
            lcout => \eeprom.i2c.n11_adj_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i56_3_lut_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__5724\,
            in1 => \N__5516\,
            in2 => \_gnd_net_\,
            in3 => \N__5837\,
            lcout => \eeprom.i2c.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__5840\,
            in1 => \N__5618\,
            in2 => \N__5539\,
            in3 => \N__5727\,
            lcout => n11_adj_399,
            ltout => \n11_adj_399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1673_2_lut_3_lut_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4924\,
            in2 => \N__4743\,
            in3 => \N__4958\,
            lcout => n2569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_adj_9_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4986\,
            in1 => \N__5617\,
            in2 => \_gnd_net_\,
            in3 => \N__4731\,
            lcout => \eeprom.i2c.n1669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_4_lut_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110010"
        )
    port map (
            in0 => \N__5725\,
            in1 => \N__5515\,
            in2 => \N__5648\,
            in3 => \N__5838\,
            lcout => \eeprom.i2c.n37\,
            ltout => \eeprom.i2c.n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_adj_8_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5615\,
            in2 => \N__4734\,
            in3 => \N__4730\,
            lcout => \eeprom.i2c.n39\,
            ltout => \eeprom.i2c.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1692_4_lut_4_lut_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__5619\,
            in1 => \N__4798\,
            in2 => \N__4722\,
            in3 => \N__5839\,
            lcout => \eeprom.i2c.n1027\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.sda_out_133_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__5874\,
            in1 => \N__4866\,
            in2 => \N__4803\,
            in3 => \N__5768\,
            lcout => sda_out,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.sda_out_133C_net\,
            ce => \N__4998\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5147\,
            in2 => \_gnd_net_\,
            in3 => \N__5195\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4_4_lut_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5210\,
            in1 => \N__5180\,
            in2 => \N__4782\,
            in3 => \N__5165\,
            lcout => \eeprom.i2c.counter2_7__N_256\,
            ltout => \eeprom.i2c.counter2_7__N_256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6117\,
            in2 => \N__4779\,
            in3 => \N__4849\,
            lcout => \eeprom.i2c.n1580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.enable_slow_121_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5065\,
            lcout => \state_7_N_269_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5132\,
            ce => \N__4776\,
            sr => \N__4856\
        );

    \eeprom.i2c.state_i0_i0_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111111"
        )
    port map (
            in0 => \N__5776\,
            in1 => \N__5250\,
            in2 => \N__5457\,
            in3 => \N__4884\,
            lcout => state_0_adj_397,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.saved_addr__i1_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__5909\,
            in1 => \N__5264\,
            in2 => \N__4770\,
            in3 => \N__5040\,
            lcout => saved_addr_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1004_2_lut_3_lut_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__5637\,
            in1 => \N__5772\,
            in2 => \_gnd_net_\,
            in3 => \N__5857\,
            lcout => n1835,
            ltout => \n1835_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__5354\,
            in1 => \_gnd_net_\,
            in2 => \N__4752\,
            in3 => \N__5537\,
            lcout => n949,
            ltout => \n949_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i2_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100000111"
        )
    port map (
            in0 => \N__5456\,
            in1 => \N__4749\,
            in2 => \N__4887\,
            in3 => \N__5859\,
            lcout => state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1630_4_lut_4_lut_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001011"
        )
    port map (
            in0 => \N__5858\,
            in1 => \N__5638\,
            in2 => \N__5778\,
            in3 => \N__5538\,
            lcout => OPEN,
            ltout => \n2547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i1_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001011"
        )
    port map (
            in0 => \N__5639\,
            in1 => \N__4883\,
            in2 => \N__4872\,
            in3 => \N__5010\,
            lcout => state_1_adj_396,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1667_2_lut_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5038\,
            in2 => \_gnd_net_\,
            in3 => \N__6379\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n2574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1666_4_lut_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000000000"
        )
    port map (
            in0 => \N__6347\,
            in1 => \N__5335\,
            in2 => \N__4869\,
            in3 => \N__5623\,
            lcout => \eeprom.i2c.n2557\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2_4_lut_4_lut_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101011101"
        )
    port map (
            in0 => \N__5624\,
            in1 => \N__5758\,
            in2 => \N__4860\,
            in3 => \N__6245\,
            lcout => OPEN,
            ltout => \n2538_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__6246\,
            in1 => \N__5021\,
            in2 => \N__4824\,
            in3 => \N__5392\,
            lcout => OPEN,
            ltout => \n4_adj_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__5625\,
            in1 => \N__4809\,
            in2 => \N__4821\,
            in3 => \N__5759\,
            lcout => OPEN,
            ltout => \n2507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i3_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111000"
        )
    port map (
            in0 => \N__5536\,
            in1 => \N__4818\,
            in2 => \N__4812\,
            in3 => \N__5355\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_142_i10_2_lut_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5535\,
            in2 => \_gnd_net_\,
            in3 => \N__5860\,
            lcout => n10_adj_394,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1674_3_lut_4_lut_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__5039\,
            in1 => \N__4923\,
            in2 => \N__5025\,
            in3 => \N__4959\,
            lcout => n2566,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1686_4_lut_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001100"
        )
    port map (
            in0 => \N__5651\,
            in1 => \N__5004\,
            in2 => \N__4968\,
            in3 => \N__5870\,
            lcout => \eeprom.i2c.n2406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5872\,
            in1 => \N__5767\,
            in2 => \_gnd_net_\,
            in3 => \N__5523\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n1051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i17_4_lut_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011111000"
        )
    port map (
            in0 => \N__4985\,
            in1 => \N__5403\,
            in2 => \N__4971\,
            in3 => \N__4896\,
            lcout => \eeprom.i2c.n1548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_2_lut_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5765\,
            in2 => \_gnd_net_\,
            in3 => \N__5521\,
            lcout => \eeprom.i2c.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i463_2_lut_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4957\,
            in2 => \_gnd_net_\,
            in3 => \N__4928\,
            lcout => \state_7_N_285_3\,
            ltout => \state_7_N_285_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1558_3_lut_4_lut_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__5871\,
            in1 => \N__5217\,
            in2 => \N__4899\,
            in3 => \N__5522\,
            lcout => \eeprom.i2c.n2475\,
            ltout => \eeprom.i2c.n2475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1545_2_lut_4_lut_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__5769\,
            in2 => \N__4890\,
            in3 => \N__5873\,
            lcout => \eeprom.i2c.n1655\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_142_i9_2_lut_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5766\,
            in2 => \_gnd_net_\,
            in3 => \N__5652\,
            lcout => \eeprom.i2c.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter2_364_365__i1_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5211\,
            in2 => \_gnd_net_\,
            in3 => \N__5199\,
            lcout => \eeprom.i2c.counter2_0\,
            ltout => OPEN,
            carryin => \bfn_21_18_0_\,
            carryout => \eeprom.i2c.n2319\,
            clk => \N__5133\,
            ce => 'H',
            sr => \N__5070\
        );

    \eeprom.i2c.counter2_364_365__i2_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5196\,
            in2 => \_gnd_net_\,
            in3 => \N__5184\,
            lcout => \eeprom.i2c.counter2_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2319\,
            carryout => \eeprom.i2c.n2320\,
            clk => \N__5133\,
            ce => 'H',
            sr => \N__5070\
        );

    \eeprom.i2c.counter2_364_365__i3_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5181\,
            in2 => \_gnd_net_\,
            in3 => \N__5169\,
            lcout => \eeprom.i2c.counter2_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2320\,
            carryout => \eeprom.i2c.n2321\,
            clk => \N__5133\,
            ce => 'H',
            sr => \N__5070\
        );

    \eeprom.i2c.counter2_364_365__i4_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5166\,
            in2 => \_gnd_net_\,
            in3 => \N__5154\,
            lcout => \eeprom.i2c.counter2_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2321\,
            carryout => \eeprom.i2c.n2322\,
            clk => \N__5133\,
            ce => 'H',
            sr => \N__5070\
        );

    \eeprom.i2c.counter2_364_365__i5_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5148\,
            in2 => \_gnd_net_\,
            in3 => \N__5151\,
            lcout => \eeprom.i2c.counter2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5133\,
            ce => 'H',
            sr => \N__5070\
        );

    \eeprom.i2c.data_out_i0_i7_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__5430\,
            in1 => \N__6424\,
            in2 => \N__5049\,
            in3 => \N__6269\,
            lcout => n306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_25_i11_2_lut_3_lut_4_lut_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5741\,
            in1 => \N__5525\,
            in2 => \N__5649\,
            in3 => \N__5841\,
            lcout => n15_adj_393,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__5843\,
            in1 => \N__5742\,
            in2 => \N__5650\,
            in3 => \N__5533\,
            lcout => n11_adj_400,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_4_lut_adj_12_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__5745\,
            in1 => \N__5343\,
            in2 => \N__5397\,
            in3 => \N__5631\,
            lcout => n1518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5842\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5532\,
            lcout => n10_adj_398,
            ltout => \n10_adj_398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_4_lut_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__5744\,
            in1 => \N__5342\,
            in2 => \N__5268\,
            in3 => \N__5630\,
            lcout => n1523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_3_lut_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__5844\,
            in1 => \N__5265\,
            in2 => \_gnd_net_\,
            in3 => \N__5534\,
            lcout => OPEN,
            ltout => \n2460_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1676_4_lut_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__5743\,
            in1 => \N__5372\,
            in2 => \N__5253\,
            in3 => \N__5629\,
            lcout => n2560,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i6_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__6258\,
            in1 => \N__5241\,
            in2 => \N__6312\,
            in3 => \N__5429\,
            lcout => n308,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i0_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__5414\,
            in1 => \N__6306\,
            in2 => \N__5235\,
            in3 => \N__6256\,
            lcout => n320,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i1_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__6257\,
            in1 => \N__6433\,
            in2 => \N__5226\,
            in3 => \N__5415\,
            lcout => n318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_50_i4_2_lut_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6346\,
            in2 => \_gnd_net_\,
            in3 => \N__6380\,
            lcout => n4_adj_408,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i986_2_lut_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6348\,
            lcout => n1817,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i5_4_lut_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5334\,
            in1 => \N__6050\,
            in2 => \N__5288\,
            in3 => \N__5303\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i6_4_lut_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6014\,
            in1 => \N__6032\,
            in2 => \N__5418\,
            in3 => \N__5413\,
            lcout => \eeprom.i2c.n942\,
            ltout => \eeprom.i2c.n942_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__5396\,
            in1 => \N__5373\,
            in2 => \N__5358\,
            in3 => \N__5760\,
            lcout => n1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter_i0_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5336\,
            in2 => \_gnd_net_\,
            in3 => \N__5313\,
            lcout => \eeprom.i2c.counter_0\,
            ltout => OPEN,
            carryin => \bfn_21_22_0_\,
            carryout => \eeprom.i2c.n2256\,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \eeprom.i2c.counter_i1_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6382\,
            in2 => \N__5986\,
            in3 => \N__5310\,
            lcout => \eeprom.i2c.counter_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2256\,
            carryout => \eeprom.i2c.n2257\,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \eeprom.i2c.counter_i2_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5976\,
            in2 => \N__6354\,
            in3 => \N__5307\,
            lcout => \eeprom.i2c.counter_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2257\,
            carryout => \eeprom.i2c.n2258\,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \eeprom.i2c.counter_i3_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5304\,
            in2 => \N__5987\,
            in3 => \N__5292\,
            lcout => \eeprom.i2c.counter_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2258\,
            carryout => \eeprom.i2c.n2259\,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \eeprom.i2c.counter_i4_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5980\,
            in2 => \N__5289\,
            in3 => \N__5271\,
            lcout => \eeprom.i2c.counter_4\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2259\,
            carryout => \eeprom.i2c.n2260\,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \eeprom.i2c.counter_i5_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6051\,
            in2 => \N__5988\,
            in3 => \N__6039\,
            lcout => \eeprom.i2c.counter_5\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2260\,
            carryout => \eeprom.i2c.n2261\,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \eeprom.i2c.counter_i6_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5984\,
            in2 => \N__6036\,
            in3 => \N__6021\,
            lcout => \eeprom.i2c.counter_6\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2261\,
            carryout => \eeprom.i2c.n2262\,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \eeprom.i2c.counter_i7_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__5985\,
            in1 => \N__6015\,
            in2 => \_gnd_net_\,
            in3 => \N__6018\,
            lcout => \eeprom.i2c.counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6169\,
            ce => \N__6003\,
            sr => \N__5997\
        );

    \CONSTANT_ONE_LUT4_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i26_2_lut_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5770\,
            in2 => \_gnd_net_\,
            in3 => \N__5548\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_scl_enable_124_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__5908\,
            in1 => \N__5653\,
            in2 => \N__5880\,
            in3 => \N__5875\,
            lcout => scl_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.i2c_scl_enable_124C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i995_3_lut_4_lut_4_lut_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111011111"
        )
    port map (
            in0 => \N__5876\,
            in1 => \N__5771\,
            in2 => \N__5660\,
            in3 => \N__5549\,
            lcout => n1826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i3_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__6266\,
            in1 => \N__6318\,
            in2 => \N__5439\,
            in3 => \N__6434\,
            lcout => n314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_45_i4_2_lut_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6383\,
            in2 => \_gnd_net_\,
            in3 => \N__6352\,
            lcout => n4_adj_395,
            ltout => \n4_adj_395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i5_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__6435\,
            in1 => \N__6405\,
            in2 => \N__6408\,
            in3 => \N__6268\,
            lcout => n310,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i4_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__6399\,
            in1 => \N__6311\,
            in2 => \N__6393\,
            in3 => \N__6267\,
            lcout => n312,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_48_i4_2_lut_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6384\,
            in2 => \_gnd_net_\,
            in3 => \N__6353\,
            lcout => n4,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i2_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__6213\,
            in1 => \N__6310\,
            in2 => \N__6285\,
            in3 => \N__6265\,
            lcout => n316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i989_2_lut_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__6194\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6182\,
            lcout => scl_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
