-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Feb 4 2020 19:52:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : in std_logic;
    SCL : in std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__56636\ : std_logic;
signal \N__56635\ : std_logic;
signal \N__56634\ : std_logic;
signal \N__56627\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56625\ : std_logic;
signal \N__56618\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56616\ : std_logic;
signal \N__56609\ : std_logic;
signal \N__56608\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56600\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56591\ : std_logic;
signal \N__56590\ : std_logic;
signal \N__56589\ : std_logic;
signal \N__56582\ : std_logic;
signal \N__56581\ : std_logic;
signal \N__56580\ : std_logic;
signal \N__56573\ : std_logic;
signal \N__56572\ : std_logic;
signal \N__56571\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56563\ : std_logic;
signal \N__56562\ : std_logic;
signal \N__56555\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56553\ : std_logic;
signal \N__56546\ : std_logic;
signal \N__56545\ : std_logic;
signal \N__56544\ : std_logic;
signal \N__56537\ : std_logic;
signal \N__56536\ : std_logic;
signal \N__56535\ : std_logic;
signal \N__56528\ : std_logic;
signal \N__56527\ : std_logic;
signal \N__56526\ : std_logic;
signal \N__56519\ : std_logic;
signal \N__56518\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56510\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56508\ : std_logic;
signal \N__56501\ : std_logic;
signal \N__56500\ : std_logic;
signal \N__56499\ : std_logic;
signal \N__56492\ : std_logic;
signal \N__56491\ : std_logic;
signal \N__56490\ : std_logic;
signal \N__56483\ : std_logic;
signal \N__56482\ : std_logic;
signal \N__56481\ : std_logic;
signal \N__56474\ : std_logic;
signal \N__56473\ : std_logic;
signal \N__56472\ : std_logic;
signal \N__56455\ : std_logic;
signal \N__56452\ : std_logic;
signal \N__56449\ : std_logic;
signal \N__56446\ : std_logic;
signal \N__56443\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56437\ : std_logic;
signal \N__56436\ : std_logic;
signal \N__56435\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56431\ : std_logic;
signal \N__56430\ : std_logic;
signal \N__56429\ : std_logic;
signal \N__56424\ : std_logic;
signal \N__56421\ : std_logic;
signal \N__56418\ : std_logic;
signal \N__56413\ : std_logic;
signal \N__56410\ : std_logic;
signal \N__56407\ : std_logic;
signal \N__56404\ : std_logic;
signal \N__56399\ : std_logic;
signal \N__56392\ : std_logic;
signal \N__56391\ : std_logic;
signal \N__56390\ : std_logic;
signal \N__56389\ : std_logic;
signal \N__56388\ : std_logic;
signal \N__56383\ : std_logic;
signal \N__56382\ : std_logic;
signal \N__56377\ : std_logic;
signal \N__56376\ : std_logic;
signal \N__56375\ : std_logic;
signal \N__56374\ : std_logic;
signal \N__56371\ : std_logic;
signal \N__56368\ : std_logic;
signal \N__56365\ : std_logic;
signal \N__56362\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56350\ : std_logic;
signal \N__56347\ : std_logic;
signal \N__56344\ : std_logic;
signal \N__56341\ : std_logic;
signal \N__56336\ : std_logic;
signal \N__56333\ : std_logic;
signal \N__56330\ : std_logic;
signal \N__56323\ : std_logic;
signal \N__56320\ : std_logic;
signal \N__56317\ : std_logic;
signal \N__56314\ : std_logic;
signal \N__56309\ : std_logic;
signal \N__56302\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56300\ : std_logic;
signal \N__56297\ : std_logic;
signal \N__56296\ : std_logic;
signal \N__56295\ : std_logic;
signal \N__56294\ : std_logic;
signal \N__56291\ : std_logic;
signal \N__56286\ : std_logic;
signal \N__56283\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56277\ : std_logic;
signal \N__56276\ : std_logic;
signal \N__56275\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56257\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56255\ : std_logic;
signal \N__56254\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56252\ : std_logic;
signal \N__56251\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56241\ : std_logic;
signal \N__56238\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56221\ : std_logic;
signal \N__56216\ : std_logic;
signal \N__56211\ : std_logic;
signal \N__56206\ : std_logic;
signal \N__56197\ : std_logic;
signal \N__56196\ : std_logic;
signal \N__56195\ : std_logic;
signal \N__56194\ : std_logic;
signal \N__56191\ : std_logic;
signal \N__56188\ : std_logic;
signal \N__56187\ : std_logic;
signal \N__56184\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56180\ : std_logic;
signal \N__56175\ : std_logic;
signal \N__56174\ : std_logic;
signal \N__56169\ : std_logic;
signal \N__56166\ : std_logic;
signal \N__56165\ : std_logic;
signal \N__56162\ : std_logic;
signal \N__56159\ : std_logic;
signal \N__56156\ : std_logic;
signal \N__56151\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56145\ : std_logic;
signal \N__56142\ : std_logic;
signal \N__56139\ : std_logic;
signal \N__56134\ : std_logic;
signal \N__56133\ : std_logic;
signal \N__56130\ : std_logic;
signal \N__56127\ : std_logic;
signal \N__56124\ : std_logic;
signal \N__56121\ : std_logic;
signal \N__56118\ : std_logic;
signal \N__56115\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56107\ : std_logic;
signal \N__56098\ : std_logic;
signal \N__56097\ : std_logic;
signal \N__56096\ : std_logic;
signal \N__56095\ : std_logic;
signal \N__56094\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56092\ : std_logic;
signal \N__56091\ : std_logic;
signal \N__56090\ : std_logic;
signal \N__56089\ : std_logic;
signal \N__56088\ : std_logic;
signal \N__56087\ : std_logic;
signal \N__56086\ : std_logic;
signal \N__56085\ : std_logic;
signal \N__56084\ : std_logic;
signal \N__56083\ : std_logic;
signal \N__56082\ : std_logic;
signal \N__56081\ : std_logic;
signal \N__56080\ : std_logic;
signal \N__56079\ : std_logic;
signal \N__56078\ : std_logic;
signal \N__56077\ : std_logic;
signal \N__56076\ : std_logic;
signal \N__56075\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56073\ : std_logic;
signal \N__56072\ : std_logic;
signal \N__56071\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56069\ : std_logic;
signal \N__56068\ : std_logic;
signal \N__56067\ : std_logic;
signal \N__56066\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56064\ : std_logic;
signal \N__56063\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56061\ : std_logic;
signal \N__56060\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56058\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56055\ : std_logic;
signal \N__56054\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56052\ : std_logic;
signal \N__56051\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56049\ : std_logic;
signal \N__56048\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56046\ : std_logic;
signal \N__56045\ : std_logic;
signal \N__56044\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56042\ : std_logic;
signal \N__56041\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56039\ : std_logic;
signal \N__55918\ : std_logic;
signal \N__55915\ : std_logic;
signal \N__55912\ : std_logic;
signal \N__55909\ : std_logic;
signal \N__55908\ : std_logic;
signal \N__55905\ : std_logic;
signal \N__55902\ : std_logic;
signal \N__55901\ : std_logic;
signal \N__55900\ : std_logic;
signal \N__55897\ : std_logic;
signal \N__55894\ : std_logic;
signal \N__55891\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55887\ : std_logic;
signal \N__55884\ : std_logic;
signal \N__55879\ : std_logic;
signal \N__55876\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55864\ : std_logic;
signal \N__55861\ : std_logic;
signal \N__55860\ : std_logic;
signal \N__55859\ : std_logic;
signal \N__55856\ : std_logic;
signal \N__55855\ : std_logic;
signal \N__55852\ : std_logic;
signal \N__55849\ : std_logic;
signal \N__55846\ : std_logic;
signal \N__55843\ : std_logic;
signal \N__55840\ : std_logic;
signal \N__55837\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55829\ : std_logic;
signal \N__55826\ : std_logic;
signal \N__55823\ : std_logic;
signal \N__55816\ : std_logic;
signal \N__55813\ : std_logic;
signal \N__55810\ : std_logic;
signal \N__55807\ : std_logic;
signal \N__55804\ : std_logic;
signal \N__55801\ : std_logic;
signal \N__55798\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55792\ : std_logic;
signal \N__55789\ : std_logic;
signal \N__55786\ : std_logic;
signal \N__55783\ : std_logic;
signal \N__55780\ : std_logic;
signal \N__55777\ : std_logic;
signal \N__55774\ : std_logic;
signal \N__55771\ : std_logic;
signal \N__55768\ : std_logic;
signal \N__55767\ : std_logic;
signal \N__55766\ : std_logic;
signal \N__55763\ : std_logic;
signal \N__55758\ : std_logic;
signal \N__55755\ : std_logic;
signal \N__55752\ : std_logic;
signal \N__55747\ : std_logic;
signal \N__55744\ : std_logic;
signal \N__55741\ : std_logic;
signal \N__55738\ : std_logic;
signal \N__55735\ : std_logic;
signal \N__55732\ : std_logic;
signal \N__55729\ : std_logic;
signal \N__55726\ : std_logic;
signal \N__55723\ : std_logic;
signal \N__55720\ : std_logic;
signal \N__55717\ : std_logic;
signal \N__55714\ : std_logic;
signal \N__55713\ : std_logic;
signal \N__55712\ : std_logic;
signal \N__55711\ : std_logic;
signal \N__55710\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55708\ : std_logic;
signal \N__55707\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55703\ : std_logic;
signal \N__55702\ : std_logic;
signal \N__55701\ : std_logic;
signal \N__55700\ : std_logic;
signal \N__55699\ : std_logic;
signal \N__55698\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55696\ : std_logic;
signal \N__55695\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55682\ : std_logic;
signal \N__55679\ : std_logic;
signal \N__55676\ : std_logic;
signal \N__55673\ : std_logic;
signal \N__55668\ : std_logic;
signal \N__55657\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55655\ : std_logic;
signal \N__55654\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55652\ : std_logic;
signal \N__55651\ : std_logic;
signal \N__55648\ : std_logic;
signal \N__55645\ : std_logic;
signal \N__55644\ : std_logic;
signal \N__55641\ : std_logic;
signal \N__55638\ : std_logic;
signal \N__55633\ : std_logic;
signal \N__55628\ : std_logic;
signal \N__55623\ : std_logic;
signal \N__55618\ : std_logic;
signal \N__55615\ : std_logic;
signal \N__55608\ : std_logic;
signal \N__55605\ : std_logic;
signal \N__55602\ : std_logic;
signal \N__55599\ : std_logic;
signal \N__55596\ : std_logic;
signal \N__55587\ : std_logic;
signal \N__55576\ : std_logic;
signal \N__55567\ : std_logic;
signal \N__55564\ : std_logic;
signal \N__55563\ : std_logic;
signal \N__55560\ : std_logic;
signal \N__55557\ : std_logic;
signal \N__55552\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55546\ : std_logic;
signal \N__55543\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55537\ : std_logic;
signal \N__55534\ : std_logic;
signal \N__55531\ : std_logic;
signal \N__55528\ : std_logic;
signal \N__55525\ : std_logic;
signal \N__55522\ : std_logic;
signal \N__55519\ : std_logic;
signal \N__55516\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55508\ : std_logic;
signal \N__55507\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55501\ : std_logic;
signal \N__55496\ : std_logic;
signal \N__55495\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55486\ : std_logic;
signal \N__55483\ : std_logic;
signal \N__55476\ : std_logic;
signal \N__55471\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55469\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55463\ : std_logic;
signal \N__55460\ : std_logic;
signal \N__55457\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55426\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55417\ : std_logic;
signal \N__55414\ : std_logic;
signal \N__55411\ : std_logic;
signal \N__55408\ : std_logic;
signal \N__55405\ : std_logic;
signal \N__55402\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55393\ : std_logic;
signal \N__55392\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55386\ : std_logic;
signal \N__55383\ : std_logic;
signal \N__55382\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55374\ : std_logic;
signal \N__55369\ : std_logic;
signal \N__55366\ : std_logic;
signal \N__55363\ : std_logic;
signal \N__55362\ : std_logic;
signal \N__55359\ : std_logic;
signal \N__55356\ : std_logic;
signal \N__55353\ : std_logic;
signal \N__55352\ : std_logic;
signal \N__55349\ : std_logic;
signal \N__55346\ : std_logic;
signal \N__55343\ : std_logic;
signal \N__55336\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55330\ : std_logic;
signal \N__55329\ : std_logic;
signal \N__55326\ : std_logic;
signal \N__55325\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55316\ : std_logic;
signal \N__55309\ : std_logic;
signal \N__55306\ : std_logic;
signal \N__55305\ : std_logic;
signal \N__55302\ : std_logic;
signal \N__55299\ : std_logic;
signal \N__55296\ : std_logic;
signal \N__55295\ : std_logic;
signal \N__55292\ : std_logic;
signal \N__55289\ : std_logic;
signal \N__55286\ : std_logic;
signal \N__55279\ : std_logic;
signal \N__55276\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55269\ : std_logic;
signal \N__55268\ : std_logic;
signal \N__55265\ : std_logic;
signal \N__55262\ : std_logic;
signal \N__55259\ : std_logic;
signal \N__55252\ : std_logic;
signal \N__55249\ : std_logic;
signal \N__55248\ : std_logic;
signal \N__55247\ : std_logic;
signal \N__55246\ : std_logic;
signal \N__55243\ : std_logic;
signal \N__55240\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55236\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55233\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55229\ : std_logic;
signal \N__55228\ : std_logic;
signal \N__55227\ : std_logic;
signal \N__55226\ : std_logic;
signal \N__55225\ : std_logic;
signal \N__55224\ : std_logic;
signal \N__55223\ : std_logic;
signal \N__55222\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55219\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55216\ : std_logic;
signal \N__55215\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55213\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55211\ : std_logic;
signal \N__55210\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55202\ : std_logic;
signal \N__55193\ : std_logic;
signal \N__55192\ : std_logic;
signal \N__55191\ : std_logic;
signal \N__55190\ : std_logic;
signal \N__55189\ : std_logic;
signal \N__55188\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55185\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55175\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55173\ : std_logic;
signal \N__55172\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55168\ : std_logic;
signal \N__55167\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55161\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55153\ : std_logic;
signal \N__55146\ : std_logic;
signal \N__55145\ : std_logic;
signal \N__55142\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55140\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55136\ : std_logic;
signal \N__55135\ : std_logic;
signal \N__55134\ : std_logic;
signal \N__55133\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55131\ : std_logic;
signal \N__55130\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55128\ : std_logic;
signal \N__55127\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55122\ : std_logic;
signal \N__55121\ : std_logic;
signal \N__55118\ : std_logic;
signal \N__55117\ : std_logic;
signal \N__55114\ : std_logic;
signal \N__55113\ : std_logic;
signal \N__55110\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55106\ : std_logic;
signal \N__55103\ : std_logic;
signal \N__55102\ : std_logic;
signal \N__55099\ : std_logic;
signal \N__55098\ : std_logic;
signal \N__55095\ : std_logic;
signal \N__55094\ : std_logic;
signal \N__55091\ : std_logic;
signal \N__55090\ : std_logic;
signal \N__55089\ : std_logic;
signal \N__55088\ : std_logic;
signal \N__55087\ : std_logic;
signal \N__55086\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55084\ : std_logic;
signal \N__55083\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55081\ : std_logic;
signal \N__55080\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55078\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55073\ : std_logic;
signal \N__55072\ : std_logic;
signal \N__55071\ : std_logic;
signal \N__55070\ : std_logic;
signal \N__55069\ : std_logic;
signal \N__55068\ : std_logic;
signal \N__55067\ : std_logic;
signal \N__55066\ : std_logic;
signal \N__55065\ : std_logic;
signal \N__55064\ : std_logic;
signal \N__55063\ : std_logic;
signal \N__55062\ : std_logic;
signal \N__55061\ : std_logic;
signal \N__55060\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55054\ : std_logic;
signal \N__55047\ : std_logic;
signal \N__55044\ : std_logic;
signal \N__55041\ : std_logic;
signal \N__55038\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55034\ : std_logic;
signal \N__55031\ : std_logic;
signal \N__55026\ : std_logic;
signal \N__55019\ : std_logic;
signal \N__55010\ : std_logic;
signal \N__55001\ : std_logic;
signal \N__54998\ : std_logic;
signal \N__54997\ : std_logic;
signal \N__54996\ : std_logic;
signal \N__54995\ : std_logic;
signal \N__54994\ : std_logic;
signal \N__54993\ : std_logic;
signal \N__54992\ : std_logic;
signal \N__54991\ : std_logic;
signal \N__54990\ : std_logic;
signal \N__54989\ : std_logic;
signal \N__54988\ : std_logic;
signal \N__54987\ : std_logic;
signal \N__54986\ : std_logic;
signal \N__54985\ : std_logic;
signal \N__54984\ : std_logic;
signal \N__54983\ : std_logic;
signal \N__54982\ : std_logic;
signal \N__54981\ : std_logic;
signal \N__54980\ : std_logic;
signal \N__54979\ : std_logic;
signal \N__54978\ : std_logic;
signal \N__54977\ : std_logic;
signal \N__54976\ : std_logic;
signal \N__54975\ : std_logic;
signal \N__54968\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54952\ : std_logic;
signal \N__54951\ : std_logic;
signal \N__54950\ : std_logic;
signal \N__54949\ : std_logic;
signal \N__54948\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54946\ : std_logic;
signal \N__54945\ : std_logic;
signal \N__54942\ : std_logic;
signal \N__54941\ : std_logic;
signal \N__54940\ : std_logic;
signal \N__54939\ : std_logic;
signal \N__54938\ : std_logic;
signal \N__54937\ : std_logic;
signal \N__54936\ : std_logic;
signal \N__54935\ : std_logic;
signal \N__54934\ : std_logic;
signal \N__54931\ : std_logic;
signal \N__54928\ : std_logic;
signal \N__54927\ : std_logic;
signal \N__54926\ : std_logic;
signal \N__54925\ : std_logic;
signal \N__54924\ : std_logic;
signal \N__54923\ : std_logic;
signal \N__54922\ : std_logic;
signal \N__54921\ : std_logic;
signal \N__54920\ : std_logic;
signal \N__54917\ : std_logic;
signal \N__54914\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54905\ : std_logic;
signal \N__54902\ : std_logic;
signal \N__54899\ : std_logic;
signal \N__54896\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54890\ : std_logic;
signal \N__54889\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54887\ : std_logic;
signal \N__54886\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54883\ : std_logic;
signal \N__54882\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54880\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54878\ : std_logic;
signal \N__54877\ : std_logic;
signal \N__54876\ : std_logic;
signal \N__54875\ : std_logic;
signal \N__54874\ : std_logic;
signal \N__54873\ : std_logic;
signal \N__54872\ : std_logic;
signal \N__54871\ : std_logic;
signal \N__54870\ : std_logic;
signal \N__54869\ : std_logic;
signal \N__54868\ : std_logic;
signal \N__54867\ : std_logic;
signal \N__54866\ : std_logic;
signal \N__54865\ : std_logic;
signal \N__54848\ : std_logic;
signal \N__54831\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54827\ : std_logic;
signal \N__54824\ : std_logic;
signal \N__54823\ : std_logic;
signal \N__54820\ : std_logic;
signal \N__54819\ : std_logic;
signal \N__54816\ : std_logic;
signal \N__54815\ : std_logic;
signal \N__54812\ : std_logic;
signal \N__54809\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54803\ : std_logic;
signal \N__54800\ : std_logic;
signal \N__54797\ : std_logic;
signal \N__54794\ : std_logic;
signal \N__54791\ : std_logic;
signal \N__54788\ : std_logic;
signal \N__54785\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54779\ : std_logic;
signal \N__54774\ : std_logic;
signal \N__54773\ : std_logic;
signal \N__54772\ : std_logic;
signal \N__54771\ : std_logic;
signal \N__54770\ : std_logic;
signal \N__54769\ : std_logic;
signal \N__54768\ : std_logic;
signal \N__54767\ : std_logic;
signal \N__54762\ : std_logic;
signal \N__54759\ : std_logic;
signal \N__54756\ : std_logic;
signal \N__54749\ : std_logic;
signal \N__54748\ : std_logic;
signal \N__54745\ : std_logic;
signal \N__54744\ : std_logic;
signal \N__54743\ : std_logic;
signal \N__54742\ : std_logic;
signal \N__54741\ : std_logic;
signal \N__54740\ : std_logic;
signal \N__54739\ : std_logic;
signal \N__54738\ : std_logic;
signal \N__54735\ : std_logic;
signal \N__54734\ : std_logic;
signal \N__54733\ : std_logic;
signal \N__54732\ : std_logic;
signal \N__54731\ : std_logic;
signal \N__54730\ : std_logic;
signal \N__54729\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54727\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54717\ : std_logic;
signal \N__54712\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54701\ : std_logic;
signal \N__54700\ : std_logic;
signal \N__54699\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54689\ : std_logic;
signal \N__54686\ : std_logic;
signal \N__54683\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54679\ : std_logic;
signal \N__54678\ : std_logic;
signal \N__54677\ : std_logic;
signal \N__54676\ : std_logic;
signal \N__54673\ : std_logic;
signal \N__54670\ : std_logic;
signal \N__54669\ : std_logic;
signal \N__54668\ : std_logic;
signal \N__54665\ : std_logic;
signal \N__54662\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54650\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54646\ : std_logic;
signal \N__54643\ : std_logic;
signal \N__54640\ : std_logic;
signal \N__54637\ : std_logic;
signal \N__54634\ : std_logic;
signal \N__54631\ : std_logic;
signal \N__54628\ : std_logic;
signal \N__54625\ : std_logic;
signal \N__54622\ : std_logic;
signal \N__54621\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54619\ : std_logic;
signal \N__54618\ : std_logic;
signal \N__54617\ : std_logic;
signal \N__54616\ : std_logic;
signal \N__54615\ : std_logic;
signal \N__54614\ : std_logic;
signal \N__54613\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54611\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54606\ : std_logic;
signal \N__54605\ : std_logic;
signal \N__54604\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54598\ : std_logic;
signal \N__54597\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54595\ : std_logic;
signal \N__54594\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54590\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54584\ : std_logic;
signal \N__54583\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54570\ : std_logic;
signal \N__54567\ : std_logic;
signal \N__54560\ : std_logic;
signal \N__54549\ : std_logic;
signal \N__54546\ : std_logic;
signal \N__54539\ : std_logic;
signal \N__54536\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54532\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54521\ : std_logic;
signal \N__54520\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54518\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54514\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54510\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54506\ : std_logic;
signal \N__54505\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54498\ : std_logic;
signal \N__54495\ : std_logic;
signal \N__54488\ : std_logic;
signal \N__54479\ : std_logic;
signal \N__54472\ : std_logic;
signal \N__54471\ : std_logic;
signal \N__54468\ : std_logic;
signal \N__54465\ : std_logic;
signal \N__54462\ : std_logic;
signal \N__54459\ : std_logic;
signal \N__54456\ : std_logic;
signal \N__54453\ : std_logic;
signal \N__54450\ : std_logic;
signal \N__54447\ : std_logic;
signal \N__54444\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54438\ : std_logic;
signal \N__54435\ : std_logic;
signal \N__54432\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54428\ : std_logic;
signal \N__54425\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54413\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54407\ : std_logic;
signal \N__54404\ : std_logic;
signal \N__54403\ : std_logic;
signal \N__54400\ : std_logic;
signal \N__54397\ : std_logic;
signal \N__54394\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54358\ : std_logic;
signal \N__54347\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54345\ : std_logic;
signal \N__54344\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54342\ : std_logic;
signal \N__54341\ : std_logic;
signal \N__54340\ : std_logic;
signal \N__54339\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54322\ : std_logic;
signal \N__54321\ : std_logic;
signal \N__54318\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54299\ : std_logic;
signal \N__54292\ : std_logic;
signal \N__54287\ : std_logic;
signal \N__54284\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54272\ : std_logic;
signal \N__54267\ : std_logic;
signal \N__54266\ : std_logic;
signal \N__54263\ : std_logic;
signal \N__54260\ : std_logic;
signal \N__54257\ : std_logic;
signal \N__54256\ : std_logic;
signal \N__54255\ : std_logic;
signal \N__54254\ : std_logic;
signal \N__54253\ : std_logic;
signal \N__54252\ : std_logic;
signal \N__54251\ : std_logic;
signal \N__54250\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54248\ : std_logic;
signal \N__54245\ : std_logic;
signal \N__54242\ : std_logic;
signal \N__54241\ : std_logic;
signal \N__54240\ : std_logic;
signal \N__54235\ : std_logic;
signal \N__54230\ : std_logic;
signal \N__54227\ : std_logic;
signal \N__54220\ : std_logic;
signal \N__54213\ : std_logic;
signal \N__54204\ : std_logic;
signal \N__54201\ : std_logic;
signal \N__54198\ : std_logic;
signal \N__54191\ : std_logic;
signal \N__54186\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54163\ : std_logic;
signal \N__54154\ : std_logic;
signal \N__54143\ : std_logic;
signal \N__54134\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54124\ : std_logic;
signal \N__54119\ : std_logic;
signal \N__54116\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54112\ : std_logic;
signal \N__54109\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54103\ : std_logic;
signal \N__54100\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54090\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54084\ : std_logic;
signal \N__54083\ : std_logic;
signal \N__54082\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54078\ : std_logic;
signal \N__54077\ : std_logic;
signal \N__54070\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54059\ : std_logic;
signal \N__54058\ : std_logic;
signal \N__54057\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54018\ : std_logic;
signal \N__54013\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53993\ : std_logic;
signal \N__53992\ : std_logic;
signal \N__53991\ : std_logic;
signal \N__53990\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53974\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53938\ : std_logic;
signal \N__53929\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53909\ : std_logic;
signal \N__53906\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53892\ : std_logic;
signal \N__53891\ : std_logic;
signal \N__53890\ : std_logic;
signal \N__53887\ : std_logic;
signal \N__53884\ : std_logic;
signal \N__53881\ : std_logic;
signal \N__53878\ : std_logic;
signal \N__53877\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53870\ : std_logic;
signal \N__53869\ : std_logic;
signal \N__53866\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53861\ : std_logic;
signal \N__53860\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53858\ : std_logic;
signal \N__53855\ : std_logic;
signal \N__53852\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53841\ : std_logic;
signal \N__53840\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53837\ : std_logic;
signal \N__53836\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53834\ : std_logic;
signal \N__53833\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53831\ : std_logic;
signal \N__53830\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53828\ : std_logic;
signal \N__53827\ : std_logic;
signal \N__53822\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53796\ : std_logic;
signal \N__53793\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53790\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53783\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53774\ : std_logic;
signal \N__53773\ : std_logic;
signal \N__53770\ : std_logic;
signal \N__53769\ : std_logic;
signal \N__53768\ : std_logic;
signal \N__53767\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53764\ : std_logic;
signal \N__53755\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53736\ : std_logic;
signal \N__53719\ : std_logic;
signal \N__53714\ : std_logic;
signal \N__53711\ : std_logic;
signal \N__53702\ : std_logic;
signal \N__53697\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53687\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53677\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53673\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53668\ : std_logic;
signal \N__53667\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53665\ : std_logic;
signal \N__53664\ : std_logic;
signal \N__53663\ : std_logic;
signal \N__53662\ : std_logic;
signal \N__53659\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53625\ : std_logic;
signal \N__53622\ : std_logic;
signal \N__53621\ : std_logic;
signal \N__53620\ : std_logic;
signal \N__53617\ : std_logic;
signal \N__53616\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53611\ : std_logic;
signal \N__53608\ : std_logic;
signal \N__53593\ : std_logic;
signal \N__53584\ : std_logic;
signal \N__53581\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53569\ : std_logic;
signal \N__53566\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53564\ : std_logic;
signal \N__53563\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53561\ : std_logic;
signal \N__53560\ : std_logic;
signal \N__53557\ : std_logic;
signal \N__53554\ : std_logic;
signal \N__53551\ : std_logic;
signal \N__53550\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53536\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53524\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53514\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53507\ : std_logic;
signal \N__53504\ : std_logic;
signal \N__53501\ : std_logic;
signal \N__53500\ : std_logic;
signal \N__53497\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53489\ : std_logic;
signal \N__53486\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53484\ : std_logic;
signal \N__53483\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53479\ : std_logic;
signal \N__53472\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53451\ : std_logic;
signal \N__53444\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53426\ : std_logic;
signal \N__53419\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53416\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53400\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53388\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53373\ : std_logic;
signal \N__53370\ : std_logic;
signal \N__53367\ : std_logic;
signal \N__53366\ : std_logic;
signal \N__53363\ : std_logic;
signal \N__53362\ : std_logic;
signal \N__53361\ : std_logic;
signal \N__53360\ : std_logic;
signal \N__53359\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53353\ : std_logic;
signal \N__53352\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53348\ : std_logic;
signal \N__53347\ : std_logic;
signal \N__53344\ : std_logic;
signal \N__53341\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53337\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53307\ : std_logic;
signal \N__53296\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53284\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53274\ : std_logic;
signal \N__53265\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53252\ : std_logic;
signal \N__53243\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53225\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53215\ : std_logic;
signal \N__53210\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53179\ : std_logic;
signal \N__53178\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53172\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53151\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53137\ : std_logic;
signal \N__53126\ : std_logic;
signal \N__53125\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53108\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53098\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53083\ : std_logic;
signal \N__53066\ : std_logic;
signal \N__53065\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53054\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53044\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53017\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52991\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52985\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52968\ : std_logic;
signal \N__52961\ : std_logic;
signal \N__52950\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52921\ : std_logic;
signal \N__52918\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52914\ : std_logic;
signal \N__52913\ : std_logic;
signal \N__52910\ : std_logic;
signal \N__52907\ : std_logic;
signal \N__52904\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52896\ : std_logic;
signal \N__52893\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52887\ : std_logic;
signal \N__52884\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52882\ : std_logic;
signal \N__52881\ : std_logic;
signal \N__52876\ : std_logic;
signal \N__52873\ : std_logic;
signal \N__52870\ : std_logic;
signal \N__52869\ : std_logic;
signal \N__52866\ : std_logic;
signal \N__52865\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52840\ : std_logic;
signal \N__52835\ : std_logic;
signal \N__52828\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52823\ : std_logic;
signal \N__52820\ : std_logic;
signal \N__52817\ : std_logic;
signal \N__52814\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52806\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52798\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52792\ : std_logic;
signal \N__52789\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52776\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52767\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52760\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52748\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52732\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52725\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52714\ : std_logic;
signal \N__52711\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52705\ : std_logic;
signal \N__52702\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52695\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52688\ : std_logic;
signal \N__52685\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52674\ : std_logic;
signal \N__52671\ : std_logic;
signal \N__52670\ : std_logic;
signal \N__52667\ : std_logic;
signal \N__52664\ : std_logic;
signal \N__52661\ : std_logic;
signal \N__52654\ : std_logic;
signal \N__52651\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52644\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52637\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52624\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52617\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52607\ : std_logic;
signal \N__52604\ : std_logic;
signal \N__52601\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52568\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52555\ : std_logic;
signal \N__52554\ : std_logic;
signal \N__52551\ : std_logic;
signal \N__52550\ : std_logic;
signal \N__52547\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52534\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52530\ : std_logic;
signal \N__52527\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52517\ : std_logic;
signal \N__52510\ : std_logic;
signal \N__52507\ : std_logic;
signal \N__52504\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52470\ : std_logic;
signal \N__52467\ : std_logic;
signal \N__52466\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52424\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52403\ : std_logic;
signal \N__52400\ : std_logic;
signal \N__52397\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52373\ : std_logic;
signal \N__52370\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52360\ : std_logic;
signal \N__52357\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52353\ : std_logic;
signal \N__52352\ : std_logic;
signal \N__52349\ : std_logic;
signal \N__52346\ : std_logic;
signal \N__52343\ : std_logic;
signal \N__52336\ : std_logic;
signal \N__52333\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52329\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52325\ : std_logic;
signal \N__52322\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52309\ : std_logic;
signal \N__52306\ : std_logic;
signal \N__52305\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52298\ : std_logic;
signal \N__52295\ : std_logic;
signal \N__52292\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52280\ : std_logic;
signal \N__52277\ : std_logic;
signal \N__52274\ : std_logic;
signal \N__52271\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52262\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52252\ : std_logic;
signal \N__52249\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52238\ : std_logic;
signal \N__52235\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52196\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52180\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52164\ : std_logic;
signal \N__52161\ : std_logic;
signal \N__52158\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52134\ : std_logic;
signal \N__52133\ : std_logic;
signal \N__52130\ : std_logic;
signal \N__52127\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52114\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52074\ : std_logic;
signal \N__52071\ : std_logic;
signal \N__52068\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52060\ : std_logic;
signal \N__52057\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52040\ : std_logic;
signal \N__52037\ : std_logic;
signal \N__52032\ : std_logic;
signal \N__52029\ : std_logic;
signal \N__52026\ : std_logic;
signal \N__52023\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51989\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51970\ : std_logic;
signal \N__51967\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51961\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51952\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51930\ : std_logic;
signal \N__51927\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51897\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51876\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51872\ : std_logic;
signal \N__51869\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51849\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51839\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51780\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51757\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51749\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51735\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51667\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51632\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51618\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51588\ : std_logic;
signal \N__51585\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51576\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51565\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51559\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51549\ : std_logic;
signal \N__51548\ : std_logic;
signal \N__51545\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51536\ : std_logic;
signal \N__51533\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51523\ : std_logic;
signal \N__51520\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51511\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51488\ : std_logic;
signal \N__51485\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51444\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51367\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51348\ : std_logic;
signal \N__51345\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51333\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51325\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51294\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51274\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51263\ : std_logic;
signal \N__51260\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51199\ : std_logic;
signal \N__51196\ : std_logic;
signal \N__51193\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51180\ : std_logic;
signal \N__51177\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51173\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51156\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51147\ : std_logic;
signal \N__51144\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51121\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51107\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51099\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51091\ : std_logic;
signal \N__51088\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51073\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51068\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51053\ : std_logic;
signal \N__51050\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51037\ : std_logic;
signal \N__51034\ : std_logic;
signal \N__51031\ : std_logic;
signal \N__51028\ : std_logic;
signal \N__51025\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51019\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51008\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__50998\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50992\ : std_logic;
signal \N__50989\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50947\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50935\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50929\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50918\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50890\ : std_logic;
signal \N__50887\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50865\ : std_logic;
signal \N__50862\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50846\ : std_logic;
signal \N__50839\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50827\ : std_logic;
signal \N__50824\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50779\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50764\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50745\ : std_logic;
signal \N__50742\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50683\ : std_logic;
signal \N__50680\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50668\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50638\ : std_logic;
signal \N__50635\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50620\ : std_logic;
signal \N__50617\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50524\ : std_logic;
signal \N__50521\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50503\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50190\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50096\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50090\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50072\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50065\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50029\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50024\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49963\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49777\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49584\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49330\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49245\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49162\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49054\ : std_logic;
signal \N__49051\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48938\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48906\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48880\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48371\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47626\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47574\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44467\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44077\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44027\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44005\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43279\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42273\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42091\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41902\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41602\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41549\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41539\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40975\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40936\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40927\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40840\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40768\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40366\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39874\ : std_logic;
signal \N__39871\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39781\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39703\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39154\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38569\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38543\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37447\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37411\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37102\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36313\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36261\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34924\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_17_0_\ : std_logic;
signal n12257 : std_logic;
signal n12258 : std_logic;
signal n12259 : std_logic;
signal n12260 : std_logic;
signal n12261 : std_logic;
signal n12262 : std_logic;
signal n12263 : std_logic;
signal n12264 : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal n12265 : std_logic;
signal n12266 : std_logic;
signal n12267 : std_logic;
signal n12268 : std_logic;
signal n12269 : std_logic;
signal n12270 : std_logic;
signal n12271 : std_logic;
signal n12272 : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal n12273 : std_logic;
signal n12274 : std_logic;
signal n12275 : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal n12239 : std_logic;
signal n12240 : std_logic;
signal n12241 : std_logic;
signal n12242 : std_logic;
signal n12243 : std_logic;
signal n12244 : std_logic;
signal n12245 : std_logic;
signal n12246 : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal n12247 : std_logic;
signal n12248 : std_logic;
signal n12249 : std_logic;
signal n12250 : std_logic;
signal n12251 : std_logic;
signal n12252 : std_logic;
signal n12253 : std_logic;
signal n12254 : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal n12255 : std_logic;
signal n12256 : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal n12206 : std_logic;
signal n12207 : std_logic;
signal n12208 : std_logic;
signal n12209 : std_logic;
signal n12210 : std_logic;
signal n12211 : std_logic;
signal n12212 : std_logic;
signal n12213 : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal n12214 : std_logic;
signal n12215 : std_logic;
signal n12216 : std_logic;
signal n12217 : std_logic;
signal n12218 : std_logic;
signal n12219 : std_logic;
signal n12220 : std_logic;
signal n12221 : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal \bfn_1_26_0_\ : std_logic;
signal n12177 : std_logic;
signal n12178 : std_logic;
signal n12179 : std_logic;
signal n12180 : std_logic;
signal n12181 : std_logic;
signal n12182 : std_logic;
signal n12183 : std_logic;
signal n12184 : std_logic;
signal \bfn_1_27_0_\ : std_logic;
signal n12185 : std_logic;
signal n12186 : std_logic;
signal n12187 : std_logic;
signal n12188 : std_logic;
signal n12189 : std_logic;
signal n12190 : std_logic;
signal \n1427_cascade_\ : std_logic;
signal \n1430_cascade_\ : std_logic;
signal n11638 : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal \debounce.n12654\ : std_logic;
signal \debounce.n12655\ : std_logic;
signal \debounce.n12656\ : std_logic;
signal \debounce.n12657\ : std_logic;
signal \debounce.n12658\ : std_logic;
signal \debounce.n12659\ : std_logic;
signal \debounce.n12660\ : std_logic;
signal \debounce.n12661\ : std_logic;
signal \bfn_1_30_0_\ : std_logic;
signal \debounce.n12662\ : std_logic;
signal \bfn_1_31_0_\ : std_logic;
signal n12122 : std_logic;
signal n12123 : std_logic;
signal n12124 : std_logic;
signal n12125 : std_logic;
signal n12126 : std_logic;
signal n12127 : std_logic;
signal n12128 : std_logic;
signal n12129 : std_logic;
signal \bfn_1_32_0_\ : std_logic;
signal n12130 : std_logic;
signal \debounce.cnt_reg_3\ : std_logic;
signal \debounce.cnt_reg_9\ : std_logic;
signal \debounce.cnt_reg_5\ : std_logic;
signal \debounce.cnt_reg_8\ : std_logic;
signal \debounce.cnt_reg_1\ : std_logic;
signal \debounce.cnt_reg_2\ : std_logic;
signal \debounce.n14472_cascade_\ : std_logic;
signal n2095 : std_logic;
signal n2094 : std_logic;
signal n2101 : std_logic;
signal n2200 : std_logic;
signal \n2133_cascade_\ : std_logic;
signal \n2232_cascade_\ : std_logic;
signal \n2331_cascade_\ : std_logic;
signal n2089 : std_logic;
signal n2188 : std_logic;
signal \n2121_cascade_\ : std_logic;
signal \n2220_cascade_\ : std_logic;
signal \n2319_cascade_\ : std_logic;
signal n2097 : std_logic;
signal \n2049_cascade_\ : std_logic;
signal n2183 : std_logic;
signal n2184 : std_logic;
signal n2084 : std_logic;
signal n2116 : std_logic;
signal n2115 : std_logic;
signal \n2116_cascade_\ : std_logic;
signal \n2148_cascade_\ : std_logic;
signal n2195 : std_logic;
signal n2087 : std_logic;
signal n2093 : std_logic;
signal n2085 : std_logic;
signal n2117 : std_logic;
signal \bfn_2_21_0_\ : std_logic;
signal n12222 : std_logic;
signal n12223 : std_logic;
signal n12224 : std_logic;
signal n12225 : std_logic;
signal n12226 : std_logic;
signal n12227 : std_logic;
signal n12228 : std_logic;
signal n12229 : std_logic;
signal \bfn_2_22_0_\ : std_logic;
signal n12230 : std_logic;
signal n12231 : std_logic;
signal n12232 : std_logic;
signal n12233 : std_logic;
signal n12234 : std_logic;
signal n12235 : std_logic;
signal n12236 : std_logic;
signal n12237 : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal n12238 : std_logic;
signal n2016 : std_logic;
signal n1888 : std_logic;
signal n1985 : std_logic;
signal n2017 : std_logic;
signal n1700 : std_logic;
signal n1699 : std_logic;
signal \n1731_cascade_\ : std_logic;
signal n1697 : std_logic;
signal \n1729_cascade_\ : std_logic;
signal n1701 : std_logic;
signal \n1733_cascade_\ : std_logic;
signal n1886 : std_logic;
signal n1698 : std_logic;
signal n1696 : std_logic;
signal \n1728_cascade_\ : std_logic;
signal n1695 : std_logic;
signal n1694 : std_logic;
signal n1689 : std_logic;
signal n1630 : std_logic;
signal \n13986_cascade_\ : std_logic;
signal \n1554_cascade_\ : std_logic;
signal n1629 : std_logic;
signal n1631 : std_logic;
signal \bfn_2_27_0_\ : std_logic;
signal n12152 : std_logic;
signal n12153 : std_logic;
signal n12154 : std_logic;
signal n12155 : std_logic;
signal n12156 : std_logic;
signal n12157 : std_logic;
signal n12158 : std_logic;
signal n12159 : std_logic;
signal \bfn_2_28_0_\ : std_logic;
signal n12160 : std_logic;
signal n12161 : std_logic;
signal n12162 : std_logic;
signal n12163 : std_logic;
signal n1491 : std_logic;
signal n26_adj_678 : std_logic;
signal \bfn_2_29_0_\ : std_logic;
signal n25_adj_677 : std_logic;
signal n12717 : std_logic;
signal n24_adj_676 : std_logic;
signal n12718 : std_logic;
signal n23_adj_675 : std_logic;
signal n12719 : std_logic;
signal n22_adj_674 : std_logic;
signal n12720 : std_logic;
signal n21_adj_673 : std_logic;
signal n12721 : std_logic;
signal n20_adj_672 : std_logic;
signal n12722 : std_logic;
signal n19_adj_671 : std_logic;
signal n12723 : std_logic;
signal n12724 : std_logic;
signal n18_adj_670 : std_logic;
signal \bfn_2_30_0_\ : std_logic;
signal n17_adj_669 : std_logic;
signal n12725 : std_logic;
signal n16_adj_668 : std_logic;
signal n12726 : std_logic;
signal n15_adj_667 : std_logic;
signal n12727 : std_logic;
signal n14_adj_666 : std_logic;
signal n12728 : std_logic;
signal n13_adj_665 : std_logic;
signal n12729 : std_logic;
signal n12_adj_664 : std_logic;
signal n12730 : std_logic;
signal n11_adj_663 : std_logic;
signal n12731 : std_logic;
signal n12732 : std_logic;
signal n10_adj_662 : std_logic;
signal \bfn_2_31_0_\ : std_logic;
signal n9_adj_661 : std_logic;
signal n12733 : std_logic;
signal n8_adj_660 : std_logic;
signal n12734 : std_logic;
signal n7_adj_659 : std_logic;
signal n12735 : std_logic;
signal n6_adj_658 : std_logic;
signal n12736 : std_logic;
signal n12737 : std_logic;
signal n12738 : std_logic;
signal n12739 : std_logic;
signal n12740 : std_logic;
signal \bfn_2_32_0_\ : std_logic;
signal n12741 : std_logic;
signal \debounce.cnt_reg_4\ : std_logic;
signal \debounce.cnt_reg_6\ : std_logic;
signal \debounce.cnt_reg_0\ : std_logic;
signal \debounce.cnt_reg_7\ : std_logic;
signal \debounce.n13\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal n12296 : std_logic;
signal n12297 : std_logic;
signal n2398 : std_logic;
signal n12298 : std_logic;
signal n12299 : std_logic;
signal n12300 : std_logic;
signal n12301 : std_logic;
signal n12302 : std_logic;
signal n12303 : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal n12304 : std_logic;
signal n12305 : std_logic;
signal n12306 : std_logic;
signal n12307 : std_logic;
signal n12308 : std_logic;
signal n12309 : std_logic;
signal n2386 : std_logic;
signal n12310 : std_logic;
signal n12311 : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal n12312 : std_logic;
signal n12313 : std_logic;
signal n12314 : std_logic;
signal n12315 : std_logic;
signal n12316 : std_logic;
signal n2098 : std_logic;
signal n2392 : std_logic;
signal n2096 : std_logic;
signal n2197 : std_logic;
signal n1996 : std_logic;
signal n2196 : std_logic;
signal n2201 : std_logic;
signal n14160 : std_logic;
signal n2186 : std_logic;
signal n2028 : std_logic;
signal n1989 : std_logic;
signal n1998 : std_logic;
signal n1994 : std_logic;
signal n2026 : std_logic;
signal n1887 : std_logic;
signal n1986 : std_logic;
signal \n1919_cascade_\ : std_logic;
signal n2018 : std_logic;
signal n1988 : std_logic;
signal n2020 : std_logic;
signal n1987 : std_logic;
signal n1991 : std_logic;
signal n1892 : std_logic;
signal n1924 : std_logic;
signal \n1924_cascade_\ : std_logic;
signal n1893 : std_logic;
signal n1891 : std_logic;
signal \n1923_cascade_\ : std_logic;
signal n1896 : std_logic;
signal n1899 : std_logic;
signal \n1822_cascade_\ : std_logic;
signal n1894 : std_logic;
signal n1688 : std_logic;
signal \n1720_cascade_\ : std_logic;
signal n1820 : std_logic;
signal \n1752_cascade_\ : std_logic;
signal n1821 : std_logic;
signal n13343 : std_logic;
signal \n14110_cascade_\ : std_logic;
signal \n1653_cascade_\ : std_logic;
signal n1691 : std_logic;
signal n13962 : std_logic;
signal n11694 : std_logic;
signal \n13968_cascade_\ : std_logic;
signal n14116 : std_logic;
signal n13972 : std_logic;
signal n1690 : std_logic;
signal n1628 : std_logic;
signal n14104 : std_logic;
signal n1624 : std_logic;
signal n1692 : std_logic;
signal n1626 : std_logic;
signal n1693 : std_logic;
signal n1632 : std_logic;
signal \n1632_cascade_\ : std_logic;
signal n1633 : std_logic;
signal n11634 : std_logic;
signal n1625 : std_logic;
signal n1623 : std_logic;
signal n1499 : std_logic;
signal \n1531_cascade_\ : std_logic;
signal n11698 : std_logic;
signal n1627 : std_logic;
signal n1430 : std_logic;
signal n1497 : std_logic;
signal n1498 : std_logic;
signal n1622 : std_logic;
signal n300 : std_logic;
signal n1501 : std_logic;
signal \n300_cascade_\ : std_logic;
signal n1490 : std_logic;
signal \n1522_cascade_\ : std_logic;
signal n1621 : std_logic;
signal n1495 : std_logic;
signal n1496 : std_logic;
signal \n1528_cascade_\ : std_logic;
signal \n13978_cascade_\ : std_logic;
signal n13984 : std_logic;
signal n1432 : std_logic;
signal n14088 : std_logic;
signal n1433 : std_logic;
signal \n1433_cascade_\ : std_logic;
signal n1500 : std_logic;
signal n1401 : std_logic;
signal \bfn_3_29_0_\ : std_logic;
signal n1400 : std_logic;
signal n12141 : std_logic;
signal n12142 : std_logic;
signal n1398 : std_logic;
signal n12143 : std_logic;
signal n12144 : std_logic;
signal n12145 : std_logic;
signal n1395 : std_logic;
signal n12146 : std_logic;
signal n12147 : std_logic;
signal n12148 : std_logic;
signal \bfn_3_30_0_\ : std_logic;
signal n12149 : std_logic;
signal n12150 : std_logic;
signal n12151 : std_logic;
signal \bfn_3_31_0_\ : std_logic;
signal n12131 : std_logic;
signal n1299 : std_logic;
signal n12132 : std_logic;
signal n1298 : std_logic;
signal n12133 : std_logic;
signal n12134 : std_logic;
signal n12135 : std_logic;
signal n12136 : std_logic;
signal n12137 : std_logic;
signal n12138 : std_logic;
signal \bfn_3_32_0_\ : std_logic;
signal n12139 : std_logic;
signal n12140 : std_logic;
signal \reg_B_2\ : std_logic;
signal \debounce.n6\ : std_logic;
signal \debounce.reg_A_2\ : std_logic;
signal \debounce.cnt_next_9__N_418\ : std_logic;
signal n1193 : std_logic;
signal n2198 : std_logic;
signal \n2230_cascade_\ : std_logic;
signal n2189 : std_logic;
signal \n2221_cascade_\ : std_logic;
signal \n2320_cascade_\ : std_logic;
signal n2387 : std_logic;
signal n2399 : std_logic;
signal n2397 : std_logic;
signal \n2429_cascade_\ : std_logic;
signal \n14210_cascade_\ : std_logic;
signal \n14214_cascade_\ : std_logic;
signal n13423 : std_logic;
signal n2396 : std_logic;
signal n2329 : std_logic;
signal \n14016_cascade_\ : std_logic;
signal \n14022_cascade_\ : std_logic;
signal n2395 : std_logic;
signal \n2346_cascade_\ : std_logic;
signal n2384 : std_logic;
signal n2385 : std_logic;
signal n2389 : std_logic;
signal n2317 : std_logic;
signal n14410 : std_logic;
signal \n11774_cascade_\ : std_logic;
signal \n14188_cascade_\ : std_logic;
signal n2187 : std_logic;
signal \n2219_cascade_\ : std_logic;
signal n2318 : std_logic;
signal n2330 : std_logic;
signal n2099 : std_logic;
signal n1997 : std_logic;
signal n2029 : std_logic;
signal n2030 : std_logic;
signal \n2029_cascade_\ : std_logic;
signal n14154 : std_logic;
signal n1990 : std_logic;
signal n1923 : std_logic;
signal n2022 : std_logic;
signal \n2022_cascade_\ : std_logic;
signal n14146 : std_logic;
signal n14152 : std_logic;
signal n1928 : std_logic;
signal n1995 : std_logic;
signal n2027 : std_logic;
signal n2023 : std_logic;
signal n2090 : std_logic;
signal n2122 : std_logic;
signal n2128 : std_logic;
signal \n2122_cascade_\ : std_logic;
signal n1918 : std_logic;
signal n1919 : std_logic;
signal n1926 : std_logic;
signal \n1950_cascade_\ : std_logic;
signal n1993 : std_logic;
signal n1999 : std_logic;
signal n2031 : std_logic;
signal \n2031_cascade_\ : std_logic;
signal n11680 : std_logic;
signal n1992 : std_logic;
signal n1925 : std_logic;
signal n1819 : std_logic;
signal n14134 : std_logic;
signal \n1851_cascade_\ : std_logic;
signal n1895 : std_logic;
signal n1927 : std_logic;
signal n1890 : std_logic;
signal n1922 : std_logic;
signal n13772 : std_logic;
signal \n1922_cascade_\ : std_logic;
signal n13770 : std_logic;
signal n1920 : std_logic;
signal \n13778_cascade_\ : std_logic;
signal n13782 : std_logic;
signal \bfn_4_24_0_\ : std_logic;
signal n1733 : std_logic;
signal n1800 : std_logic;
signal n12191 : std_logic;
signal n1732 : std_logic;
signal n1799 : std_logic;
signal n12192 : std_logic;
signal n1731 : std_logic;
signal n1798 : std_logic;
signal n12193 : std_logic;
signal n1730 : std_logic;
signal n1797 : std_logic;
signal n12194 : std_logic;
signal n12195 : std_logic;
signal n1728 : std_logic;
signal n1795 : std_logic;
signal n12196 : std_logic;
signal n1727 : std_logic;
signal n1794 : std_logic;
signal n12197 : std_logic;
signal n12198 : std_logic;
signal \bfn_4_25_0_\ : std_logic;
signal n1725 : std_logic;
signal n1792 : std_logic;
signal n12199 : std_logic;
signal n12200 : std_logic;
signal n1723 : std_logic;
signal n1790 : std_logic;
signal n12201 : std_logic;
signal n1722 : std_logic;
signal n1789 : std_logic;
signal n12202 : std_logic;
signal n1721 : std_logic;
signal n1788 : std_logic;
signal n12203 : std_logic;
signal n1720 : std_logic;
signal n1787 : std_logic;
signal n12204 : std_logic;
signal n1719 : std_logic;
signal n12205 : std_logic;
signal n1601 : std_logic;
signal \bfn_4_26_0_\ : std_logic;
signal n1533 : std_logic;
signal n1600 : std_logic;
signal n12164 : std_logic;
signal n1532 : std_logic;
signal n1599 : std_logic;
signal n12165 : std_logic;
signal n1531 : std_logic;
signal n1598 : std_logic;
signal n12166 : std_logic;
signal n1530 : std_logic;
signal n1597 : std_logic;
signal n12167 : std_logic;
signal n1529 : std_logic;
signal n1596 : std_logic;
signal n12168 : std_logic;
signal n1528 : std_logic;
signal n1595 : std_logic;
signal n12169 : std_logic;
signal n1527 : std_logic;
signal n1594 : std_logic;
signal n12170 : std_logic;
signal n12171 : std_logic;
signal n1593 : std_logic;
signal \bfn_4_27_0_\ : std_logic;
signal n1592 : std_logic;
signal n12172 : std_logic;
signal n1591 : std_logic;
signal n12173 : std_logic;
signal n1523 : std_logic;
signal n1590 : std_logic;
signal n12174 : std_logic;
signal n1522 : std_logic;
signal n1589 : std_logic;
signal n12175 : std_logic;
signal n1521 : std_logic;
signal n12176 : std_logic;
signal n1620 : std_logic;
signal n1427 : std_logic;
signal n1494 : std_logic;
signal n1526 : std_logic;
signal n1493 : std_logic;
signal n1525 : std_logic;
signal n1396 : std_logic;
signal n1428 : std_logic;
signal n1393 : std_logic;
signal n1394 : std_logic;
signal n1426 : std_logic;
signal n1399 : std_logic;
signal n1431 : std_logic;
signal n1391 : std_logic;
signal n1423 : std_logic;
signal n1422 : std_logic;
signal n13334 : std_logic;
signal \n1423_cascade_\ : std_logic;
signal n14094 : std_logic;
signal n1425 : std_logic;
signal \n1455_cascade_\ : std_logic;
signal n1492 : std_logic;
signal n1524 : std_logic;
signal n1301 : std_logic;
signal n1333 : std_logic;
signal \n1333_cascade_\ : std_logic;
signal \n11640_cascade_\ : std_logic;
signal n1331 : std_logic;
signal n1323 : std_logic;
signal \n13315_cascade_\ : std_logic;
signal \n1356_cascade_\ : std_logic;
signal n1392 : std_logic;
signal n1424 : std_logic;
signal n299 : std_logic;
signal n1330 : std_logic;
signal n1397 : std_logic;
signal n1429 : std_logic;
signal n1297 : std_logic;
signal n1329 : std_logic;
signal n1295 : std_logic;
signal n1294 : std_logic;
signal n1224 : std_logic;
signal \n1257_cascade_\ : std_logic;
signal n1201 : std_logic;
signal n1300 : std_logic;
signal \n1233_cascade_\ : std_logic;
signal n1332 : std_logic;
signal n1296 : std_logic;
signal n1194 : std_logic;
signal n1200 : std_logic;
signal n1225 : std_logic;
signal n1292 : std_logic;
signal n1324 : std_logic;
signal \n1158_cascade_\ : std_logic;
signal n1199 : std_logic;
signal n1197 : std_logic;
signal n1130 : std_logic;
signal \n1130_cascade_\ : std_logic;
signal n14068 : std_logic;
signal n11706 : std_logic;
signal \n2527_cascade_\ : std_logic;
signal n13798 : std_logic;
signal \n13796_cascade_\ : std_logic;
signal \n14354_cascade_\ : std_logic;
signal n14220 : std_logic;
signal \n14224_cascade_\ : std_logic;
signal \n2445_cascade_\ : std_logic;
signal \n2517_cascade_\ : std_logic;
signal n13804 : std_logic;
signal n2185 : std_logic;
signal n2390 : std_logic;
signal n2401 : std_logic;
signal \n2433_cascade_\ : std_logic;
signal n11670 : std_logic;
signal n2383 : std_logic;
signal n2314 : std_logic;
signal n2381 : std_logic;
signal \n2314_cascade_\ : std_logic;
signal \n2326_cascade_\ : std_logic;
signal n2393 : std_logic;
signal n2400 : std_logic;
signal n14194 : std_logic;
signal \n2247_cascade_\ : std_logic;
signal n2333 : std_logic;
signal n2332 : std_logic;
signal \n2333_cascade_\ : std_logic;
signal n2331 : std_logic;
signal n11766 : std_logic;
signal n2190 : std_logic;
signal n2133 : std_logic;
signal n2129 : std_logic;
signal n2130 : std_logic;
signal \n11616_cascade_\ : std_logic;
signal n2131 : std_logic;
signal n2001 : std_logic;
signal n2033 : std_logic;
signal n2100 : std_logic;
signal \n2033_cascade_\ : std_logic;
signal n2132 : std_logic;
signal n2199 : std_logic;
signal \n2132_cascade_\ : std_logic;
signal n2000 : std_logic;
signal n2032 : std_logic;
signal n2091 : std_logic;
signal n2024 : std_logic;
signal n2123 : std_logic;
signal \n2123_cascade_\ : std_logic;
signal n2121 : std_logic;
signal \n13746_cascade_\ : std_logic;
signal n13748 : std_logic;
signal n2119 : std_logic;
signal \n13754_cascade_\ : std_logic;
signal n13382 : std_logic;
signal n13760 : std_logic;
signal n1822 : std_logic;
signal n1889 : std_logic;
signal n1921 : std_logic;
signal n1900 : std_logic;
signal n1932 : std_logic;
signal \n1932_cascade_\ : std_logic;
signal n1931 : std_logic;
signal n11686 : std_logic;
signal n1897 : std_logic;
signal n1929 : std_logic;
signal \n1929_cascade_\ : std_logic;
signal n14136 : std_logic;
signal n1901 : std_logic;
signal n1933 : std_logic;
signal n1898 : std_logic;
signal n1930 : std_logic;
signal n1885 : std_logic;
signal n1818 : std_logic;
signal n1917 : std_logic;
signal n1791 : std_logic;
signal n1724 : std_logic;
signal n1823 : std_logic;
signal n1824 : std_logic;
signal \n1823_cascade_\ : std_logic;
signal n1830 : std_logic;
signal n1829 : std_logic;
signal \n14126_cascade_\ : std_logic;
signal n14128 : std_logic;
signal n1793 : std_logic;
signal n1726 : std_logic;
signal n1825 : std_logic;
signal n1827 : std_logic;
signal n1826 : std_logic;
signal \n1825_cascade_\ : std_logic;
signal n14122 : std_logic;
signal n1729 : std_logic;
signal n1796 : std_logic;
signal n1828 : std_logic;
signal n1832 : std_logic;
signal n1831 : std_logic;
signal n11688 : std_logic;
signal n2021 : std_logic;
signal n2088 : std_logic;
signal n2120 : std_logic;
signal n301 : std_logic;
signal n1801 : std_logic;
signal n303 : std_logic;
signal n1833 : std_logic;
signal n307 : std_logic;
signal n13490 : std_logic;
signal n306 : std_logic;
signal \n13257_cascade_\ : std_logic;
signal n302 : std_logic;
signal \bfn_5_28_0_\ : std_logic;
signal n12096 : std_logic;
signal n12097 : std_logic;
signal n2287 : std_logic;
signal n12098 : std_logic;
signal n12099 : std_logic;
signal n402 : std_logic;
signal n12100 : std_logic;
signal n2289 : std_logic;
signal \n13261_cascade_\ : std_logic;
signal n297 : std_logic;
signal \debounce.reg_A_1\ : std_logic;
signal \reg_B_1\ : std_logic;
signal \debounce.reg_A_0\ : std_logic;
signal \reg_B_0\ : std_logic;
signal n2288 : std_logic;
signal n1293 : std_logic;
signal n1325 : std_logic;
signal n1326 : std_logic;
signal n1327 : std_logic;
signal \n1325_cascade_\ : std_logic;
signal n1328 : std_logic;
signal n13734 : std_logic;
signal n298 : std_logic;
signal n1233 : std_logic;
signal \n298_cascade_\ : std_logic;
signal n1232 : std_logic;
signal n1196 : std_logic;
signal n1228 : std_logic;
signal \n1228_cascade_\ : std_logic;
signal n1226 : std_logic;
signal n14078 : std_logic;
signal n1132 : std_logic;
signal n1129 : std_logic;
signal n1133 : std_logic;
signal n1195 : std_logic;
signal n1227 : std_logic;
signal n1198 : std_logic;
signal n1230 : std_logic;
signal n1229 : std_logic;
signal n1231 : std_logic;
signal \n1230_cascade_\ : std_logic;
signal n11642 : std_logic;
signal n13318 : std_logic;
signal n1125 : std_logic;
signal n1126 : std_logic;
signal \n1126_cascade_\ : std_logic;
signal n1127 : std_logic;
signal n13994 : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal n12339 : std_logic;
signal n12340 : std_logic;
signal n12341 : std_logic;
signal n12342 : std_logic;
signal n12343 : std_logic;
signal n12344 : std_logic;
signal n12345 : std_logic;
signal n12346 : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal n12347 : std_logic;
signal n12348 : std_logic;
signal n12349 : std_logic;
signal n12350 : std_logic;
signal n12351 : std_logic;
signal n12352 : std_logic;
signal n12353 : std_logic;
signal n12354 : std_logic;
signal \bfn_6_16_0_\ : std_logic;
signal n12355 : std_logic;
signal n12356 : std_logic;
signal n12357 : std_logic;
signal n2581 : std_logic;
signal n12358 : std_logic;
signal n12359 : std_logic;
signal n12360 : std_logic;
signal n12361 : std_logic;
signal \bfn_6_17_0_\ : std_logic;
signal n12317 : std_logic;
signal n12318 : std_logic;
signal n12319 : std_logic;
signal n2430 : std_logic;
signal n2497 : std_logic;
signal n12320 : std_logic;
signal n2429 : std_logic;
signal n2496 : std_logic;
signal n12321 : std_logic;
signal n2428 : std_logic;
signal n2495 : std_logic;
signal n12322 : std_logic;
signal n2427 : std_logic;
signal n2494 : std_logic;
signal n12323 : std_logic;
signal n12324 : std_logic;
signal n2493 : std_logic;
signal \bfn_6_18_0_\ : std_logic;
signal n12325 : std_logic;
signal n12326 : std_logic;
signal n2490 : std_logic;
signal n12327 : std_logic;
signal n2422 : std_logic;
signal n2489 : std_logic;
signal n12328 : std_logic;
signal n12329 : std_logic;
signal n12330 : std_logic;
signal n2419 : std_logic;
signal n2486 : std_logic;
signal n12331 : std_logic;
signal n12332 : std_logic;
signal n2418 : std_logic;
signal n2485 : std_logic;
signal \bfn_6_19_0_\ : std_logic;
signal n12333 : std_logic;
signal n12334 : std_logic;
signal n2415 : std_logic;
signal n2482 : std_logic;
signal n12335 : std_logic;
signal n12336 : std_logic;
signal n12337 : std_logic;
signal n2412 : std_logic;
signal n12338 : std_logic;
signal n2421 : std_logic;
signal n2488 : std_logic;
signal n2126 : std_logic;
signal n2193 : std_logic;
signal n2192 : std_logic;
signal n2125 : std_logic;
signal \n2224_cascade_\ : std_logic;
signal \n14174_cascade_\ : std_logic;
signal \n14178_cascade_\ : std_logic;
signal n14184 : std_logic;
signal n2500 : std_logic;
signal n2433 : std_logic;
signal n2431 : std_logic;
signal n2498 : std_logic;
signal n2194 : std_logic;
signal n2127 : std_logic;
signal n2501 : std_logic;
signal \n2533_cascade_\ : std_logic;
signal \n11682_cascade_\ : std_logic;
signal n13397 : std_logic;
signal n2086 : std_logic;
signal n2019 : std_logic;
signal n2118 : std_logic;
signal n2432 : std_logic;
signal n2499 : std_logic;
signal n2025 : std_logic;
signal n2092 : std_logic;
signal n2124 : std_logic;
signal n2191 : std_logic;
signal \n2124_cascade_\ : std_logic;
signal \n2223_cascade_\ : std_logic;
signal n2315 : std_logic;
signal n2382 : std_logic;
signal \n2315_cascade_\ : std_logic;
signal n2414 : std_logic;
signal \n2414_cascade_\ : std_logic;
signal n2481 : std_logic;
signal \bfn_6_23_0_\ : std_logic;
signal \quad_counter0.n12623\ : std_logic;
signal \quad_counter0.n12624\ : std_logic;
signal \quad_counter0.n12625\ : std_logic;
signal \quad_counter0.n12626\ : std_logic;
signal \quad_counter0.n12627\ : std_logic;
signal \quad_counter0.n12628\ : std_logic;
signal \quad_counter0.n12629\ : std_logic;
signal \quad_counter0.n12630\ : std_logic;
signal \bfn_6_24_0_\ : std_logic;
signal \quad_counter0.n12631\ : std_logic;
signal \quad_counter0.n12632\ : std_logic;
signal \quad_counter0.n12633\ : std_logic;
signal encoder0_position_12 : std_logic;
signal \quad_counter0.n12634\ : std_logic;
signal \quad_counter0.n12635\ : std_logic;
signal \quad_counter0.n12636\ : std_logic;
signal \quad_counter0.n12637\ : std_logic;
signal \quad_counter0.n12638\ : std_logic;
signal \bfn_6_25_0_\ : std_logic;
signal encoder0_position_17 : std_logic;
signal \quad_counter0.n12639\ : std_logic;
signal encoder0_position_18 : std_logic;
signal \quad_counter0.n12640\ : std_logic;
signal encoder0_position_19 : std_logic;
signal \quad_counter0.n12641\ : std_logic;
signal encoder0_position_20 : std_logic;
signal \quad_counter0.n12642\ : std_logic;
signal encoder0_position_21 : std_logic;
signal \quad_counter0.n12643\ : std_logic;
signal encoder0_position_22 : std_logic;
signal \quad_counter0.n12644\ : std_logic;
signal \quad_counter0.n12645\ : std_logic;
signal \quad_counter0.n12646\ : std_logic;
signal \bfn_6_26_0_\ : std_logic;
signal \quad_counter0.n12647\ : std_logic;
signal \quad_counter0.n12648\ : std_logic;
signal \quad_counter0.n12649\ : std_logic;
signal \quad_counter0.n12650\ : std_logic;
signal \quad_counter0.n12651\ : std_logic;
signal \quad_counter0.n12652\ : std_logic;
signal \quad_counter0.n12653\ : std_logic;
signal encoder0_position_16 : std_logic;
signal encoder0_position_27 : std_logic;
signal n175 : std_logic;
signal encoder0_position_29 : std_logic;
signal n404 : std_logic;
signal \n14170_cascade_\ : std_logic;
signal n2285 : std_logic;
signal n293 : std_logic;
signal \n293_cascade_\ : std_logic;
signal n5_adj_697 : std_logic;
signal \n5_adj_697_cascade_\ : std_logic;
signal n2290 : std_logic;
signal \n13254_cascade_\ : std_logic;
signal n13259 : std_logic;
signal n13263 : std_logic;
signal n174 : std_logic;
signal n13254 : std_logic;
signal n2286 : std_logic;
signal \n13255_cascade_\ : std_logic;
signal encoder0_position_26 : std_logic;
signal encoder0_position_30 : std_logic;
signal n403 : std_logic;
signal \n11712_cascade_\ : std_logic;
signal \n861_cascade_\ : std_logic;
signal encoder0_position_24 : std_logic;
signal n1101 : std_logic;
signal \bfn_6_31_0_\ : std_logic;
signal n1100 : std_logic;
signal n12114 : std_logic;
signal n12115 : std_logic;
signal n1098 : std_logic;
signal n12116 : std_logic;
signal n1097 : std_logic;
signal n12117 : std_logic;
signal n12118 : std_logic;
signal n1095 : std_logic;
signal n12119 : std_logic;
signal n1094 : std_logic;
signal n12120 : std_logic;
signal n12121 : std_logic;
signal \bfn_6_32_0_\ : std_logic;
signal n1093 : std_logic;
signal n1096 : std_logic;
signal n1128 : std_logic;
signal n1028 : std_logic;
signal n1027 : std_logic;
signal \n1059_cascade_\ : std_logic;
signal n1099 : std_logic;
signal n1131 : std_logic;
signal encoder0_position_23 : std_logic;
signal n2590 : std_logic;
signal n2592 : std_logic;
signal n2525 : std_logic;
signal n2517 : std_logic;
signal n2584 : std_logic;
signal n2595 : std_logic;
signal n2528 : std_logic;
signal n2491 : std_logic;
signal n2424 : std_logic;
signal n2523 : std_logic;
signal n2583 : std_logic;
signal n2596 : std_logic;
signal n2529 : std_logic;
signal \n2628_cascade_\ : std_logic;
signal n2585 : std_logic;
signal n2518 : std_logic;
signal n2417 : std_logic;
signal n2484 : std_logic;
signal n2516 : std_logic;
signal n2514 : std_logic;
signal \n2516_cascade_\ : std_logic;
signal n13810 : std_logic;
signal \n13816_cascade_\ : std_logic;
signal n2511 : std_logic;
signal n2582 : std_logic;
signal \n2544_cascade_\ : std_logic;
signal n2579 : std_logic;
signal n2425 : std_logic;
signal n2492 : std_logic;
signal n2524 : std_logic;
signal n2591 : std_logic;
signal \n2524_cascade_\ : std_logic;
signal n2391 : std_logic;
signal n2423 : std_logic;
signal n2601 : std_logic;
signal n2394 : std_logic;
signal n2426 : std_logic;
signal n2480 : std_logic;
signal n2413 : std_logic;
signal n2512 : std_logic;
signal n2388 : std_logic;
signal n2420 : std_logic;
signal n2487 : std_logic;
signal \n2420_cascade_\ : std_logic;
signal n2519 : std_logic;
signal \n2519_cascade_\ : std_logic;
signal n2586 : std_logic;
signal n2532 : std_logic;
signal n2599 : std_logic;
signal n2483 : std_logic;
signal n2416 : std_logic;
signal n2515 : std_logic;
signal n2301 : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal n2233 : std_logic;
signal n2300 : std_logic;
signal n12276 : std_logic;
signal n2232 : std_logic;
signal n2299 : std_logic;
signal n12277 : std_logic;
signal n2231 : std_logic;
signal n2298 : std_logic;
signal n12278 : std_logic;
signal n2230 : std_logic;
signal n2297 : std_logic;
signal n12279 : std_logic;
signal n2229 : std_logic;
signal n2296 : std_logic;
signal n12280 : std_logic;
signal n12281 : std_logic;
signal n2227 : std_logic;
signal n2294 : std_logic;
signal n12282 : std_logic;
signal n12283 : std_logic;
signal n2226 : std_logic;
signal n2293 : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal n12284 : std_logic;
signal n12285 : std_logic;
signal n2223 : std_logic;
signal n2290_adj_604 : std_logic;
signal n12286 : std_logic;
signal n2222 : std_logic;
signal n2289_adj_603 : std_logic;
signal n12287 : std_logic;
signal n2221 : std_logic;
signal n2288_adj_602 : std_logic;
signal n12288 : std_logic;
signal n2220 : std_logic;
signal n2287_adj_601 : std_logic;
signal n12289 : std_logic;
signal n2219 : std_logic;
signal n2286_adj_600 : std_logic;
signal n12290 : std_logic;
signal n12291 : std_logic;
signal n2218 : std_logic;
signal n2285_adj_599 : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal n12292 : std_logic;
signal n2216 : std_logic;
signal n2283 : std_logic;
signal n12293 : std_logic;
signal n2215 : std_logic;
signal n2282 : std_logic;
signal n12294 : std_logic;
signal n2214 : std_logic;
signal n12295 : std_logic;
signal n2313 : std_logic;
signal n2225 : std_logic;
signal n2292 : std_logic;
signal n2224 : std_logic;
signal n2291 : std_logic;
signal n2295 : std_logic;
signal n2228 : std_logic;
signal encoder0_position_2 : std_logic;
signal n2321 : std_logic;
signal n2324 : std_logic;
signal n2328 : std_logic;
signal n2327 : std_logic;
signal n2322 : std_logic;
signal n2326 : std_logic;
signal n2325 : std_logic;
signal n2323 : std_logic;
signal encoder0_position_3 : std_logic;
signal encoder0_position_11 : std_logic;
signal n308 : std_logic;
signal encoder0_position_8 : std_logic;
signal n311 : std_logic;
signal encoder0_position_5 : std_logic;
signal encoder0_position_15 : std_logic;
signal n304 : std_logic;
signal n2320 : std_logic;
signal n2319 : std_logic;
signal n14008 : std_logic;
signal n14006 : std_logic;
signal n14014 : std_logic;
signal encoder0_position_1 : std_logic;
signal encoder0_position_0 : std_logic;
signal n33_adj_657 : std_logic;
signal n33 : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal n32_adj_656 : std_logic;
signal n32 : std_logic;
signal n12575 : std_logic;
signal n31_adj_655 : std_logic;
signal n31 : std_logic;
signal n12576 : std_logic;
signal n30_adj_654 : std_logic;
signal n30 : std_logic;
signal n12577 : std_logic;
signal n29_adj_653 : std_logic;
signal n12578 : std_logic;
signal n28_adj_652 : std_logic;
signal n28 : std_logic;
signal n12579 : std_logic;
signal n27 : std_logic;
signal n12580 : std_logic;
signal n26_adj_650 : std_logic;
signal n12581 : std_logic;
signal n12582 : std_logic;
signal n25_adj_649 : std_logic;
signal n25 : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal n24_adj_648 : std_logic;
signal n12583 : std_logic;
signal n23_adj_647 : std_logic;
signal n12584 : std_logic;
signal n22_adj_646 : std_logic;
signal n22 : std_logic;
signal n12585 : std_logic;
signal n21_adj_645 : std_logic;
signal n21 : std_logic;
signal n12586 : std_logic;
signal n20 : std_logic;
signal n12587 : std_logic;
signal n19_adj_643 : std_logic;
signal n12588 : std_logic;
signal n18_adj_642 : std_logic;
signal n18 : std_logic;
signal n12589 : std_logic;
signal n12590 : std_logic;
signal n17_adj_641 : std_logic;
signal n17 : std_logic;
signal \bfn_7_27_0_\ : std_logic;
signal n16_adj_640 : std_logic;
signal n16 : std_logic;
signal n12591 : std_logic;
signal n15_adj_639 : std_logic;
signal n15 : std_logic;
signal n12592 : std_logic;
signal n14_adj_638 : std_logic;
signal n14 : std_logic;
signal n12593 : std_logic;
signal n13_adj_637 : std_logic;
signal n13 : std_logic;
signal n12594 : std_logic;
signal n12_adj_636 : std_logic;
signal n12 : std_logic;
signal n12595 : std_logic;
signal n11_adj_635 : std_logic;
signal n11 : std_logic;
signal n12596 : std_logic;
signal n10_adj_634 : std_logic;
signal n10 : std_logic;
signal n12597 : std_logic;
signal n12598 : std_logic;
signal n9_adj_633 : std_logic;
signal n9 : std_logic;
signal \bfn_7_28_0_\ : std_logic;
signal n8_adj_632 : std_logic;
signal n12599 : std_logic;
signal n7_adj_631 : std_logic;
signal n7 : std_logic;
signal n12600 : std_logic;
signal n6_adj_630 : std_logic;
signal n6 : std_logic;
signal n12601 : std_logic;
signal n5 : std_logic;
signal n12602 : std_logic;
signal n4_adj_628 : std_logic;
signal n4 : std_logic;
signal n12603 : std_logic;
signal n3_adj_627 : std_logic;
signal n3_adj_567 : std_logic;
signal n12604 : std_logic;
signal n12605 : std_logic;
signal n2_adj_568 : std_logic;
signal n901 : std_logic;
signal \bfn_7_29_0_\ : std_logic;
signal n12101 : std_logic;
signal n832 : std_logic;
signal n899 : std_logic;
signal n12102 : std_logic;
signal n12103 : std_logic;
signal n830 : std_logic;
signal n897 : std_logic;
signal n12104 : std_logic;
signal n829 : std_logic;
signal n896 : std_logic;
signal n12105 : std_logic;
signal n828 : std_logic;
signal n12106 : std_logic;
signal n900 : std_logic;
signal n833 : std_logic;
signal \bfn_7_30_0_\ : std_logic;
signal n12107 : std_logic;
signal n12108 : std_logic;
signal n12109 : std_logic;
signal n12110 : std_logic;
signal n996 : std_logic;
signal n12111 : std_logic;
signal n995 : std_logic;
signal n12112 : std_logic;
signal n12113 : std_logic;
signal n1026 : std_logic;
signal n997 : std_logic;
signal n999 : std_logic;
signal n932 : std_logic;
signal n898 : std_logic;
signal n831 : std_logic;
signal n861 : std_logic;
signal n930 : std_logic;
signal \n930_cascade_\ : std_logic;
signal n929 : std_logic;
signal n927 : std_logic;
signal n928 : std_logic;
signal \n13726_cascade_\ : std_logic;
signal n11710 : std_logic;
signal n1000 : std_logic;
signal \n960_cascade_\ : std_logic;
signal n933 : std_logic;
signal n295 : std_logic;
signal n1001 : std_logic;
signal n931 : std_logic;
signal n960 : std_logic;
signal n998 : std_logic;
signal n1032 : std_logic;
signal n296 : std_logic;
signal n1033 : std_logic;
signal n1031 : std_logic;
signal n1029 : std_logic;
signal \n11646_cascade_\ : std_logic;
signal n1030 : std_logic;
signal n13323 : std_logic;
signal n2531 : std_logic;
signal n2598 : std_logic;
signal \n2630_cascade_\ : std_logic;
signal \n14288_cascade_\ : std_logic;
signal n2527 : std_logic;
signal n2594 : std_logic;
signal \n2626_cascade_\ : std_logic;
signal n14278 : std_logic;
signal \n14280_cascade_\ : std_logic;
signal n14286 : std_logic;
signal n2522 : std_logic;
signal n2589 : std_logic;
signal n2597 : std_logic;
signal n2530 : std_logic;
signal n2520 : std_logic;
signal n2587 : std_logic;
signal n2580 : std_logic;
signal n2513 : std_logic;
signal \n2721_cascade_\ : std_logic;
signal n2526 : std_logic;
signal n2593 : std_logic;
signal \n2625_cascade_\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal n12362 : std_logic;
signal n12363 : std_logic;
signal n12364 : std_logic;
signal n12365 : std_logic;
signal n12366 : std_logic;
signal n12367 : std_logic;
signal n12368 : std_logic;
signal n12369 : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal n2625 : std_logic;
signal n2692 : std_logic;
signal n12370 : std_logic;
signal n12371 : std_logic;
signal n12372 : std_logic;
signal n2622 : std_logic;
signal n2689 : std_logic;
signal n12373 : std_logic;
signal n12374 : std_logic;
signal n12375 : std_logic;
signal n12376 : std_logic;
signal n12377 : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal n12378 : std_logic;
signal n12379 : std_logic;
signal n12380 : std_logic;
signal n12381 : std_logic;
signal n12382 : std_logic;
signal n12383 : std_logic;
signal n12384 : std_logic;
signal n12385 : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \n11750_cascade_\ : std_logic;
signal \n13900_cascade_\ : std_logic;
signal \n3232_cascade_\ : std_logic;
signal n13906 : std_logic;
signal \n13912_cascade_\ : std_logic;
signal \n3138_cascade_\ : std_logic;
signal \n3229_cascade_\ : std_logic;
signal n11658 : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal n12552 : std_logic;
signal n12553 : std_logic;
signal n12554 : std_logic;
signal n12555 : std_logic;
signal n12556 : std_logic;
signal n12557 : std_logic;
signal n15437 : std_logic;
signal n12558 : std_logic;
signal n12559 : std_logic;
signal n15401 : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal n15375 : std_logic;
signal n2445 : std_logic;
signal n12560 : std_logic;
signal n15348 : std_logic;
signal n2346 : std_logic;
signal n12561 : std_logic;
signal n15322 : std_logic;
signal n12562 : std_logic;
signal n15059 : std_logic;
signal n2148 : std_logic;
signal n12563 : std_logic;
signal n15035 : std_logic;
signal n2049 : std_logic;
signal n12564 : std_logic;
signal n15012 : std_logic;
signal n1950 : std_logic;
signal n12565 : std_logic;
signal n14990 : std_logic;
signal n1851 : std_logic;
signal n12566 : std_logic;
signal n12567 : std_logic;
signal n14969 : std_logic;
signal n1752 : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal n14949 : std_logic;
signal n1653 : std_logic;
signal n12568 : std_logic;
signal n15292 : std_logic;
signal n1554 : std_logic;
signal n12569 : std_logic;
signal n15276 : std_logic;
signal n1455 : std_logic;
signal n12570 : std_logic;
signal n15259 : std_logic;
signal n1356 : std_logic;
signal n12571 : std_logic;
signal n15243 : std_logic;
signal n1257 : std_logic;
signal n12572 : std_logic;
signal n15224 : std_logic;
signal n1158 : std_logic;
signal n12573 : std_logic;
signal n2_adj_626 : std_logic;
signal n12574 : std_logic;
signal encoder0_position_scaled_17 : std_logic;
signal encoder0_position_scaled_20 : std_logic;
signal encoder0_position_25 : std_logic;
signal n8 : std_logic;
signal n294 : std_logic;
signal encoder0_position_scaled_23 : std_logic;
signal \ENCODER0_A_N\ : std_logic;
signal n1059 : std_logic;
signal n15210 : std_logic;
signal \n14536_cascade_\ : std_logic;
signal blink_counter_25 : std_logic;
signal \LED_c\ : std_logic;
signal blink_counter_24 : std_logic;
signal blink_counter_21 : std_logic;
signal blink_counter_22 : std_logic;
signal blink_counter_23 : std_logic;
signal n14535 : std_logic;
signal n14294 : std_logic;
signal n2693 : std_logic;
signal n2626 : std_logic;
signal \n2725_cascade_\ : std_logic;
signal \n14040_cascade_\ : std_logic;
signal n2629 : std_logic;
signal n2696 : std_logic;
signal n2630 : std_logic;
signal n2697 : std_logic;
signal n2695 : std_logic;
signal n2628 : std_logic;
signal n2619 : std_logic;
signal n2686 : std_logic;
signal n2627 : std_logic;
signal n2694 : std_logic;
signal n2521 : std_logic;
signal n2588 : std_logic;
signal n2620 : std_logic;
signal n2687 : std_logic;
signal \n2620_cascade_\ : std_logic;
signal n2610 : std_logic;
signal n14300 : std_logic;
signal n2621 : std_logic;
signal \n2643_cascade_\ : std_logic;
signal n2688 : std_logic;
signal \n2720_cascade_\ : std_logic;
signal \n14038_cascade_\ : std_logic;
signal n14042 : std_logic;
signal n2614 : std_logic;
signal n2681 : std_logic;
signal n2685 : std_logic;
signal n2618 : std_logic;
signal encoder0_position_6 : std_logic;
signal n27_adj_651 : std_logic;
signal n24 : std_logic;
signal encoder0_position_9 : std_logic;
signal n310 : std_logic;
signal n19 : std_logic;
signal encoder0_position_14 : std_logic;
signal n305 : std_logic;
signal n23 : std_logic;
signal encoder0_position_10 : std_logic;
signal n309 : std_logic;
signal n2616 : std_logic;
signal n2683 : std_logic;
signal \n13884_cascade_\ : std_logic;
signal \n3117_cascade_\ : std_logic;
signal n13888 : std_logic;
signal n13886 : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal n12437 : std_logic;
signal n12438 : std_logic;
signal n12439 : std_logic;
signal n12440 : std_logic;
signal n12441 : std_logic;
signal n12442 : std_logic;
signal n12443 : std_logic;
signal n12444 : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal n12445 : std_logic;
signal n12446 : std_logic;
signal n12447 : std_logic;
signal n12448 : std_logic;
signal n12449 : std_logic;
signal n12450 : std_logic;
signal n12451 : std_logic;
signal n12452 : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal n12453 : std_logic;
signal n12454 : std_logic;
signal n12455 : std_logic;
signal n12456 : std_logic;
signal n12457 : std_logic;
signal n12458 : std_logic;
signal n12459 : std_logic;
signal n12460 : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal n12461 : std_logic;
signal n12462 : std_logic;
signal n12463 : std_logic;
signal n15197 : std_logic;
signal \n11593_cascade_\ : std_logic;
signal \n59_cascade_\ : std_logic;
signal n11838 : std_logic;
signal encoder0_position_scaled_0 : std_logic;
signal encoder0_position_scaled_15 : std_logic;
signal encoder0_position_scaled_12 : std_logic;
signal encoder0_position_scaled_2 : std_logic;
signal encoder0_position_scaled_4 : std_logic;
signal \dti_N_333_cascade_\ : std_logic;
signal encoder0_position_scaled_22 : std_logic;
signal n26 : std_logic;
signal encoder0_position_7 : std_logic;
signal encoder0_position_scaled_19 : std_logic;
signal encoder0_position_scaled_21 : std_logic;
signal encoder0_position_scaled_13 : std_logic;
signal n4828 : std_logic;
signal encoder0_position_13 : std_logic;
signal n20_adj_644 : std_logic;
signal encoder0_position_28 : std_logic;
signal n5_adj_629 : std_logic;
signal encoder0_position_scaled_9 : std_logic;
signal encoder0_position_scaled_10 : std_logic;
signal h2 : std_logic;
signal h3 : std_logic;
signal h1 : std_logic;
signal n6_adj_592 : std_logic;
signal \commutation_state_7__N_261\ : std_logic;
signal \n41_cascade_\ : std_logic;
signal n41 : std_logic;
signal \n14715_cascade_\ : std_logic;
signal n40 : std_logic;
signal \n14866_cascade_\ : std_logic;
signal \n12_adj_598_cascade_\ : std_logic;
signal \n45_cascade_\ : std_logic;
signal n16_adj_614 : std_logic;
signal \n14843_cascade_\ : std_logic;
signal n24_adj_619 : std_logic;
signal \n14711_cascade_\ : std_logic;
signal n8_adj_607 : std_logic;
signal n45 : std_logic;
signal \n14826_cascade_\ : std_logic;
signal n14779 : std_logic;
signal n14864 : std_logic;
signal n43 : std_logic;
signal n14713 : std_logic;
signal n2700 : std_logic;
signal \n2732_cascade_\ : std_logic;
signal \n11666_cascade_\ : std_logic;
signal n2691 : std_logic;
signal n2624 : std_logic;
signal n2617 : std_logic;
signal n2684 : std_logic;
signal n2701 : std_logic;
signal n2613 : std_logic;
signal n2680 : std_logic;
signal n2611 : std_logic;
signal n2678 : std_logic;
signal n2615 : std_logic;
signal n2682 : std_logic;
signal \n2714_cascade_\ : std_logic;
signal n2623 : std_logic;
signal n2690 : std_logic;
signal n2698 : std_logic;
signal n2699 : std_logic;
signal n2217 : std_logic;
signal n2284 : std_logic;
signal n2247 : std_logic;
signal n2316 : std_logic;
signal n2533 : std_logic;
signal n2600 : std_logic;
signal n2544 : std_logic;
signal n2632 : std_logic;
signal n312 : std_logic;
signal n2633 : std_logic;
signal \n2632_cascade_\ : std_logic;
signal n2631 : std_logic;
signal n11760 : std_logic;
signal \n2817_cascade_\ : std_logic;
signal n3000 : std_logic;
signal \n3032_cascade_\ : std_logic;
signal \n11660_cascade_\ : std_logic;
signal n2986 : std_logic;
signal n2997 : std_logic;
signal \n3029_cascade_\ : std_logic;
signal encoder0_position_31 : std_logic;
signal n29 : std_logic;
signal encoder0_position_4 : std_logic;
signal n3001 : std_logic;
signal \n315_cascade_\ : std_logic;
signal n2998 : std_logic;
signal \n3115_cascade_\ : std_logic;
signal n13894 : std_logic;
signal n13898 : std_logic;
signal n2988 : std_logic;
signal n2987 : std_logic;
signal \n3019_cascade_\ : std_logic;
signal n2983 : std_logic;
signal n2981 : std_logic;
signal n2984 : std_logic;
signal \n2912_cascade_\ : std_logic;
signal n2979 : std_logic;
signal n2975 : std_logic;
signal n2980 : std_logic;
signal n2976 : std_logic;
signal n2978 : std_logic;
signal \n3010_cascade_\ : std_logic;
signal n15090 : std_logic;
signal \n14392_cascade_\ : std_logic;
signal n13470 : std_logic;
signal \n14380_cascade_\ : std_logic;
signal n14386 : std_logic;
signal n14398 : std_logic;
signal \n3237_cascade_\ : std_logic;
signal n61 : std_logic;
signal \n13856_cascade_\ : std_logic;
signal \n13858_cascade_\ : std_logic;
signal \n13860_cascade_\ : std_logic;
signal \n13862_cascade_\ : std_logic;
signal \n13864_cascade_\ : std_logic;
signal n13866 : std_logic;
signal encoder0_position_scaled_5 : std_logic;
signal encoder0_position_scaled_8 : std_logic;
signal encoder0_position_scaled_11 : std_logic;
signal encoder0_position_scaled_7 : std_logic;
signal encoder0_position_scaled_1 : std_logic;
signal \n4_adj_698_cascade_\ : std_logic;
signal pwm_setpoint_21 : std_logic;
signal encoder0_position_scaled_14 : std_logic;
signal encoder0_position_scaled_16 : std_logic;
signal encoder0_position_scaled_18 : std_logic;
signal commutation_state_prev_2 : std_logic;
signal \bfn_11_29_0_\ : std_logic;
signal \PWM.n12686\ : std_logic;
signal \PWM.n12687\ : std_logic;
signal \PWM.n12688\ : std_logic;
signal pwm_counter_4 : std_logic;
signal \PWM.n12689\ : std_logic;
signal \PWM.n12690\ : std_logic;
signal \PWM.n12691\ : std_logic;
signal \PWM.n12692\ : std_logic;
signal \PWM.n12693\ : std_logic;
signal \bfn_11_30_0_\ : std_logic;
signal \PWM.n12694\ : std_logic;
signal \PWM.n12695\ : std_logic;
signal pwm_counter_11 : std_logic;
signal \PWM.n12696\ : std_logic;
signal \PWM.n12697\ : std_logic;
signal \PWM.n12698\ : std_logic;
signal \PWM.n12699\ : std_logic;
signal \PWM.n12700\ : std_logic;
signal \PWM.n12701\ : std_logic;
signal \bfn_11_31_0_\ : std_logic;
signal \PWM.n12702\ : std_logic;
signal \PWM.n12703\ : std_logic;
signal \PWM.n12704\ : std_logic;
signal pwm_counter_20 : std_logic;
signal \PWM.n12705\ : std_logic;
signal pwm_counter_21 : std_logic;
signal \PWM.n12706\ : std_logic;
signal pwm_counter_22 : std_logic;
signal \PWM.n12707\ : std_logic;
signal \PWM.n12708\ : std_logic;
signal \PWM.n12709\ : std_logic;
signal pwm_counter_24 : std_logic;
signal \bfn_11_32_0_\ : std_logic;
signal pwm_counter_25 : std_logic;
signal \PWM.n12710\ : std_logic;
signal pwm_counter_26 : std_logic;
signal \PWM.n12711\ : std_logic;
signal pwm_counter_27 : std_logic;
signal \PWM.n12712\ : std_logic;
signal pwm_counter_28 : std_logic;
signal \PWM.n12713\ : std_logic;
signal pwm_counter_29 : std_logic;
signal \PWM.n12714\ : std_logic;
signal pwm_counter_30 : std_logic;
signal \PWM.n12715\ : std_logic;
signal \PWM.n12716\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal n12386 : std_logic;
signal n12387 : std_logic;
signal n12388 : std_logic;
signal n12389 : std_logic;
signal n12390 : std_logic;
signal n12391 : std_logic;
signal n12392 : std_logic;
signal n12393 : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal n12394 : std_logic;
signal n12395 : std_logic;
signal n12396 : std_logic;
signal n12397 : std_logic;
signal n2721 : std_logic;
signal n2788 : std_logic;
signal n12398 : std_logic;
signal n12399 : std_logic;
signal n12400 : std_logic;
signal n12401 : std_logic;
signal n2718 : std_logic;
signal n2785 : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal n2717 : std_logic;
signal n2784 : std_logic;
signal n12402 : std_logic;
signal n12403 : std_logic;
signal n12404 : std_logic;
signal n2781 : std_logic;
signal n12405 : std_logic;
signal n12406 : std_logic;
signal n12407 : std_logic;
signal n12408 : std_logic;
signal n12409 : std_logic;
signal n2777 : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal n12410 : std_logic;
signal n2985 : std_logic;
signal \n3017_cascade_\ : std_logic;
signal n2977 : std_logic;
signal n2993 : std_logic;
signal n2911 : std_logic;
signal n2912 : std_logic;
signal \n13948_cascade_\ : std_logic;
signal \n13954_cascade_\ : std_logic;
signal n2999 : std_logic;
signal \n2940_cascade_\ : std_logic;
signal n2996 : std_logic;
signal \n14340_cascade_\ : std_logic;
signal n2908 : std_logic;
signal n14344 : std_logic;
signal \n3039_cascade_\ : std_logic;
signal n13466 : std_logic;
signal n14334 : std_logic;
signal \n3121_cascade_\ : std_logic;
signal \n3112_cascade_\ : std_logic;
signal \n23_adj_707_cascade_\ : std_logic;
signal \n25_adj_708_cascade_\ : std_logic;
signal \n13832_cascade_\ : std_logic;
signal n13828 : std_logic;
signal n13826 : std_logic;
signal \n13840_cascade_\ : std_logic;
signal n13846 : std_logic;
signal \n13848_cascade_\ : std_logic;
signal n5_adj_713 : std_logic;
signal \n13850_cascade_\ : std_logic;
signal n11656 : std_logic;
signal \n13852_cascade_\ : std_logic;
signal n13854 : std_logic;
signal n37_adj_710 : std_logic;
signal n7_adj_703 : std_logic;
signal \n14_adj_679_cascade_\ : std_logic;
signal \n4781_cascade_\ : std_logic;
signal n14700 : std_logic;
signal n1259 : std_logic;
signal dti_counter_0 : std_logic;
signal \bfn_12_27_0_\ : std_logic;
signal n14693 : std_logic;
signal n12742 : std_logic;
signal n14692 : std_logic;
signal n12743 : std_logic;
signal n14691 : std_logic;
signal dti_counter_3 : std_logic;
signal n12744 : std_logic;
signal n14690 : std_logic;
signal dti_counter_4 : std_logic;
signal n12745 : std_logic;
signal n12746 : std_logic;
signal n14688 : std_logic;
signal dti_counter_6 : std_logic;
signal n12747 : std_logic;
signal n14687 : std_logic;
signal n11202 : std_logic;
signal n12748 : std_logic;
signal dti_counter_7 : std_logic;
signal pwm_setpoint_4 : std_logic;
signal pwm_counter_2 : std_logic;
signal pwm_counter_3 : std_logic;
signal pwm_setpoint_3 : std_logic;
signal n4_adj_698 : std_logic;
signal dti_counter_5 : std_logic;
signal commutation_state_prev_0 : std_logic;
signal n14689 : std_logic;
signal pwm_setpoint_2 : std_logic;
signal pwm_setpoint_11 : std_logic;
signal pwm_setpoint_8 : std_logic;
signal pwm_counter_10 : std_logic;
signal \n21_adj_617_cascade_\ : std_logic;
signal n6_adj_606 : std_logic;
signal n14842 : std_logic;
signal pwm_setpoint_10 : std_logic;
signal \n11_adj_610_cascade_\ : std_logic;
signal pwm_setpoint_5 : std_logic;
signal pwm_setpoint_6 : std_logic;
signal n4825 : std_logic;
signal n13_adj_612 : std_logic;
signal n11_adj_610 : std_logic;
signal n14745 : std_logic;
signal pwm_setpoint_20 : std_logic;
signal pwm_counter_5 : std_logic;
signal pwm_counter_6 : std_logic;
signal \PWM.n13596_cascade_\ : std_logic;
signal pwm_counter_8 : std_logic;
signal \PWM.n26\ : std_logic;
signal n4823 : std_logic;
signal \PWM.n17_cascade_\ : std_logic;
signal pwm_counter_31 : std_logic;
signal \PWM.n29_cascade_\ : std_logic;
signal \PWM.n27\ : std_logic;
signal \PWM.pwm_counter_31__N_401\ : std_logic;
signal pwm_counter_19 : std_logic;
signal n39 : std_logic;
signal pwm_setpoint_19 : std_logic;
signal \n39_cascade_\ : std_logic;
signal n14883 : std_logic;
signal pwm_counter_9 : std_logic;
signal n14804 : std_logic;
signal \n19_adj_616_cascade_\ : std_logic;
signal n15_adj_613 : std_logic;
signal n23_adj_618 : std_logic;
signal \n14800_cascade_\ : std_logic;
signal n19_adj_616 : std_logic;
signal n17_adj_615 : std_logic;
signal n9_adj_608 : std_logic;
signal n21_adj_617 : std_logic;
signal n14734 : std_logic;
signal n14874 : std_logic;
signal pwm_setpoint_12 : std_logic;
signal pwm_counter_12 : std_logic;
signal n25_adj_620 : std_logic;
signal n2723 : std_logic;
signal n2790 : std_logic;
signal n2725 : std_logic;
signal n2792 : std_logic;
signal n13403 : std_logic;
signal n14048 : std_logic;
signal n2714 : std_logic;
signal \n14054_cascade_\ : std_logic;
signal n2710 : std_logic;
signal \n14060_cascade_\ : std_logic;
signal n2709 : std_logic;
signal n2798 : std_logic;
signal \n2742_cascade_\ : std_logic;
signal n2731 : std_logic;
signal n2728 : std_logic;
signal n2795 : std_logic;
signal \n14238_cascade_\ : std_logic;
signal \n14240_cascade_\ : std_logic;
signal n2720 : std_logic;
signal n2787 : std_logic;
signal n2789 : std_logic;
signal n2722 : std_logic;
signal n2797 : std_logic;
signal n2730 : std_logic;
signal n2724 : std_logic;
signal n2791 : std_logic;
signal n2786 : std_logic;
signal n2719 : std_logic;
signal n2921 : std_logic;
signal \n2921_cascade_\ : std_logic;
signal n2778 : std_logic;
signal n2917 : std_logic;
signal n2918 : std_logic;
signal n13926 : std_logic;
signal \n2917_cascade_\ : std_logic;
signal n2916 : std_logic;
signal \n13934_cascade_\ : std_logic;
signal n13942 : std_logic;
signal n2679 : std_logic;
signal n2612 : std_logic;
signal n2643 : std_logic;
signal n2711 : std_logic;
signal n15467 : std_logic;
signal n2909 : std_logic;
signal n2713 : std_logic;
signal n2780 : std_logic;
signal \n14322_cascade_\ : std_logic;
signal n14328 : std_logic;
signal n2992 : std_logic;
signal n2991 : std_logic;
signal \n3023_cascade_\ : std_logic;
signal n14320 : std_logic;
signal n2995 : std_logic;
signal n2994 : std_logic;
signal n2913 : std_logic;
signal n2990 : std_logic;
signal n2982 : std_logic;
signal n2915 : std_logic;
signal \n3014_cascade_\ : std_logic;
signal n14408 : std_logic;
signal n2940 : std_logic;
signal n2989 : std_logic;
signal \n3021_cascade_\ : std_logic;
signal n319 : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal n318 : std_logic;
signal n3301 : std_logic;
signal n12521 : std_logic;
signal n3233 : std_logic;
signal n3300 : std_logic;
signal n12522 : std_logic;
signal n3232 : std_logic;
signal n3299 : std_logic;
signal n12523 : std_logic;
signal n3231 : std_logic;
signal n12524 : std_logic;
signal n3298 : std_logic;
signal n3230 : std_logic;
signal n14697 : std_logic;
signal n12525 : std_logic;
signal n12526 : std_logic;
signal n12527 : std_logic;
signal n12528 : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal n3293 : std_logic;
signal n12529 : std_logic;
signal n12530 : std_logic;
signal n3291 : std_logic;
signal n12531 : std_logic;
signal n3290 : std_logic;
signal n12532 : std_logic;
signal n12533 : std_logic;
signal n3288 : std_logic;
signal n12534 : std_logic;
signal n12535 : std_logic;
signal n12536 : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal n3285 : std_logic;
signal n12537 : std_logic;
signal n3217 : std_logic;
signal n3284 : std_logic;
signal n12538 : std_logic;
signal n3216 : std_logic;
signal n3283 : std_logic;
signal n12539 : std_logic;
signal n3215 : std_logic;
signal n3282 : std_logic;
signal n12540 : std_logic;
signal n3214 : std_logic;
signal n3281 : std_logic;
signal n12541 : std_logic;
signal n3280 : std_logic;
signal n12542 : std_logic;
signal n3212 : std_logic;
signal n3279 : std_logic;
signal n12543 : std_logic;
signal n12544 : std_logic;
signal n3211 : std_logic;
signal n3278 : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal n3210 : std_logic;
signal n3277 : std_logic;
signal n12545 : std_logic;
signal n3276 : std_logic;
signal n12546 : std_logic;
signal n3208 : std_logic;
signal n3275 : std_logic;
signal n12547 : std_logic;
signal n3207 : std_logic;
signal n3274 : std_logic;
signal n12548 : std_logic;
signal n3206 : std_logic;
signal n3273 : std_logic;
signal n12549 : std_logic;
signal n3205 : std_logic;
signal n3272 : std_logic;
signal n12550 : std_logic;
signal n15163 : std_logic;
signal n12551 : std_logic;
signal n14461 : std_logic;
signal encoder0_position_scaled_3 : std_logic;
signal dti_counter_2 : std_logic;
signal dti_counter_1 : std_logic;
signal n10_adj_680 : std_logic;
signal n25_adj_591 : std_logic;
signal \bfn_13_28_0_\ : std_logic;
signal n12050 : std_logic;
signal n23_adj_589 : std_logic;
signal \pwm_setpoint_23_N_171_2\ : std_logic;
signal n12051 : std_logic;
signal \pwm_setpoint_23_N_171_3\ : std_logic;
signal n12052 : std_logic;
signal n21_adj_587 : std_logic;
signal \pwm_setpoint_23_N_171_4\ : std_logic;
signal n12053 : std_logic;
signal n20_adj_586 : std_logic;
signal \pwm_setpoint_23_N_171_5\ : std_logic;
signal n12054 : std_logic;
signal n19_adj_585 : std_logic;
signal \pwm_setpoint_23_N_171_6\ : std_logic;
signal n12055 : std_logic;
signal n18_adj_584 : std_logic;
signal n12056 : std_logic;
signal n12057 : std_logic;
signal \pwm_setpoint_23_N_171_8\ : std_logic;
signal \bfn_13_29_0_\ : std_logic;
signal n12058 : std_logic;
signal n15_adj_581 : std_logic;
signal \pwm_setpoint_23_N_171_10\ : std_logic;
signal n12059 : std_logic;
signal n14_adj_580 : std_logic;
signal \pwm_setpoint_23_N_171_11\ : std_logic;
signal n12060 : std_logic;
signal \pwm_setpoint_23_N_171_12\ : std_logic;
signal n12061 : std_logic;
signal n12062 : std_logic;
signal n11_adj_577 : std_logic;
signal n12063 : std_logic;
signal n12064 : std_logic;
signal n12065 : std_logic;
signal \bfn_13_30_0_\ : std_logic;
signal n12066 : std_logic;
signal n12067 : std_logic;
signal \pwm_setpoint_23_N_171_19\ : std_logic;
signal n12068 : std_logic;
signal \pwm_setpoint_23_N_171_20\ : std_logic;
signal n12069 : std_logic;
signal n4_adj_570 : std_logic;
signal \pwm_setpoint_23_N_171_21\ : std_logic;
signal n12070 : std_logic;
signal n12071 : std_logic;
signal n12072 : std_logic;
signal pwm_setpoint_23 : std_logic;
signal \pwm_setpoint_23_N_171_15\ : std_logic;
signal \pwm_setpoint_23_N_171_18\ : std_logic;
signal pwm_counter_23 : std_logic;
signal \PWM.n28\ : std_logic;
signal pwm_counter_15 : std_logic;
signal pwm_counter_18 : std_logic;
signal n37 : std_logic;
signal pwm_setpoint_18 : std_logic;
signal \n37_cascade_\ : std_logic;
signal n14887 : std_logic;
signal \pwm_setpoint_23_N_171_22\ : std_logic;
signal pwm_setpoint_22 : std_logic;
signal \pwm_setpoint_23_N_171_17\ : std_logic;
signal n14870 : std_logic;
signal n14832 : std_logic;
signal pwm_counter_17 : std_logic;
signal n2712 : std_logic;
signal n2779 : std_logic;
signal \n2811_cascade_\ : std_logic;
signal n2794 : std_logic;
signal n2727 : std_logic;
signal n2716 : std_logic;
signal n2783 : std_logic;
signal n2782 : std_logic;
signal n2715 : std_logic;
signal \n2814_cascade_\ : std_logic;
signal n14260 : std_logic;
signal n2796 : std_logic;
signal n2729 : std_logic;
signal n2800 : std_logic;
signal n2733 : std_logic;
signal n2799 : std_logic;
signal n2732 : std_logic;
signal n14246 : std_logic;
signal \n14248_cascade_\ : std_logic;
signal \n14254_cascade_\ : std_logic;
signal n14266 : std_logic;
signal \n2841_cascade_\ : std_logic;
signal n2923 : std_logic;
signal \n13932_cascade_\ : std_logic;
signal n13936 : std_logic;
signal n2926 : std_logic;
signal n2920 : std_logic;
signal n2927 : std_logic;
signal n2919 : std_logic;
signal n2928 : std_logic;
signal n2922 : std_logic;
signal n2793 : std_logic;
signal n2726 : std_logic;
signal \n2825_cascade_\ : std_logic;
signal n2924 : std_logic;
signal n2925 : std_logic;
signal \n3122_cascade_\ : std_logic;
signal n2914 : std_logic;
signal n316 : std_logic;
signal n3101 : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal n3033 : std_logic;
signal n3100 : std_logic;
signal n12464 : std_logic;
signal n3032 : std_logic;
signal n3099 : std_logic;
signal n12465 : std_logic;
signal n3031 : std_logic;
signal n3098 : std_logic;
signal n12466 : std_logic;
signal n3030 : std_logic;
signal n3097 : std_logic;
signal n12467 : std_logic;
signal n3029 : std_logic;
signal n3096 : std_logic;
signal n12468 : std_logic;
signal n3028 : std_logic;
signal n3095 : std_logic;
signal n12469 : std_logic;
signal n3027 : std_logic;
signal n3094 : std_logic;
signal n12470 : std_logic;
signal n12471 : std_logic;
signal n3026 : std_logic;
signal n3093 : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal n3025 : std_logic;
signal n3092 : std_logic;
signal n12472 : std_logic;
signal n3024 : std_logic;
signal n3091 : std_logic;
signal n12473 : std_logic;
signal n3023 : std_logic;
signal n3090 : std_logic;
signal n12474 : std_logic;
signal n3022 : std_logic;
signal n3089 : std_logic;
signal n12475 : std_logic;
signal n3021 : std_logic;
signal n3088 : std_logic;
signal n12476 : std_logic;
signal n3020 : std_logic;
signal n3087 : std_logic;
signal n12477 : std_logic;
signal n3019 : std_logic;
signal n3086 : std_logic;
signal n12478 : std_logic;
signal n12479 : std_logic;
signal n3018 : std_logic;
signal n3085 : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal n3017 : std_logic;
signal n3084 : std_logic;
signal n12480 : std_logic;
signal n3016 : std_logic;
signal n3083 : std_logic;
signal n12481 : std_logic;
signal n12482 : std_logic;
signal n3014 : std_logic;
signal n3081 : std_logic;
signal n12483 : std_logic;
signal n3013 : std_logic;
signal n3080 : std_logic;
signal n12484 : std_logic;
signal n3012 : std_logic;
signal n3079 : std_logic;
signal n12485 : std_logic;
signal n12486 : std_logic;
signal n12487 : std_logic;
signal n3010 : std_logic;
signal n3077 : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal n12488 : std_logic;
signal n3008 : std_logic;
signal n3075 : std_logic;
signal n12489 : std_logic;
signal n3007 : std_logic;
signal n3074 : std_logic;
signal n12490 : std_logic;
signal n3006 : std_logic;
signal n15123 : std_logic;
signal n12491 : std_logic;
signal n3295 : std_logic;
signal n3294 : std_logic;
signal n3221 : std_logic;
signal n3218 : std_logic;
signal \n14368_cascade_\ : std_logic;
signal n14374 : std_logic;
signal n3228 : std_logic;
signal \n3228_cascade_\ : std_logic;
signal n3224 : std_logic;
signal n14362 : std_logic;
signal n3223 : std_logic;
signal n14366 : std_logic;
signal n3227 : std_logic;
signal n25_adj_545 : std_logic;
signal \bfn_14_26_0_\ : std_logic;
signal n24_adj_546 : std_logic;
signal n12073 : std_logic;
signal n23_adj_547 : std_logic;
signal duty_2 : std_logic;
signal n12074 : std_logic;
signal n22_adj_548 : std_logic;
signal n12075 : std_logic;
signal n21_adj_549 : std_logic;
signal duty_4 : std_logic;
signal n12076 : std_logic;
signal n20_adj_550 : std_logic;
signal duty_5 : std_logic;
signal n12077 : std_logic;
signal duty_6 : std_logic;
signal n12078 : std_logic;
signal n18_adj_552 : std_logic;
signal n12079 : std_logic;
signal n12080 : std_logic;
signal n17_adj_553 : std_logic;
signal \bfn_14_27_0_\ : std_logic;
signal n16_adj_554 : std_logic;
signal n12081 : std_logic;
signal n15_adj_555 : std_logic;
signal duty_10 : std_logic;
signal n12082 : std_logic;
signal n14_adj_556 : std_logic;
signal duty_11 : std_logic;
signal n12083 : std_logic;
signal n13_adj_557 : std_logic;
signal n12084 : std_logic;
signal n12_adj_558 : std_logic;
signal n12085 : std_logic;
signal n11_adj_559 : std_logic;
signal n12086 : std_logic;
signal n10_adj_560 : std_logic;
signal n12087 : std_logic;
signal n12088 : std_logic;
signal n9_adj_561 : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal n8_adj_562 : std_logic;
signal n12089 : std_logic;
signal n7_adj_563 : std_logic;
signal n12090 : std_logic;
signal n6_adj_564 : std_logic;
signal n12091 : std_logic;
signal n5_adj_565 : std_logic;
signal n12092 : std_logic;
signal n4_adj_566 : std_logic;
signal duty_21 : std_logic;
signal n12093 : std_logic;
signal n3 : std_logic;
signal n12094 : std_logic;
signal n2 : std_logic;
signal n12095 : std_logic;
signal \pwm_setpoint_23_N_171_13\ : std_logic;
signal duty_15 : std_logic;
signal n10_adj_576 : std_logic;
signal duty_14 : std_logic;
signal \pwm_setpoint_23_N_171_14\ : std_logic;
signal pwm_counter_1 : std_logic;
signal pwm_counter_0 : std_logic;
signal n16_adj_582 : std_logic;
signal duty_13 : std_logic;
signal n12_adj_578 : std_logic;
signal \pwm_setpoint_23_N_171_0\ : std_logic;
signal duty_0 : std_logic;
signal pwm_setpoint_0 : std_logic;
signal duty_12 : std_logic;
signal n13_adj_579 : std_logic;
signal pwm_counter_14 : std_logic;
signal pwm_counter_13 : std_logic;
signal n27_adj_621 : std_logic;
signal pwm_setpoint_13 : std_logic;
signal \n27_adj_621_cascade_\ : std_logic;
signal n4_adj_605 : std_logic;
signal pwm_setpoint_14 : std_logic;
signal \n14840_cascade_\ : std_logic;
signal duty_22 : std_logic;
signal n3_adj_569 : std_logic;
signal n9_adj_575 : std_logic;
signal duty_16 : std_logic;
signal \pwm_setpoint_23_N_171_16\ : std_logic;
signal duty_20 : std_logic;
signal n5_adj_571 : std_logic;
signal pwm_counter_7 : std_logic;
signal n10_adj_609 : std_logic;
signal \n14722_cascade_\ : std_logic;
signal \n14876_cascade_\ : std_logic;
signal n14886 : std_logic;
signal pwm_setpoint_15 : std_logic;
signal n14841 : std_logic;
signal n14781 : std_logic;
signal \pwm_setpoint_23_N_171_7\ : std_logic;
signal duty_7 : std_logic;
signal pwm_setpoint_7 : std_logic;
signal pwm_setpoint_17 : std_logic;
signal \n12_adj_611_cascade_\ : std_logic;
signal n35 : std_logic;
signal n30_adj_623 : std_logic;
signal pwm_setpoint_16 : std_logic;
signal pwm_counter_16 : std_logic;
signal n33_adj_625 : std_logic;
signal n31_adj_624 : std_logic;
signal n14728 : std_logic;
signal \n33_adj_625_cascade_\ : std_logic;
signal n29_adj_622 : std_logic;
signal n14724 : std_logic;
signal duty_17 : std_logic;
signal n8_adj_574 : std_logic;
signal n28_adj_597 : std_logic;
signal n31_adj_594 : std_logic;
signal \n32_adj_593_cascade_\ : std_logic;
signal n2910 : std_logic;
signal n30_adj_595 : std_logic;
signal n29_adj_596 : std_logic;
signal n2801 : std_logic;
signal n313 : std_logic;
signal n2742 : std_logic;
signal \n2833_cascade_\ : std_logic;
signal n11756 : std_logic;
signal n2932 : std_logic;
signal n315 : std_logic;
signal \n2932_cascade_\ : std_logic;
signal n2933 : std_logic;
signal n2930 : std_logic;
signal n2931 : std_logic;
signal n2929 : std_logic;
signal \n2930_cascade_\ : std_logic;
signal n11662 : std_logic;
signal n13417 : std_logic;
signal n314 : std_logic;
signal n2901 : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal n2833 : std_logic;
signal n2900 : std_logic;
signal n12411 : std_logic;
signal n2832 : std_logic;
signal n2899 : std_logic;
signal n12412 : std_logic;
signal n2831 : std_logic;
signal n2898 : std_logic;
signal n12413 : std_logic;
signal n2830 : std_logic;
signal n2897 : std_logic;
signal n12414 : std_logic;
signal n2829 : std_logic;
signal n2896 : std_logic;
signal n12415 : std_logic;
signal n2828 : std_logic;
signal n2895 : std_logic;
signal n12416 : std_logic;
signal n2827 : std_logic;
signal n2894 : std_logic;
signal n12417 : std_logic;
signal n12418 : std_logic;
signal n2826 : std_logic;
signal n2893 : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal n2825 : std_logic;
signal n2892 : std_logic;
signal n12419 : std_logic;
signal n2824 : std_logic;
signal n2891 : std_logic;
signal n12420 : std_logic;
signal n2823 : std_logic;
signal n2890 : std_logic;
signal n12421 : std_logic;
signal n2822 : std_logic;
signal n2889 : std_logic;
signal n12422 : std_logic;
signal n2821 : std_logic;
signal n2888 : std_logic;
signal n12423 : std_logic;
signal n2820 : std_logic;
signal n2887 : std_logic;
signal n12424 : std_logic;
signal n2819 : std_logic;
signal n2886 : std_logic;
signal n12425 : std_logic;
signal n12426 : std_logic;
signal n2818 : std_logic;
signal n2885 : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal n2817 : std_logic;
signal n2884 : std_logic;
signal n12427 : std_logic;
signal n2816 : std_logic;
signal n2883 : std_logic;
signal n12428 : std_logic;
signal n2815 : std_logic;
signal n2882 : std_logic;
signal n12429 : std_logic;
signal n2814 : std_logic;
signal n2881 : std_logic;
signal n12430 : std_logic;
signal n2813 : std_logic;
signal n2880 : std_logic;
signal n12431 : std_logic;
signal n2812 : std_logic;
signal n2879 : std_logic;
signal n12432 : std_logic;
signal n2811 : std_logic;
signal n2878 : std_logic;
signal n12433 : std_logic;
signal n12434 : std_logic;
signal n2810 : std_logic;
signal n2877 : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal n2809 : std_logic;
signal n2876 : std_logic;
signal n12435 : std_logic;
signal n12436 : std_logic;
signal n2808 : std_logic;
signal n2875 : std_logic;
signal n2907 : std_logic;
signal n3220 : std_logic;
signal n3287 : std_logic;
signal n17_adj_705 : std_logic;
signal n3296 : std_logic;
signal \n13822_cascade_\ : std_logic;
signal n3229 : std_logic;
signal n15_adj_704 : std_logic;
signal \n13834_cascade_\ : std_logic;
signal n13842 : std_logic;
signal n3222 : std_logic;
signal n3289 : std_logic;
signal n3286 : std_logic;
signal \n27_adj_709_cascade_\ : std_logic;
signal n3219 : std_logic;
signal n13830 : std_logic;
signal n3292 : std_logic;
signal n3225 : std_logic;
signal n3237 : std_logic;
signal n21_adj_706 : std_logic;
signal n3011 : std_logic;
signal n3078 : std_logic;
signal \n3110_cascade_\ : std_logic;
signal n3209 : std_logic;
signal n3226 : std_logic;
signal n2841 : std_logic;
signal n14921 : std_logic;
signal n3009 : std_logic;
signal n3076 : std_logic;
signal \ENCODER0_B_N\ : std_logic;
signal n3015 : std_logic;
signal n3082 : std_logic;
signal n3039 : std_logic;
signal n3138 : std_logic;
signal \n3114_cascade_\ : std_logic;
signal n3213 : std_logic;
signal \n7_adj_712_cascade_\ : std_logic;
signal n8_adj_711 : std_logic;
signal \quad_counter0.direction_N_530\ : std_logic;
signal n13676 : std_logic;
signal \n10_adj_714_cascade_\ : std_logic;
signal \n16_adj_702_cascade_\ : std_logic;
signal n19_adj_701 : std_logic;
signal n24_adj_590 : std_logic;
signal duty_3 : std_logic;
signal n22_adj_588 : std_logic;
signal \n21_adj_700_cascade_\ : std_logic;
signal n22_adj_699 : std_logic;
signal duty_1 : std_logic;
signal \pwm_setpoint_23_N_171_1\ : std_logic;
signal pwm_setpoint_1 : std_logic;
signal \quad_counter0.a_prev_N_537_cascade_\ : std_logic;
signal \quad_counter0.direction_N_534_cascade_\ : std_logic;
signal \quad_counter0.a_prev_N_537\ : std_logic;
signal \quad_counter0.a_prev\ : std_logic;
signal \quad_counter0.b_new_1\ : std_logic;
signal \quad_counter0.b_new_0\ : std_logic;
signal \quad_counter0.debounce_cnt\ : std_logic;
signal \direction_N_531\ : std_logic;
signal b_prev : std_logic;
signal n1185 : std_logic;
signal \quad_counter0.a_new_0\ : std_logic;
signal a_new_1 : std_logic;
signal duty_19 : std_logic;
signal n6_adj_572 : std_logic;
signal duty_18 : std_logic;
signal n7_adj_573 : std_logic;
signal sweep_counter_0 : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal sweep_counter_1 : std_logic;
signal n12606 : std_logic;
signal sweep_counter_2 : std_logic;
signal n12607 : std_logic;
signal sweep_counter_3 : std_logic;
signal n12608 : std_logic;
signal sweep_counter_4 : std_logic;
signal n12609 : std_logic;
signal sweep_counter_5 : std_logic;
signal n12610 : std_logic;
signal sweep_counter_6 : std_logic;
signal n12611 : std_logic;
signal sweep_counter_7 : std_logic;
signal n12612 : std_logic;
signal n12613 : std_logic;
signal sweep_counter_8 : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal sweep_counter_9 : std_logic;
signal n12614 : std_logic;
signal sweep_counter_10 : std_logic;
signal n12615 : std_logic;
signal sweep_counter_11 : std_logic;
signal n12616 : std_logic;
signal sweep_counter_12 : std_logic;
signal n12617 : std_logic;
signal sweep_counter_13 : std_logic;
signal n12618 : std_logic;
signal sweep_counter_14 : std_logic;
signal n12619 : std_logic;
signal sweep_counter_15 : std_logic;
signal n12620 : std_logic;
signal n12621 : std_logic;
signal sweep_counter_16 : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal n12622 : std_logic;
signal sweep_counter_17 : std_logic;
signal n317 : std_logic;
signal n3201 : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal n3133 : std_logic;
signal n3200 : std_logic;
signal n12492 : std_logic;
signal n3132 : std_logic;
signal n3199 : std_logic;
signal n12493 : std_logic;
signal n3131 : std_logic;
signal n3198 : std_logic;
signal n12494 : std_logic;
signal n3130 : std_logic;
signal n3197 : std_logic;
signal n12495 : std_logic;
signal n3129 : std_logic;
signal n3196 : std_logic;
signal n12496 : std_logic;
signal n3128 : std_logic;
signal n3195 : std_logic;
signal n12497 : std_logic;
signal n3127 : std_logic;
signal n3194 : std_logic;
signal n12498 : std_logic;
signal n12499 : std_logic;
signal n3126 : std_logic;
signal n3193 : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal n3125 : std_logic;
signal n3192 : std_logic;
signal n12500 : std_logic;
signal n3124 : std_logic;
signal n3191 : std_logic;
signal n12501 : std_logic;
signal n3123 : std_logic;
signal n3190 : std_logic;
signal n12502 : std_logic;
signal n3122 : std_logic;
signal n3189 : std_logic;
signal n12503 : std_logic;
signal n3121 : std_logic;
signal n3188 : std_logic;
signal n12504 : std_logic;
signal n3120 : std_logic;
signal n3187 : std_logic;
signal n12505 : std_logic;
signal n3119 : std_logic;
signal n3186 : std_logic;
signal n12506 : std_logic;
signal n12507 : std_logic;
signal n3118 : std_logic;
signal n3185 : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal n3117 : std_logic;
signal n3184 : std_logic;
signal n12508 : std_logic;
signal n3116 : std_logic;
signal n3183 : std_logic;
signal n12509 : std_logic;
signal n3115 : std_logic;
signal n3182 : std_logic;
signal n12510 : std_logic;
signal n3114 : std_logic;
signal n3181 : std_logic;
signal n12511 : std_logic;
signal n3113 : std_logic;
signal n3180 : std_logic;
signal n12512 : std_logic;
signal n3112 : std_logic;
signal n3179 : std_logic;
signal n12513 : std_logic;
signal n3111 : std_logic;
signal n3178 : std_logic;
signal n12514 : std_logic;
signal n12515 : std_logic;
signal n3110 : std_logic;
signal n3177 : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal n3109 : std_logic;
signal n3176 : std_logic;
signal n12516 : std_logic;
signal n3108 : std_logic;
signal n3175 : std_logic;
signal n12517 : std_logic;
signal n3107 : std_logic;
signal n3174 : std_logic;
signal n12518 : std_logic;
signal n3106 : std_logic;
signal n3173 : std_logic;
signal n12519 : std_logic;
signal n15158 : std_logic;
signal n3105 : std_logic;
signal n12520 : std_logic;
signal n3204 : std_logic;
signal encoder0_position_target_0 : std_logic;
signal \bfn_16_26_0_\ : std_logic;
signal encoder0_position_target_1 : std_logic;
signal n12663 : std_logic;
signal encoder0_position_target_2 : std_logic;
signal n12664 : std_logic;
signal encoder0_position_target_3 : std_logic;
signal n12665 : std_logic;
signal encoder0_position_target_4 : std_logic;
signal n12666 : std_logic;
signal encoder0_position_target_5 : std_logic;
signal n12667 : std_logic;
signal encoder0_position_target_6 : std_logic;
signal n12668 : std_logic;
signal encoder0_position_target_7 : std_logic;
signal n12669 : std_logic;
signal n12670 : std_logic;
signal encoder0_position_target_8 : std_logic;
signal \bfn_16_27_0_\ : std_logic;
signal encoder0_position_target_9 : std_logic;
signal n12671 : std_logic;
signal encoder0_position_target_10 : std_logic;
signal n12672 : std_logic;
signal encoder0_position_target_11 : std_logic;
signal n12673 : std_logic;
signal encoder0_position_target_12 : std_logic;
signal n12674 : std_logic;
signal encoder0_position_target_13 : std_logic;
signal n12675 : std_logic;
signal encoder0_position_target_14 : std_logic;
signal n12676 : std_logic;
signal encoder0_position_target_15 : std_logic;
signal n12677 : std_logic;
signal n12678 : std_logic;
signal encoder0_position_target_16 : std_logic;
signal \bfn_16_28_0_\ : std_logic;
signal encoder0_position_target_17 : std_logic;
signal n12679 : std_logic;
signal encoder0_position_target_18 : std_logic;
signal n12680 : std_logic;
signal encoder0_position_target_19 : std_logic;
signal n12681 : std_logic;
signal encoder0_position_target_20 : std_logic;
signal n12682 : std_logic;
signal encoder0_position_target_21 : std_logic;
signal n12683 : std_logic;
signal encoder0_position_target_22 : std_logic;
signal n12684 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n12685 : std_logic;
signal encoder0_position_target_23 : std_logic;
signal n4856 : std_logic;
signal n4890 : std_logic;
signal \pwm_setpoint_23_N_171_9\ : std_logic;
signal duty_9 : std_logic;
signal pwm_setpoint_9 : std_logic;
signal duty_8 : std_logic;
signal n17_adj_583 : std_logic;
signal commutation_state_prev_1 : std_logic;
signal duty_23 : std_logic;
signal \pwm_setpoint_23__N_195\ : std_logic;
signal encoder0_position_scaled_6 : std_logic;
signal n19_adj_551 : std_logic;
signal dti : std_logic;
signal n4781 : std_logic;
signal \INLC_c_0\ : std_logic;
signal \INLA_c_0\ : std_logic;
signal \INLB_c_0\ : std_logic;
signal dir : std_logic;
signal commutation_state_1 : std_logic;
signal commutation_state_0 : std_logic;
signal commutation_state_2 : std_logic;
signal \CLK_N\ : std_logic;
signal n4842 : std_logic;
signal n4886 : std_logic;
signal \GHA\ : std_logic;
signal \INHA_c_0\ : std_logic;
signal \GHC\ : std_logic;
signal \INHC_c_0\ : std_logic;
signal \GHB\ : std_logic;
signal pwm_out : std_logic;
signal \INHB_c_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \ENCODER0_A_wire\ : std_logic;
signal \ENCODER0_B_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \HALL1_wire\ : std_logic;
signal \HALL2_wire\ : std_logic;
signal \HALL3_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    \ENCODER0_A_wire\ <= ENCODER0_A;
    \ENCODER0_B_wire\ <= ENCODER0_B;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \HALL1_wire\ <= HALL1;
    \HALL2_wire\ <= HALL2;
    \HALL3_wire\ <= HALL3;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56636\,
            DIN => \N__56635\,
            DOUT => \N__56634\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56636\,
            PADOUT => \N__56635\,
            PADIN => \N__56634\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56627\,
            DIN => \N__56626\,
            DOUT => \N__56625\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56627\,
            PADOUT => \N__56626\,
            PADIN => \N__56625\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56618\,
            DIN => \N__56617\,
            DOUT => \N__56616\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56618\,
            PADOUT => \N__56617\,
            PADIN => \N__56616\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ENCODER0_A_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56609\,
            DIN => \N__56608\,
            DOUT => \N__56607\,
            PACKAGEPIN => \ENCODER0_A_wire\
        );

    \ENCODER0_A_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56609\,
            PADOUT => \N__56608\,
            PADIN => \N__56607\,
            CLOCKENABLE => 'H',
            DIN0 => \ENCODER0_A_N\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ENCODER0_B_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56600\,
            DIN => \N__56599\,
            DOUT => \N__56598\,
            PACKAGEPIN => \ENCODER0_B_wire\
        );

    \ENCODER0_B_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56600\,
            PADOUT => \N__56599\,
            PADIN => \N__56598\,
            CLOCKENABLE => 'H',
            DIN0 => \ENCODER0_B_N\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56591\,
            DIN => \N__56590\,
            DOUT => \N__56589\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56591\,
            PADOUT => \N__56590\,
            PADIN => \N__56589\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55810\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56582\,
            DIN => \N__56581\,
            DOUT => \N__56580\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56582\,
            PADOUT => \N__56581\,
            PADIN => \N__56580\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55744\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56573\,
            DIN => \N__56572\,
            DOUT => \N__56571\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56573\,
            PADOUT => \N__56572\,
            PADIN => \N__56571\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55789\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56564\,
            DIN => \N__56563\,
            DOUT => \N__56562\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56564\,
            PADOUT => \N__56563\,
            PADIN => \N__56562\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55411\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56555\,
            DIN => \N__56554\,
            DOUT => \N__56553\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56555\,
            PADOUT => \N__56554\,
            PADIN => \N__56553\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__56455\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56546\,
            DIN => \N__56545\,
            DOUT => \N__56544\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56546\,
            PADOUT => \N__56545\,
            PADIN => \N__56544\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55426\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56537\,
            DIN => \N__56536\,
            DOUT => \N__56535\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56537\,
            PADOUT => \N__56536\,
            PADIN => \N__56535\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36871\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56528\,
            DIN => \N__56527\,
            DOUT => \N__56526\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56528\,
            PADOUT => \N__56527\,
            PADIN => \N__56526\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56519\,
            DIN => \N__56518\,
            DOUT => \N__56517\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56519\,
            PADOUT => \N__56518\,
            PADIN => \N__56517\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56510\,
            DIN => \N__56509\,
            DOUT => \N__56508\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56510\,
            PADOUT => \N__56509\,
            PADIN => \N__56508\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall1_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56501\,
            DIN => \N__56500\,
            DOUT => \N__56499\,
            PACKAGEPIN => \HALL1_wire\
        );

    \hall1_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56501\,
            PADOUT => \N__56500\,
            PADIN => \N__56499\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_2\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__56041\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall2_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56492\,
            DIN => \N__56491\,
            DOUT => \N__56490\,
            PACKAGEPIN => \HALL2_wire\
        );

    \hall2_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56492\,
            PADOUT => \N__56491\,
            PADIN => \N__56490\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_1\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__56039\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall3_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56483\,
            DIN => \N__56482\,
            DOUT => \N__56481\,
            PACKAGEPIN => \HALL3_wire\
        );

    \hall3_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56483\,
            PADOUT => \N__56482\,
            PADIN => \N__56481\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_0\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__56039\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56474\,
            DIN => \N__56473\,
            DOUT => \N__56472\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56474\,
            PADOUT => \N__56473\,
            PADIN => \N__56472\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__13460\ : IoInMux
    port map (
            O => \N__56455\,
            I => \N__56452\
        );

    \I__13459\ : LocalMux
    port map (
            O => \N__56452\,
            I => \N__56449\
        );

    \I__13458\ : IoSpan4Mux
    port map (
            O => \N__56449\,
            I => \N__56446\
        );

    \I__13457\ : Span4Mux_s1_v
    port map (
            O => \N__56446\,
            I => \N__56443\
        );

    \I__13456\ : Span4Mux_h
    port map (
            O => \N__56443\,
            I => \N__56440\
        );

    \I__13455\ : Odrv4
    port map (
            O => \N__56440\,
            I => \INLB_c_0\
        );

    \I__13454\ : InMux
    port map (
            O => \N__56437\,
            I => \N__56431\
        );

    \I__13453\ : InMux
    port map (
            O => \N__56436\,
            I => \N__56424\
        );

    \I__13452\ : InMux
    port map (
            O => \N__56435\,
            I => \N__56424\
        );

    \I__13451\ : CascadeMux
    port map (
            O => \N__56434\,
            I => \N__56421\
        );

    \I__13450\ : LocalMux
    port map (
            O => \N__56431\,
            I => \N__56418\
        );

    \I__13449\ : InMux
    port map (
            O => \N__56430\,
            I => \N__56413\
        );

    \I__13448\ : InMux
    port map (
            O => \N__56429\,
            I => \N__56413\
        );

    \I__13447\ : LocalMux
    port map (
            O => \N__56424\,
            I => \N__56410\
        );

    \I__13446\ : InMux
    port map (
            O => \N__56421\,
            I => \N__56407\
        );

    \I__13445\ : Span4Mux_s2_v
    port map (
            O => \N__56418\,
            I => \N__56404\
        );

    \I__13444\ : LocalMux
    port map (
            O => \N__56413\,
            I => \N__56399\
        );

    \I__13443\ : Span4Mux_s2_v
    port map (
            O => \N__56410\,
            I => \N__56399\
        );

    \I__13442\ : LocalMux
    port map (
            O => \N__56407\,
            I => dir
        );

    \I__13441\ : Odrv4
    port map (
            O => \N__56404\,
            I => dir
        );

    \I__13440\ : Odrv4
    port map (
            O => \N__56399\,
            I => dir
        );

    \I__13439\ : InMux
    port map (
            O => \N__56392\,
            I => \N__56383\
        );

    \I__13438\ : InMux
    port map (
            O => \N__56391\,
            I => \N__56383\
        );

    \I__13437\ : InMux
    port map (
            O => \N__56390\,
            I => \N__56377\
        );

    \I__13436\ : InMux
    port map (
            O => \N__56389\,
            I => \N__56377\
        );

    \I__13435\ : InMux
    port map (
            O => \N__56388\,
            I => \N__56371\
        );

    \I__13434\ : LocalMux
    port map (
            O => \N__56383\,
            I => \N__56368\
        );

    \I__13433\ : InMux
    port map (
            O => \N__56382\,
            I => \N__56365\
        );

    \I__13432\ : LocalMux
    port map (
            O => \N__56377\,
            I => \N__56362\
        );

    \I__13431\ : InMux
    port map (
            O => \N__56376\,
            I => \N__56359\
        );

    \I__13430\ : InMux
    port map (
            O => \N__56375\,
            I => \N__56354\
        );

    \I__13429\ : InMux
    port map (
            O => \N__56374\,
            I => \N__56354\
        );

    \I__13428\ : LocalMux
    port map (
            O => \N__56371\,
            I => \N__56350\
        );

    \I__13427\ : Span4Mux_v
    port map (
            O => \N__56368\,
            I => \N__56347\
        );

    \I__13426\ : LocalMux
    port map (
            O => \N__56365\,
            I => \N__56344\
        );

    \I__13425\ : Span4Mux_v
    port map (
            O => \N__56362\,
            I => \N__56341\
        );

    \I__13424\ : LocalMux
    port map (
            O => \N__56359\,
            I => \N__56336\
        );

    \I__13423\ : LocalMux
    port map (
            O => \N__56354\,
            I => \N__56336\
        );

    \I__13422\ : CascadeMux
    port map (
            O => \N__56353\,
            I => \N__56333\
        );

    \I__13421\ : Span4Mux_h
    port map (
            O => \N__56350\,
            I => \N__56330\
        );

    \I__13420\ : Span4Mux_h
    port map (
            O => \N__56347\,
            I => \N__56323\
        );

    \I__13419\ : Span4Mux_v
    port map (
            O => \N__56344\,
            I => \N__56323\
        );

    \I__13418\ : Span4Mux_h
    port map (
            O => \N__56341\,
            I => \N__56323\
        );

    \I__13417\ : Span4Mux_v
    port map (
            O => \N__56336\,
            I => \N__56320\
        );

    \I__13416\ : InMux
    port map (
            O => \N__56333\,
            I => \N__56317\
        );

    \I__13415\ : Span4Mux_v
    port map (
            O => \N__56330\,
            I => \N__56314\
        );

    \I__13414\ : Sp12to4
    port map (
            O => \N__56323\,
            I => \N__56309\
        );

    \I__13413\ : Sp12to4
    port map (
            O => \N__56320\,
            I => \N__56309\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__56317\,
            I => commutation_state_1
        );

    \I__13411\ : Odrv4
    port map (
            O => \N__56314\,
            I => commutation_state_1
        );

    \I__13410\ : Odrv12
    port map (
            O => \N__56309\,
            I => commutation_state_1
        );

    \I__13409\ : CascadeMux
    port map (
            O => \N__56302\,
            I => \N__56297\
        );

    \I__13408\ : InMux
    port map (
            O => \N__56301\,
            I => \N__56291\
        );

    \I__13407\ : InMux
    port map (
            O => \N__56300\,
            I => \N__56286\
        );

    \I__13406\ : InMux
    port map (
            O => \N__56297\,
            I => \N__56286\
        );

    \I__13405\ : InMux
    port map (
            O => \N__56296\,
            I => \N__56283\
        );

    \I__13404\ : InMux
    port map (
            O => \N__56295\,
            I => \N__56278\
        );

    \I__13403\ : InMux
    port map (
            O => \N__56294\,
            I => \N__56278\
        );

    \I__13402\ : LocalMux
    port map (
            O => \N__56291\,
            I => \N__56272\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__56286\,
            I => \N__56265\
        );

    \I__13400\ : LocalMux
    port map (
            O => \N__56283\,
            I => \N__56265\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__56278\,
            I => \N__56265\
        );

    \I__13398\ : InMux
    port map (
            O => \N__56277\,
            I => \N__56260\
        );

    \I__13397\ : InMux
    port map (
            O => \N__56276\,
            I => \N__56260\
        );

    \I__13396\ : InMux
    port map (
            O => \N__56275\,
            I => \N__56257\
        );

    \I__13395\ : Sp12to4
    port map (
            O => \N__56272\,
            I => \N__56247\
        );

    \I__13394\ : Span4Mux_s3_v
    port map (
            O => \N__56265\,
            I => \N__56244\
        );

    \I__13393\ : LocalMux
    port map (
            O => \N__56260\,
            I => \N__56241\
        );

    \I__13392\ : LocalMux
    port map (
            O => \N__56257\,
            I => \N__56238\
        );

    \I__13391\ : InMux
    port map (
            O => \N__56256\,
            I => \N__56227\
        );

    \I__13390\ : InMux
    port map (
            O => \N__56255\,
            I => \N__56227\
        );

    \I__13389\ : InMux
    port map (
            O => \N__56254\,
            I => \N__56227\
        );

    \I__13388\ : InMux
    port map (
            O => \N__56253\,
            I => \N__56227\
        );

    \I__13387\ : InMux
    port map (
            O => \N__56252\,
            I => \N__56227\
        );

    \I__13386\ : InMux
    port map (
            O => \N__56251\,
            I => \N__56224\
        );

    \I__13385\ : InMux
    port map (
            O => \N__56250\,
            I => \N__56221\
        );

    \I__13384\ : Span12Mux_s3_v
    port map (
            O => \N__56247\,
            I => \N__56216\
        );

    \I__13383\ : Sp12to4
    port map (
            O => \N__56244\,
            I => \N__56216\
        );

    \I__13382\ : Span4Mux_v
    port map (
            O => \N__56241\,
            I => \N__56211\
        );

    \I__13381\ : Span4Mux_v
    port map (
            O => \N__56238\,
            I => \N__56211\
        );

    \I__13380\ : LocalMux
    port map (
            O => \N__56227\,
            I => \N__56206\
        );

    \I__13379\ : LocalMux
    port map (
            O => \N__56224\,
            I => \N__56206\
        );

    \I__13378\ : LocalMux
    port map (
            O => \N__56221\,
            I => commutation_state_0
        );

    \I__13377\ : Odrv12
    port map (
            O => \N__56216\,
            I => commutation_state_0
        );

    \I__13376\ : Odrv4
    port map (
            O => \N__56211\,
            I => commutation_state_0
        );

    \I__13375\ : Odrv4
    port map (
            O => \N__56206\,
            I => commutation_state_0
        );

    \I__13374\ : CascadeMux
    port map (
            O => \N__56197\,
            I => \N__56191\
        );

    \I__13373\ : CascadeMux
    port map (
            O => \N__56196\,
            I => \N__56188\
        );

    \I__13372\ : CascadeMux
    port map (
            O => \N__56195\,
            I => \N__56184\
        );

    \I__13371\ : CascadeMux
    port map (
            O => \N__56194\,
            I => \N__56181\
        );

    \I__13370\ : InMux
    port map (
            O => \N__56191\,
            I => \N__56175\
        );

    \I__13369\ : InMux
    port map (
            O => \N__56188\,
            I => \N__56175\
        );

    \I__13368\ : InMux
    port map (
            O => \N__56187\,
            I => \N__56169\
        );

    \I__13367\ : InMux
    port map (
            O => \N__56184\,
            I => \N__56169\
        );

    \I__13366\ : InMux
    port map (
            O => \N__56181\,
            I => \N__56166\
        );

    \I__13365\ : CascadeMux
    port map (
            O => \N__56180\,
            I => \N__56162\
        );

    \I__13364\ : LocalMux
    port map (
            O => \N__56175\,
            I => \N__56159\
        );

    \I__13363\ : CascadeMux
    port map (
            O => \N__56174\,
            I => \N__56156\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__56169\,
            I => \N__56151\
        );

    \I__13361\ : LocalMux
    port map (
            O => \N__56166\,
            I => \N__56151\
        );

    \I__13360\ : InMux
    port map (
            O => \N__56165\,
            I => \N__56146\
        );

    \I__13359\ : InMux
    port map (
            O => \N__56162\,
            I => \N__56146\
        );

    \I__13358\ : Span4Mux_h
    port map (
            O => \N__56159\,
            I => \N__56142\
        );

    \I__13357\ : InMux
    port map (
            O => \N__56156\,
            I => \N__56139\
        );

    \I__13356\ : Span4Mux_h
    port map (
            O => \N__56151\,
            I => \N__56134\
        );

    \I__13355\ : LocalMux
    port map (
            O => \N__56146\,
            I => \N__56134\
        );

    \I__13354\ : InMux
    port map (
            O => \N__56145\,
            I => \N__56130\
        );

    \I__13353\ : Span4Mux_h
    port map (
            O => \N__56142\,
            I => \N__56127\
        );

    \I__13352\ : LocalMux
    port map (
            O => \N__56139\,
            I => \N__56124\
        );

    \I__13351\ : Span4Mux_h
    port map (
            O => \N__56134\,
            I => \N__56121\
        );

    \I__13350\ : InMux
    port map (
            O => \N__56133\,
            I => \N__56118\
        );

    \I__13349\ : LocalMux
    port map (
            O => \N__56130\,
            I => \N__56115\
        );

    \I__13348\ : Span4Mux_h
    port map (
            O => \N__56127\,
            I => \N__56112\
        );

    \I__13347\ : Span4Mux_h
    port map (
            O => \N__56124\,
            I => \N__56107\
        );

    \I__13346\ : Span4Mux_h
    port map (
            O => \N__56121\,
            I => \N__56107\
        );

    \I__13345\ : LocalMux
    port map (
            O => \N__56118\,
            I => commutation_state_2
        );

    \I__13344\ : Odrv4
    port map (
            O => \N__56115\,
            I => commutation_state_2
        );

    \I__13343\ : Odrv4
    port map (
            O => \N__56112\,
            I => commutation_state_2
        );

    \I__13342\ : Odrv4
    port map (
            O => \N__56107\,
            I => commutation_state_2
        );

    \I__13341\ : ClkMux
    port map (
            O => \N__56098\,
            I => \N__55918\
        );

    \I__13340\ : ClkMux
    port map (
            O => \N__56097\,
            I => \N__55918\
        );

    \I__13339\ : ClkMux
    port map (
            O => \N__56096\,
            I => \N__55918\
        );

    \I__13338\ : ClkMux
    port map (
            O => \N__56095\,
            I => \N__55918\
        );

    \I__13337\ : ClkMux
    port map (
            O => \N__56094\,
            I => \N__55918\
        );

    \I__13336\ : ClkMux
    port map (
            O => \N__56093\,
            I => \N__55918\
        );

    \I__13335\ : ClkMux
    port map (
            O => \N__56092\,
            I => \N__55918\
        );

    \I__13334\ : ClkMux
    port map (
            O => \N__56091\,
            I => \N__55918\
        );

    \I__13333\ : ClkMux
    port map (
            O => \N__56090\,
            I => \N__55918\
        );

    \I__13332\ : ClkMux
    port map (
            O => \N__56089\,
            I => \N__55918\
        );

    \I__13331\ : ClkMux
    port map (
            O => \N__56088\,
            I => \N__55918\
        );

    \I__13330\ : ClkMux
    port map (
            O => \N__56087\,
            I => \N__55918\
        );

    \I__13329\ : ClkMux
    port map (
            O => \N__56086\,
            I => \N__55918\
        );

    \I__13328\ : ClkMux
    port map (
            O => \N__56085\,
            I => \N__55918\
        );

    \I__13327\ : ClkMux
    port map (
            O => \N__56084\,
            I => \N__55918\
        );

    \I__13326\ : ClkMux
    port map (
            O => \N__56083\,
            I => \N__55918\
        );

    \I__13325\ : ClkMux
    port map (
            O => \N__56082\,
            I => \N__55918\
        );

    \I__13324\ : ClkMux
    port map (
            O => \N__56081\,
            I => \N__55918\
        );

    \I__13323\ : ClkMux
    port map (
            O => \N__56080\,
            I => \N__55918\
        );

    \I__13322\ : ClkMux
    port map (
            O => \N__56079\,
            I => \N__55918\
        );

    \I__13321\ : ClkMux
    port map (
            O => \N__56078\,
            I => \N__55918\
        );

    \I__13320\ : ClkMux
    port map (
            O => \N__56077\,
            I => \N__55918\
        );

    \I__13319\ : ClkMux
    port map (
            O => \N__56076\,
            I => \N__55918\
        );

    \I__13318\ : ClkMux
    port map (
            O => \N__56075\,
            I => \N__55918\
        );

    \I__13317\ : ClkMux
    port map (
            O => \N__56074\,
            I => \N__55918\
        );

    \I__13316\ : ClkMux
    port map (
            O => \N__56073\,
            I => \N__55918\
        );

    \I__13315\ : ClkMux
    port map (
            O => \N__56072\,
            I => \N__55918\
        );

    \I__13314\ : ClkMux
    port map (
            O => \N__56071\,
            I => \N__55918\
        );

    \I__13313\ : ClkMux
    port map (
            O => \N__56070\,
            I => \N__55918\
        );

    \I__13312\ : ClkMux
    port map (
            O => \N__56069\,
            I => \N__55918\
        );

    \I__13311\ : ClkMux
    port map (
            O => \N__56068\,
            I => \N__55918\
        );

    \I__13310\ : ClkMux
    port map (
            O => \N__56067\,
            I => \N__55918\
        );

    \I__13309\ : ClkMux
    port map (
            O => \N__56066\,
            I => \N__55918\
        );

    \I__13308\ : ClkMux
    port map (
            O => \N__56065\,
            I => \N__55918\
        );

    \I__13307\ : ClkMux
    port map (
            O => \N__56064\,
            I => \N__55918\
        );

    \I__13306\ : ClkMux
    port map (
            O => \N__56063\,
            I => \N__55918\
        );

    \I__13305\ : ClkMux
    port map (
            O => \N__56062\,
            I => \N__55918\
        );

    \I__13304\ : ClkMux
    port map (
            O => \N__56061\,
            I => \N__55918\
        );

    \I__13303\ : ClkMux
    port map (
            O => \N__56060\,
            I => \N__55918\
        );

    \I__13302\ : ClkMux
    port map (
            O => \N__56059\,
            I => \N__55918\
        );

    \I__13301\ : ClkMux
    port map (
            O => \N__56058\,
            I => \N__55918\
        );

    \I__13300\ : ClkMux
    port map (
            O => \N__56057\,
            I => \N__55918\
        );

    \I__13299\ : ClkMux
    port map (
            O => \N__56056\,
            I => \N__55918\
        );

    \I__13298\ : ClkMux
    port map (
            O => \N__56055\,
            I => \N__55918\
        );

    \I__13297\ : ClkMux
    port map (
            O => \N__56054\,
            I => \N__55918\
        );

    \I__13296\ : ClkMux
    port map (
            O => \N__56053\,
            I => \N__55918\
        );

    \I__13295\ : ClkMux
    port map (
            O => \N__56052\,
            I => \N__55918\
        );

    \I__13294\ : ClkMux
    port map (
            O => \N__56051\,
            I => \N__55918\
        );

    \I__13293\ : ClkMux
    port map (
            O => \N__56050\,
            I => \N__55918\
        );

    \I__13292\ : ClkMux
    port map (
            O => \N__56049\,
            I => \N__55918\
        );

    \I__13291\ : ClkMux
    port map (
            O => \N__56048\,
            I => \N__55918\
        );

    \I__13290\ : ClkMux
    port map (
            O => \N__56047\,
            I => \N__55918\
        );

    \I__13289\ : ClkMux
    port map (
            O => \N__56046\,
            I => \N__55918\
        );

    \I__13288\ : ClkMux
    port map (
            O => \N__56045\,
            I => \N__55918\
        );

    \I__13287\ : ClkMux
    port map (
            O => \N__56044\,
            I => \N__55918\
        );

    \I__13286\ : ClkMux
    port map (
            O => \N__56043\,
            I => \N__55918\
        );

    \I__13285\ : ClkMux
    port map (
            O => \N__56042\,
            I => \N__55918\
        );

    \I__13284\ : ClkMux
    port map (
            O => \N__56041\,
            I => \N__55918\
        );

    \I__13283\ : ClkMux
    port map (
            O => \N__56040\,
            I => \N__55918\
        );

    \I__13282\ : ClkMux
    port map (
            O => \N__56039\,
            I => \N__55918\
        );

    \I__13281\ : GlobalMux
    port map (
            O => \N__55918\,
            I => \N__55915\
        );

    \I__13280\ : gio2CtrlBuf
    port map (
            O => \N__55915\,
            I => \CLK_N\
        );

    \I__13279\ : CEMux
    port map (
            O => \N__55912\,
            I => \N__55909\
        );

    \I__13278\ : LocalMux
    port map (
            O => \N__55909\,
            I => \N__55905\
        );

    \I__13277\ : CEMux
    port map (
            O => \N__55908\,
            I => \N__55902\
        );

    \I__13276\ : Span4Mux_v
    port map (
            O => \N__55905\,
            I => \N__55897\
        );

    \I__13275\ : LocalMux
    port map (
            O => \N__55902\,
            I => \N__55894\
        );

    \I__13274\ : CEMux
    port map (
            O => \N__55901\,
            I => \N__55891\
        );

    \I__13273\ : CEMux
    port map (
            O => \N__55900\,
            I => \N__55888\
        );

    \I__13272\ : Span4Mux_s1_v
    port map (
            O => \N__55897\,
            I => \N__55884\
        );

    \I__13271\ : Sp12to4
    port map (
            O => \N__55894\,
            I => \N__55879\
        );

    \I__13270\ : LocalMux
    port map (
            O => \N__55891\,
            I => \N__55879\
        );

    \I__13269\ : LocalMux
    port map (
            O => \N__55888\,
            I => \N__55876\
        );

    \I__13268\ : InMux
    port map (
            O => \N__55887\,
            I => \N__55873\
        );

    \I__13267\ : Odrv4
    port map (
            O => \N__55884\,
            I => n4842
        );

    \I__13266\ : Odrv12
    port map (
            O => \N__55879\,
            I => n4842
        );

    \I__13265\ : Odrv4
    port map (
            O => \N__55876\,
            I => n4842
        );

    \I__13264\ : LocalMux
    port map (
            O => \N__55873\,
            I => n4842
        );

    \I__13263\ : SRMux
    port map (
            O => \N__55864\,
            I => \N__55861\
        );

    \I__13262\ : LocalMux
    port map (
            O => \N__55861\,
            I => \N__55856\
        );

    \I__13261\ : SRMux
    port map (
            O => \N__55860\,
            I => \N__55852\
        );

    \I__13260\ : SRMux
    port map (
            O => \N__55859\,
            I => \N__55849\
        );

    \I__13259\ : Span4Mux_h
    port map (
            O => \N__55856\,
            I => \N__55846\
        );

    \I__13258\ : SRMux
    port map (
            O => \N__55855\,
            I => \N__55843\
        );

    \I__13257\ : LocalMux
    port map (
            O => \N__55852\,
            I => \N__55840\
        );

    \I__13256\ : LocalMux
    port map (
            O => \N__55849\,
            I => \N__55837\
        );

    \I__13255\ : Span4Mux_h
    port map (
            O => \N__55846\,
            I => \N__55832\
        );

    \I__13254\ : LocalMux
    port map (
            O => \N__55843\,
            I => \N__55832\
        );

    \I__13253\ : Span4Mux_h
    port map (
            O => \N__55840\,
            I => \N__55829\
        );

    \I__13252\ : Span4Mux_h
    port map (
            O => \N__55837\,
            I => \N__55826\
        );

    \I__13251\ : Span4Mux_s2_v
    port map (
            O => \N__55832\,
            I => \N__55823\
        );

    \I__13250\ : Odrv4
    port map (
            O => \N__55829\,
            I => n4886
        );

    \I__13249\ : Odrv4
    port map (
            O => \N__55826\,
            I => n4886
        );

    \I__13248\ : Odrv4
    port map (
            O => \N__55823\,
            I => n4886
        );

    \I__13247\ : InMux
    port map (
            O => \N__55816\,
            I => \N__55813\
        );

    \I__13246\ : LocalMux
    port map (
            O => \N__55813\,
            I => \GHA\
        );

    \I__13245\ : IoInMux
    port map (
            O => \N__55810\,
            I => \N__55807\
        );

    \I__13244\ : LocalMux
    port map (
            O => \N__55807\,
            I => \N__55804\
        );

    \I__13243\ : IoSpan4Mux
    port map (
            O => \N__55804\,
            I => \N__55801\
        );

    \I__13242\ : Span4Mux_s0_v
    port map (
            O => \N__55801\,
            I => \N__55798\
        );

    \I__13241\ : Odrv4
    port map (
            O => \N__55798\,
            I => \INHA_c_0\
        );

    \I__13240\ : InMux
    port map (
            O => \N__55795\,
            I => \N__55792\
        );

    \I__13239\ : LocalMux
    port map (
            O => \N__55792\,
            I => \GHC\
        );

    \I__13238\ : IoInMux
    port map (
            O => \N__55789\,
            I => \N__55786\
        );

    \I__13237\ : LocalMux
    port map (
            O => \N__55786\,
            I => \N__55783\
        );

    \I__13236\ : Span12Mux_s2_v
    port map (
            O => \N__55783\,
            I => \N__55780\
        );

    \I__13235\ : Odrv12
    port map (
            O => \N__55780\,
            I => \INHC_c_0\
        );

    \I__13234\ : InMux
    port map (
            O => \N__55777\,
            I => \N__55774\
        );

    \I__13233\ : LocalMux
    port map (
            O => \N__55774\,
            I => \GHB\
        );

    \I__13232\ : InMux
    port map (
            O => \N__55771\,
            I => \N__55768\
        );

    \I__13231\ : LocalMux
    port map (
            O => \N__55768\,
            I => \N__55763\
        );

    \I__13230\ : InMux
    port map (
            O => \N__55767\,
            I => \N__55758\
        );

    \I__13229\ : InMux
    port map (
            O => \N__55766\,
            I => \N__55758\
        );

    \I__13228\ : Span4Mux_s2_v
    port map (
            O => \N__55763\,
            I => \N__55755\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__55758\,
            I => \N__55752\
        );

    \I__13226\ : Sp12to4
    port map (
            O => \N__55755\,
            I => \N__55747\
        );

    \I__13225\ : Sp12to4
    port map (
            O => \N__55752\,
            I => \N__55747\
        );

    \I__13224\ : Odrv12
    port map (
            O => \N__55747\,
            I => pwm_out
        );

    \I__13223\ : IoInMux
    port map (
            O => \N__55744\,
            I => \N__55741\
        );

    \I__13222\ : LocalMux
    port map (
            O => \N__55741\,
            I => \N__55738\
        );

    \I__13221\ : Span4Mux_s2_v
    port map (
            O => \N__55738\,
            I => \N__55735\
        );

    \I__13220\ : Span4Mux_h
    port map (
            O => \N__55735\,
            I => \N__55732\
        );

    \I__13219\ : Odrv4
    port map (
            O => \N__55732\,
            I => \INHB_c_0\
        );

    \I__13218\ : InMux
    port map (
            O => \N__55729\,
            I => \N__55726\
        );

    \I__13217\ : LocalMux
    port map (
            O => \N__55726\,
            I => \N__55723\
        );

    \I__13216\ : Span4Mux_h
    port map (
            O => \N__55723\,
            I => \N__55720\
        );

    \I__13215\ : Span4Mux_h
    port map (
            O => \N__55720\,
            I => \N__55717\
        );

    \I__13214\ : Odrv4
    port map (
            O => \N__55717\,
            I => commutation_state_prev_1
        );

    \I__13213\ : CascadeMux
    port map (
            O => \N__55714\,
            I => \N__55703\
        );

    \I__13212\ : InMux
    port map (
            O => \N__55713\,
            I => \N__55685\
        );

    \I__13211\ : InMux
    port map (
            O => \N__55712\,
            I => \N__55685\
        );

    \I__13210\ : InMux
    port map (
            O => \N__55711\,
            I => \N__55685\
        );

    \I__13209\ : InMux
    port map (
            O => \N__55710\,
            I => \N__55685\
        );

    \I__13208\ : InMux
    port map (
            O => \N__55709\,
            I => \N__55682\
        );

    \I__13207\ : InMux
    port map (
            O => \N__55708\,
            I => \N__55679\
        );

    \I__13206\ : InMux
    port map (
            O => \N__55707\,
            I => \N__55676\
        );

    \I__13205\ : InMux
    port map (
            O => \N__55706\,
            I => \N__55673\
        );

    \I__13204\ : InMux
    port map (
            O => \N__55703\,
            I => \N__55668\
        );

    \I__13203\ : InMux
    port map (
            O => \N__55702\,
            I => \N__55668\
        );

    \I__13202\ : InMux
    port map (
            O => \N__55701\,
            I => \N__55657\
        );

    \I__13201\ : InMux
    port map (
            O => \N__55700\,
            I => \N__55657\
        );

    \I__13200\ : InMux
    port map (
            O => \N__55699\,
            I => \N__55657\
        );

    \I__13199\ : InMux
    port map (
            O => \N__55698\,
            I => \N__55657\
        );

    \I__13198\ : InMux
    port map (
            O => \N__55697\,
            I => \N__55657\
        );

    \I__13197\ : InMux
    port map (
            O => \N__55696\,
            I => \N__55648\
        );

    \I__13196\ : InMux
    port map (
            O => \N__55695\,
            I => \N__55645\
        );

    \I__13195\ : InMux
    port map (
            O => \N__55694\,
            I => \N__55641\
        );

    \I__13194\ : LocalMux
    port map (
            O => \N__55685\,
            I => \N__55638\
        );

    \I__13193\ : LocalMux
    port map (
            O => \N__55682\,
            I => \N__55633\
        );

    \I__13192\ : LocalMux
    port map (
            O => \N__55679\,
            I => \N__55633\
        );

    \I__13191\ : LocalMux
    port map (
            O => \N__55676\,
            I => \N__55628\
        );

    \I__13190\ : LocalMux
    port map (
            O => \N__55673\,
            I => \N__55628\
        );

    \I__13189\ : LocalMux
    port map (
            O => \N__55668\,
            I => \N__55623\
        );

    \I__13188\ : LocalMux
    port map (
            O => \N__55657\,
            I => \N__55623\
        );

    \I__13187\ : InMux
    port map (
            O => \N__55656\,
            I => \N__55618\
        );

    \I__13186\ : InMux
    port map (
            O => \N__55655\,
            I => \N__55618\
        );

    \I__13185\ : InMux
    port map (
            O => \N__55654\,
            I => \N__55615\
        );

    \I__13184\ : InMux
    port map (
            O => \N__55653\,
            I => \N__55608\
        );

    \I__13183\ : InMux
    port map (
            O => \N__55652\,
            I => \N__55608\
        );

    \I__13182\ : InMux
    port map (
            O => \N__55651\,
            I => \N__55608\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__55648\,
            I => \N__55605\
        );

    \I__13180\ : LocalMux
    port map (
            O => \N__55645\,
            I => \N__55602\
        );

    \I__13179\ : InMux
    port map (
            O => \N__55644\,
            I => \N__55599\
        );

    \I__13178\ : LocalMux
    port map (
            O => \N__55641\,
            I => \N__55596\
        );

    \I__13177\ : Span4Mux_h
    port map (
            O => \N__55638\,
            I => \N__55587\
        );

    \I__13176\ : Span4Mux_v
    port map (
            O => \N__55633\,
            I => \N__55587\
        );

    \I__13175\ : Span4Mux_v
    port map (
            O => \N__55628\,
            I => \N__55587\
        );

    \I__13174\ : Span4Mux_v
    port map (
            O => \N__55623\,
            I => \N__55587\
        );

    \I__13173\ : LocalMux
    port map (
            O => \N__55618\,
            I => \N__55576\
        );

    \I__13172\ : LocalMux
    port map (
            O => \N__55615\,
            I => \N__55576\
        );

    \I__13171\ : LocalMux
    port map (
            O => \N__55608\,
            I => \N__55576\
        );

    \I__13170\ : Span4Mux_h
    port map (
            O => \N__55605\,
            I => \N__55576\
        );

    \I__13169\ : Span4Mux_h
    port map (
            O => \N__55602\,
            I => \N__55576\
        );

    \I__13168\ : LocalMux
    port map (
            O => \N__55599\,
            I => duty_23
        );

    \I__13167\ : Odrv12
    port map (
            O => \N__55596\,
            I => duty_23
        );

    \I__13166\ : Odrv4
    port map (
            O => \N__55587\,
            I => duty_23
        );

    \I__13165\ : Odrv4
    port map (
            O => \N__55576\,
            I => duty_23
        );

    \I__13164\ : SRMux
    port map (
            O => \N__55567\,
            I => \N__55564\
        );

    \I__13163\ : LocalMux
    port map (
            O => \N__55564\,
            I => \N__55560\
        );

    \I__13162\ : InMux
    port map (
            O => \N__55563\,
            I => \N__55557\
        );

    \I__13161\ : Sp12to4
    port map (
            O => \N__55560\,
            I => \N__55552\
        );

    \I__13160\ : LocalMux
    port map (
            O => \N__55557\,
            I => \N__55552\
        );

    \I__13159\ : Span12Mux_s5_v
    port map (
            O => \N__55552\,
            I => \N__55549\
        );

    \I__13158\ : Odrv12
    port map (
            O => \N__55549\,
            I => \pwm_setpoint_23__N_195\
        );

    \I__13157\ : InMux
    port map (
            O => \N__55546\,
            I => \N__55543\
        );

    \I__13156\ : LocalMux
    port map (
            O => \N__55543\,
            I => \N__55540\
        );

    \I__13155\ : Span4Mux_v
    port map (
            O => \N__55540\,
            I => \N__55537\
        );

    \I__13154\ : Sp12to4
    port map (
            O => \N__55537\,
            I => \N__55534\
        );

    \I__13153\ : Odrv12
    port map (
            O => \N__55534\,
            I => encoder0_position_scaled_6
        );

    \I__13152\ : CascadeMux
    port map (
            O => \N__55531\,
            I => \N__55528\
        );

    \I__13151\ : InMux
    port map (
            O => \N__55528\,
            I => \N__55525\
        );

    \I__13150\ : LocalMux
    port map (
            O => \N__55525\,
            I => \N__55522\
        );

    \I__13149\ : Span4Mux_v
    port map (
            O => \N__55522\,
            I => \N__55519\
        );

    \I__13148\ : Odrv4
    port map (
            O => \N__55519\,
            I => n19_adj_551
        );

    \I__13147\ : InMux
    port map (
            O => \N__55516\,
            I => \N__55512\
        );

    \I__13146\ : InMux
    port map (
            O => \N__55515\,
            I => \N__55509\
        );

    \I__13145\ : LocalMux
    port map (
            O => \N__55512\,
            I => \N__55501\
        );

    \I__13144\ : LocalMux
    port map (
            O => \N__55509\,
            I => \N__55501\
        );

    \I__13143\ : InMux
    port map (
            O => \N__55508\,
            I => \N__55496\
        );

    \I__13142\ : InMux
    port map (
            O => \N__55507\,
            I => \N__55496\
        );

    \I__13141\ : InMux
    port map (
            O => \N__55506\,
            I => \N__55492\
        );

    \I__13140\ : Span4Mux_v
    port map (
            O => \N__55501\,
            I => \N__55489\
        );

    \I__13139\ : LocalMux
    port map (
            O => \N__55496\,
            I => \N__55486\
        );

    \I__13138\ : InMux
    port map (
            O => \N__55495\,
            I => \N__55483\
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__55492\,
            I => \N__55476\
        );

    \I__13136\ : Span4Mux_h
    port map (
            O => \N__55489\,
            I => \N__55476\
        );

    \I__13135\ : Span4Mux_v
    port map (
            O => \N__55486\,
            I => \N__55476\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__55483\,
            I => dti
        );

    \I__13133\ : Odrv4
    port map (
            O => \N__55476\,
            I => dti
        );

    \I__13132\ : InMux
    port map (
            O => \N__55471\,
            I => \N__55466\
        );

    \I__13131\ : InMux
    port map (
            O => \N__55470\,
            I => \N__55463\
        );

    \I__13130\ : InMux
    port map (
            O => \N__55469\,
            I => \N__55460\
        );

    \I__13129\ : LocalMux
    port map (
            O => \N__55466\,
            I => \N__55457\
        );

    \I__13128\ : LocalMux
    port map (
            O => \N__55463\,
            I => \N__55454\
        );

    \I__13127\ : LocalMux
    port map (
            O => \N__55460\,
            I => \N__55451\
        );

    \I__13126\ : Span4Mux_s3_v
    port map (
            O => \N__55457\,
            I => \N__55448\
        );

    \I__13125\ : Span4Mux_h
    port map (
            O => \N__55454\,
            I => \N__55444\
        );

    \I__13124\ : Span4Mux_h
    port map (
            O => \N__55451\,
            I => \N__55441\
        );

    \I__13123\ : Span4Mux_h
    port map (
            O => \N__55448\,
            I => \N__55438\
        );

    \I__13122\ : InMux
    port map (
            O => \N__55447\,
            I => \N__55435\
        );

    \I__13121\ : Odrv4
    port map (
            O => \N__55444\,
            I => n4781
        );

    \I__13120\ : Odrv4
    port map (
            O => \N__55441\,
            I => n4781
        );

    \I__13119\ : Odrv4
    port map (
            O => \N__55438\,
            I => n4781
        );

    \I__13118\ : LocalMux
    port map (
            O => \N__55435\,
            I => n4781
        );

    \I__13117\ : IoInMux
    port map (
            O => \N__55426\,
            I => \N__55423\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__55423\,
            I => \N__55420\
        );

    \I__13115\ : Span12Mux_s1_v
    port map (
            O => \N__55420\,
            I => \N__55417\
        );

    \I__13114\ : Span12Mux_h
    port map (
            O => \N__55417\,
            I => \N__55414\
        );

    \I__13113\ : Odrv12
    port map (
            O => \N__55414\,
            I => \INLC_c_0\
        );

    \I__13112\ : IoInMux
    port map (
            O => \N__55411\,
            I => \N__55408\
        );

    \I__13111\ : LocalMux
    port map (
            O => \N__55408\,
            I => \N__55405\
        );

    \I__13110\ : Span4Mux_s1_v
    port map (
            O => \N__55405\,
            I => \N__55402\
        );

    \I__13109\ : Span4Mux_h
    port map (
            O => \N__55402\,
            I => \N__55399\
        );

    \I__13108\ : Odrv4
    port map (
            O => \N__55399\,
            I => \INLA_c_0\
        );

    \I__13107\ : CascadeMux
    port map (
            O => \N__55396\,
            I => \N__55393\
        );

    \I__13106\ : InMux
    port map (
            O => \N__55393\,
            I => \N__55389\
        );

    \I__13105\ : InMux
    port map (
            O => \N__55392\,
            I => \N__55386\
        );

    \I__13104\ : LocalMux
    port map (
            O => \N__55389\,
            I => \N__55383\
        );

    \I__13103\ : LocalMux
    port map (
            O => \N__55386\,
            I => \N__55377\
        );

    \I__13102\ : Span4Mux_h
    port map (
            O => \N__55383\,
            I => \N__55377\
        );

    \I__13101\ : InMux
    port map (
            O => \N__55382\,
            I => \N__55374\
        );

    \I__13100\ : Odrv4
    port map (
            O => \N__55377\,
            I => encoder0_position_target_18
        );

    \I__13099\ : LocalMux
    port map (
            O => \N__55374\,
            I => encoder0_position_target_18
        );

    \I__13098\ : InMux
    port map (
            O => \N__55369\,
            I => n12680
        );

    \I__13097\ : CascadeMux
    port map (
            O => \N__55366\,
            I => \N__55363\
        );

    \I__13096\ : InMux
    port map (
            O => \N__55363\,
            I => \N__55359\
        );

    \I__13095\ : CascadeMux
    port map (
            O => \N__55362\,
            I => \N__55356\
        );

    \I__13094\ : LocalMux
    port map (
            O => \N__55359\,
            I => \N__55353\
        );

    \I__13093\ : InMux
    port map (
            O => \N__55356\,
            I => \N__55349\
        );

    \I__13092\ : Span4Mux_h
    port map (
            O => \N__55353\,
            I => \N__55346\
        );

    \I__13091\ : InMux
    port map (
            O => \N__55352\,
            I => \N__55343\
        );

    \I__13090\ : LocalMux
    port map (
            O => \N__55349\,
            I => encoder0_position_target_19
        );

    \I__13089\ : Odrv4
    port map (
            O => \N__55346\,
            I => encoder0_position_target_19
        );

    \I__13088\ : LocalMux
    port map (
            O => \N__55343\,
            I => encoder0_position_target_19
        );

    \I__13087\ : InMux
    port map (
            O => \N__55336\,
            I => n12681
        );

    \I__13086\ : CascadeMux
    port map (
            O => \N__55333\,
            I => \N__55330\
        );

    \I__13085\ : InMux
    port map (
            O => \N__55330\,
            I => \N__55326\
        );

    \I__13084\ : InMux
    port map (
            O => \N__55329\,
            I => \N__55322\
        );

    \I__13083\ : LocalMux
    port map (
            O => \N__55326\,
            I => \N__55319\
        );

    \I__13082\ : InMux
    port map (
            O => \N__55325\,
            I => \N__55316\
        );

    \I__13081\ : LocalMux
    port map (
            O => \N__55322\,
            I => encoder0_position_target_20
        );

    \I__13080\ : Odrv4
    port map (
            O => \N__55319\,
            I => encoder0_position_target_20
        );

    \I__13079\ : LocalMux
    port map (
            O => \N__55316\,
            I => encoder0_position_target_20
        );

    \I__13078\ : InMux
    port map (
            O => \N__55309\,
            I => n12682
        );

    \I__13077\ : CascadeMux
    port map (
            O => \N__55306\,
            I => \N__55302\
        );

    \I__13076\ : CascadeMux
    port map (
            O => \N__55305\,
            I => \N__55299\
        );

    \I__13075\ : InMux
    port map (
            O => \N__55302\,
            I => \N__55296\
        );

    \I__13074\ : InMux
    port map (
            O => \N__55299\,
            I => \N__55292\
        );

    \I__13073\ : LocalMux
    port map (
            O => \N__55296\,
            I => \N__55289\
        );

    \I__13072\ : InMux
    port map (
            O => \N__55295\,
            I => \N__55286\
        );

    \I__13071\ : LocalMux
    port map (
            O => \N__55292\,
            I => encoder0_position_target_21
        );

    \I__13070\ : Odrv4
    port map (
            O => \N__55289\,
            I => encoder0_position_target_21
        );

    \I__13069\ : LocalMux
    port map (
            O => \N__55286\,
            I => encoder0_position_target_21
        );

    \I__13068\ : InMux
    port map (
            O => \N__55279\,
            I => n12683
        );

    \I__13067\ : CascadeMux
    port map (
            O => \N__55276\,
            I => \N__55273\
        );

    \I__13066\ : InMux
    port map (
            O => \N__55273\,
            I => \N__55269\
        );

    \I__13065\ : InMux
    port map (
            O => \N__55272\,
            I => \N__55265\
        );

    \I__13064\ : LocalMux
    port map (
            O => \N__55269\,
            I => \N__55262\
        );

    \I__13063\ : InMux
    port map (
            O => \N__55268\,
            I => \N__55259\
        );

    \I__13062\ : LocalMux
    port map (
            O => \N__55265\,
            I => encoder0_position_target_22
        );

    \I__13061\ : Odrv4
    port map (
            O => \N__55262\,
            I => encoder0_position_target_22
        );

    \I__13060\ : LocalMux
    port map (
            O => \N__55259\,
            I => encoder0_position_target_22
        );

    \I__13059\ : InMux
    port map (
            O => \N__55252\,
            I => n12684
        );

    \I__13058\ : CascadeMux
    port map (
            O => \N__55249\,
            I => \N__55243\
        );

    \I__13057\ : CascadeMux
    port map (
            O => \N__55248\,
            I => \N__55240\
        );

    \I__13056\ : CascadeMux
    port map (
            O => \N__55247\,
            I => \N__55237\
        );

    \I__13055\ : CascadeMux
    port map (
            O => \N__55246\,
            I => \N__55230\
        );

    \I__13054\ : InMux
    port map (
            O => \N__55243\,
            I => \N__55202\
        );

    \I__13053\ : InMux
    port map (
            O => \N__55240\,
            I => \N__55202\
        );

    \I__13052\ : InMux
    port map (
            O => \N__55237\,
            I => \N__55202\
        );

    \I__13051\ : InMux
    port map (
            O => \N__55236\,
            I => \N__55193\
        );

    \I__13050\ : InMux
    port map (
            O => \N__55235\,
            I => \N__55193\
        );

    \I__13049\ : InMux
    port map (
            O => \N__55234\,
            I => \N__55193\
        );

    \I__13048\ : InMux
    port map (
            O => \N__55233\,
            I => \N__55193\
        );

    \I__13047\ : InMux
    port map (
            O => \N__55230\,
            I => \N__55180\
        );

    \I__13046\ : InMux
    port map (
            O => \N__55229\,
            I => \N__55180\
        );

    \I__13045\ : InMux
    port map (
            O => \N__55228\,
            I => \N__55175\
        );

    \I__13044\ : InMux
    port map (
            O => \N__55227\,
            I => \N__55175\
        );

    \I__13043\ : CascadeMux
    port map (
            O => \N__55226\,
            I => \N__55169\
        );

    \I__13042\ : InMux
    port map (
            O => \N__55225\,
            I => \N__55156\
        );

    \I__13041\ : InMux
    port map (
            O => \N__55224\,
            I => \N__55156\
        );

    \I__13040\ : InMux
    port map (
            O => \N__55223\,
            I => \N__55153\
        );

    \I__13039\ : InMux
    port map (
            O => \N__55222\,
            I => \N__55146\
        );

    \I__13038\ : InMux
    port map (
            O => \N__55221\,
            I => \N__55146\
        );

    \I__13037\ : InMux
    port map (
            O => \N__55220\,
            I => \N__55146\
        );

    \I__13036\ : CascadeMux
    port map (
            O => \N__55219\,
            I => \N__55142\
        );

    \I__13035\ : CascadeMux
    port map (
            O => \N__55218\,
            I => \N__55137\
        );

    \I__13034\ : CascadeMux
    port map (
            O => \N__55217\,
            I => \N__55118\
        );

    \I__13033\ : CascadeMux
    port map (
            O => \N__55216\,
            I => \N__55114\
        );

    \I__13032\ : CascadeMux
    port map (
            O => \N__55215\,
            I => \N__55110\
        );

    \I__13031\ : CascadeMux
    port map (
            O => \N__55214\,
            I => \N__55106\
        );

    \I__13030\ : CascadeMux
    port map (
            O => \N__55213\,
            I => \N__55103\
        );

    \I__13029\ : CascadeMux
    port map (
            O => \N__55212\,
            I => \N__55099\
        );

    \I__13028\ : CascadeMux
    port map (
            O => \N__55211\,
            I => \N__55095\
        );

    \I__13027\ : CascadeMux
    port map (
            O => \N__55210\,
            I => \N__55091\
        );

    \I__13026\ : CascadeMux
    port map (
            O => \N__55209\,
            I => \N__55073\
        );

    \I__13025\ : LocalMux
    port map (
            O => \N__55202\,
            I => \N__55057\
        );

    \I__13024\ : LocalMux
    port map (
            O => \N__55193\,
            I => \N__55054\
        );

    \I__13023\ : InMux
    port map (
            O => \N__55192\,
            I => \N__55047\
        );

    \I__13022\ : InMux
    port map (
            O => \N__55191\,
            I => \N__55047\
        );

    \I__13021\ : InMux
    port map (
            O => \N__55190\,
            I => \N__55047\
        );

    \I__13020\ : CascadeMux
    port map (
            O => \N__55189\,
            I => \N__55044\
        );

    \I__13019\ : CascadeMux
    port map (
            O => \N__55188\,
            I => \N__55041\
        );

    \I__13018\ : CascadeMux
    port map (
            O => \N__55187\,
            I => \N__55038\
        );

    \I__13017\ : CascadeMux
    port map (
            O => \N__55186\,
            I => \N__55035\
        );

    \I__13016\ : CascadeMux
    port map (
            O => \N__55185\,
            I => \N__55031\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__55180\,
            I => \N__55026\
        );

    \I__13014\ : LocalMux
    port map (
            O => \N__55175\,
            I => \N__55026\
        );

    \I__13013\ : InMux
    port map (
            O => \N__55174\,
            I => \N__55019\
        );

    \I__13012\ : InMux
    port map (
            O => \N__55173\,
            I => \N__55019\
        );

    \I__13011\ : InMux
    port map (
            O => \N__55172\,
            I => \N__55019\
        );

    \I__13010\ : InMux
    port map (
            O => \N__55169\,
            I => \N__55010\
        );

    \I__13009\ : InMux
    port map (
            O => \N__55168\,
            I => \N__55010\
        );

    \I__13008\ : InMux
    port map (
            O => \N__55167\,
            I => \N__55010\
        );

    \I__13007\ : InMux
    port map (
            O => \N__55166\,
            I => \N__55010\
        );

    \I__13006\ : InMux
    port map (
            O => \N__55165\,
            I => \N__55001\
        );

    \I__13005\ : InMux
    port map (
            O => \N__55164\,
            I => \N__55001\
        );

    \I__13004\ : InMux
    port map (
            O => \N__55163\,
            I => \N__55001\
        );

    \I__13003\ : InMux
    port map (
            O => \N__55162\,
            I => \N__55001\
        );

    \I__13002\ : CascadeMux
    port map (
            O => \N__55161\,
            I => \N__54998\
        );

    \I__13001\ : LocalMux
    port map (
            O => \N__55156\,
            I => \N__54968\
        );

    \I__13000\ : LocalMux
    port map (
            O => \N__55153\,
            I => \N__54968\
        );

    \I__12999\ : LocalMux
    port map (
            O => \N__55146\,
            I => \N__54968\
        );

    \I__12998\ : InMux
    port map (
            O => \N__55145\,
            I => \N__54959\
        );

    \I__12997\ : InMux
    port map (
            O => \N__55142\,
            I => \N__54959\
        );

    \I__12996\ : InMux
    port map (
            O => \N__55141\,
            I => \N__54959\
        );

    \I__12995\ : InMux
    port map (
            O => \N__55140\,
            I => \N__54959\
        );

    \I__12994\ : InMux
    port map (
            O => \N__55137\,
            I => \N__54952\
        );

    \I__12993\ : InMux
    port map (
            O => \N__55136\,
            I => \N__54952\
        );

    \I__12992\ : InMux
    port map (
            O => \N__55135\,
            I => \N__54952\
        );

    \I__12991\ : CascadeMux
    port map (
            O => \N__55134\,
            I => \N__54942\
        );

    \I__12990\ : CascadeMux
    port map (
            O => \N__55133\,
            I => \N__54931\
        );

    \I__12989\ : CascadeMux
    port map (
            O => \N__55132\,
            I => \N__54928\
        );

    \I__12988\ : CascadeMux
    port map (
            O => \N__55131\,
            I => \N__54917\
        );

    \I__12987\ : CascadeMux
    port map (
            O => \N__55130\,
            I => \N__54914\
        );

    \I__12986\ : CascadeMux
    port map (
            O => \N__55129\,
            I => \N__54911\
        );

    \I__12985\ : CascadeMux
    port map (
            O => \N__55128\,
            I => \N__54908\
        );

    \I__12984\ : CascadeMux
    port map (
            O => \N__55127\,
            I => \N__54905\
        );

    \I__12983\ : CascadeMux
    port map (
            O => \N__55126\,
            I => \N__54902\
        );

    \I__12982\ : CascadeMux
    port map (
            O => \N__55125\,
            I => \N__54899\
        );

    \I__12981\ : CascadeMux
    port map (
            O => \N__55124\,
            I => \N__54896\
        );

    \I__12980\ : CascadeMux
    port map (
            O => \N__55123\,
            I => \N__54893\
        );

    \I__12979\ : CascadeMux
    port map (
            O => \N__55122\,
            I => \N__54890\
        );

    \I__12978\ : InMux
    port map (
            O => \N__55121\,
            I => \N__54848\
        );

    \I__12977\ : InMux
    port map (
            O => \N__55118\,
            I => \N__54848\
        );

    \I__12976\ : InMux
    port map (
            O => \N__55117\,
            I => \N__54848\
        );

    \I__12975\ : InMux
    port map (
            O => \N__55114\,
            I => \N__54848\
        );

    \I__12974\ : InMux
    port map (
            O => \N__55113\,
            I => \N__54848\
        );

    \I__12973\ : InMux
    port map (
            O => \N__55110\,
            I => \N__54848\
        );

    \I__12972\ : InMux
    port map (
            O => \N__55109\,
            I => \N__54848\
        );

    \I__12971\ : InMux
    port map (
            O => \N__55106\,
            I => \N__54848\
        );

    \I__12970\ : InMux
    port map (
            O => \N__55103\,
            I => \N__54831\
        );

    \I__12969\ : InMux
    port map (
            O => \N__55102\,
            I => \N__54831\
        );

    \I__12968\ : InMux
    port map (
            O => \N__55099\,
            I => \N__54831\
        );

    \I__12967\ : InMux
    port map (
            O => \N__55098\,
            I => \N__54831\
        );

    \I__12966\ : InMux
    port map (
            O => \N__55095\,
            I => \N__54831\
        );

    \I__12965\ : InMux
    port map (
            O => \N__55094\,
            I => \N__54831\
        );

    \I__12964\ : InMux
    port map (
            O => \N__55091\,
            I => \N__54831\
        );

    \I__12963\ : InMux
    port map (
            O => \N__55090\,
            I => \N__54831\
        );

    \I__12962\ : CascadeMux
    port map (
            O => \N__55089\,
            I => \N__54828\
        );

    \I__12961\ : CascadeMux
    port map (
            O => \N__55088\,
            I => \N__54824\
        );

    \I__12960\ : CascadeMux
    port map (
            O => \N__55087\,
            I => \N__54820\
        );

    \I__12959\ : CascadeMux
    port map (
            O => \N__55086\,
            I => \N__54816\
        );

    \I__12958\ : CascadeMux
    port map (
            O => \N__55085\,
            I => \N__54812\
        );

    \I__12957\ : CascadeMux
    port map (
            O => \N__55084\,
            I => \N__54809\
        );

    \I__12956\ : CascadeMux
    port map (
            O => \N__55083\,
            I => \N__54806\
        );

    \I__12955\ : CascadeMux
    port map (
            O => \N__55082\,
            I => \N__54803\
        );

    \I__12954\ : CascadeMux
    port map (
            O => \N__55081\,
            I => \N__54800\
        );

    \I__12953\ : CascadeMux
    port map (
            O => \N__55080\,
            I => \N__54797\
        );

    \I__12952\ : CascadeMux
    port map (
            O => \N__55079\,
            I => \N__54794\
        );

    \I__12951\ : CascadeMux
    port map (
            O => \N__55078\,
            I => \N__54791\
        );

    \I__12950\ : CascadeMux
    port map (
            O => \N__55077\,
            I => \N__54788\
        );

    \I__12949\ : CascadeMux
    port map (
            O => \N__55076\,
            I => \N__54785\
        );

    \I__12948\ : InMux
    port map (
            O => \N__55073\,
            I => \N__54779\
        );

    \I__12947\ : InMux
    port map (
            O => \N__55072\,
            I => \N__54779\
        );

    \I__12946\ : InMux
    port map (
            O => \N__55071\,
            I => \N__54774\
        );

    \I__12945\ : InMux
    port map (
            O => \N__55070\,
            I => \N__54774\
        );

    \I__12944\ : InMux
    port map (
            O => \N__55069\,
            I => \N__54762\
        );

    \I__12943\ : InMux
    port map (
            O => \N__55068\,
            I => \N__54762\
        );

    \I__12942\ : InMux
    port map (
            O => \N__55067\,
            I => \N__54759\
        );

    \I__12941\ : InMux
    port map (
            O => \N__55066\,
            I => \N__54756\
        );

    \I__12940\ : InMux
    port map (
            O => \N__55065\,
            I => \N__54749\
        );

    \I__12939\ : InMux
    port map (
            O => \N__55064\,
            I => \N__54749\
        );

    \I__12938\ : InMux
    port map (
            O => \N__55063\,
            I => \N__54749\
        );

    \I__12937\ : CascadeMux
    port map (
            O => \N__55062\,
            I => \N__54745\
        );

    \I__12936\ : CascadeMux
    port map (
            O => \N__55061\,
            I => \N__54735\
        );

    \I__12935\ : InMux
    port map (
            O => \N__55060\,
            I => \N__54724\
        );

    \I__12934\ : Span4Mux_v
    port map (
            O => \N__55057\,
            I => \N__54717\
        );

    \I__12933\ : Span4Mux_h
    port map (
            O => \N__55054\,
            I => \N__54717\
        );

    \I__12932\ : LocalMux
    port map (
            O => \N__55047\,
            I => \N__54717\
        );

    \I__12931\ : InMux
    port map (
            O => \N__55044\,
            I => \N__54712\
        );

    \I__12930\ : InMux
    port map (
            O => \N__55041\,
            I => \N__54712\
        );

    \I__12929\ : InMux
    port map (
            O => \N__55038\,
            I => \N__54703\
        );

    \I__12928\ : InMux
    port map (
            O => \N__55035\,
            I => \N__54703\
        );

    \I__12927\ : InMux
    port map (
            O => \N__55034\,
            I => \N__54703\
        );

    \I__12926\ : InMux
    port map (
            O => \N__55031\,
            I => \N__54703\
        );

    \I__12925\ : Span4Mux_s3_v
    port map (
            O => \N__55026\,
            I => \N__54694\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__55019\,
            I => \N__54694\
        );

    \I__12923\ : LocalMux
    port map (
            O => \N__55010\,
            I => \N__54689\
        );

    \I__12922\ : LocalMux
    port map (
            O => \N__55001\,
            I => \N__54689\
        );

    \I__12921\ : InMux
    port map (
            O => \N__54998\,
            I => \N__54686\
        );

    \I__12920\ : CascadeMux
    port map (
            O => \N__54997\,
            I => \N__54683\
        );

    \I__12919\ : CascadeMux
    port map (
            O => \N__54996\,
            I => \N__54680\
        );

    \I__12918\ : CascadeMux
    port map (
            O => \N__54995\,
            I => \N__54673\
        );

    \I__12917\ : CascadeMux
    port map (
            O => \N__54994\,
            I => \N__54670\
        );

    \I__12916\ : CascadeMux
    port map (
            O => \N__54993\,
            I => \N__54665\
        );

    \I__12915\ : CascadeMux
    port map (
            O => \N__54992\,
            I => \N__54662\
        );

    \I__12914\ : CascadeMux
    port map (
            O => \N__54991\,
            I => \N__54659\
        );

    \I__12913\ : CascadeMux
    port map (
            O => \N__54990\,
            I => \N__54656\
        );

    \I__12912\ : CascadeMux
    port map (
            O => \N__54989\,
            I => \N__54653\
        );

    \I__12911\ : CascadeMux
    port map (
            O => \N__54988\,
            I => \N__54650\
        );

    \I__12910\ : CascadeMux
    port map (
            O => \N__54987\,
            I => \N__54646\
        );

    \I__12909\ : CascadeMux
    port map (
            O => \N__54986\,
            I => \N__54643\
        );

    \I__12908\ : CascadeMux
    port map (
            O => \N__54985\,
            I => \N__54640\
        );

    \I__12907\ : CascadeMux
    port map (
            O => \N__54984\,
            I => \N__54637\
        );

    \I__12906\ : CascadeMux
    port map (
            O => \N__54983\,
            I => \N__54634\
        );

    \I__12905\ : CascadeMux
    port map (
            O => \N__54982\,
            I => \N__54631\
        );

    \I__12904\ : CascadeMux
    port map (
            O => \N__54981\,
            I => \N__54628\
        );

    \I__12903\ : CascadeMux
    port map (
            O => \N__54980\,
            I => \N__54625\
        );

    \I__12902\ : CascadeMux
    port map (
            O => \N__54979\,
            I => \N__54622\
        );

    \I__12901\ : CascadeMux
    port map (
            O => \N__54978\,
            I => \N__54606\
        );

    \I__12900\ : CascadeMux
    port map (
            O => \N__54977\,
            I => \N__54600\
        );

    \I__12899\ : CascadeMux
    port map (
            O => \N__54976\,
            I => \N__54590\
        );

    \I__12898\ : CascadeMux
    port map (
            O => \N__54975\,
            I => \N__54586\
        );

    \I__12897\ : Span4Mux_s2_v
    port map (
            O => \N__54968\,
            I => \N__54573\
        );

    \I__12896\ : LocalMux
    port map (
            O => \N__54959\,
            I => \N__54573\
        );

    \I__12895\ : LocalMux
    port map (
            O => \N__54952\,
            I => \N__54573\
        );

    \I__12894\ : InMux
    port map (
            O => \N__54951\,
            I => \N__54570\
        );

    \I__12893\ : InMux
    port map (
            O => \N__54950\,
            I => \N__54567\
        );

    \I__12892\ : InMux
    port map (
            O => \N__54949\,
            I => \N__54560\
        );

    \I__12891\ : InMux
    port map (
            O => \N__54948\,
            I => \N__54560\
        );

    \I__12890\ : InMux
    port map (
            O => \N__54947\,
            I => \N__54560\
        );

    \I__12889\ : InMux
    port map (
            O => \N__54946\,
            I => \N__54549\
        );

    \I__12888\ : InMux
    port map (
            O => \N__54945\,
            I => \N__54549\
        );

    \I__12887\ : InMux
    port map (
            O => \N__54942\,
            I => \N__54549\
        );

    \I__12886\ : InMux
    port map (
            O => \N__54941\,
            I => \N__54549\
        );

    \I__12885\ : InMux
    port map (
            O => \N__54940\,
            I => \N__54549\
        );

    \I__12884\ : InMux
    port map (
            O => \N__54939\,
            I => \N__54546\
        );

    \I__12883\ : InMux
    port map (
            O => \N__54938\,
            I => \N__54539\
        );

    \I__12882\ : InMux
    port map (
            O => \N__54937\,
            I => \N__54539\
        );

    \I__12881\ : InMux
    port map (
            O => \N__54936\,
            I => \N__54539\
        );

    \I__12880\ : CascadeMux
    port map (
            O => \N__54935\,
            I => \N__54536\
        );

    \I__12879\ : CascadeMux
    port map (
            O => \N__54934\,
            I => \N__54532\
        );

    \I__12878\ : InMux
    port map (
            O => \N__54931\,
            I => \N__54522\
        );

    \I__12877\ : InMux
    port map (
            O => \N__54928\,
            I => \N__54522\
        );

    \I__12876\ : InMux
    port map (
            O => \N__54927\,
            I => \N__54522\
        );

    \I__12875\ : InMux
    port map (
            O => \N__54926\,
            I => \N__54522\
        );

    \I__12874\ : CascadeMux
    port map (
            O => \N__54925\,
            I => \N__54514\
        );

    \I__12873\ : CascadeMux
    port map (
            O => \N__54924\,
            I => \N__54511\
        );

    \I__12872\ : CascadeMux
    port map (
            O => \N__54923\,
            I => \N__54506\
        );

    \I__12871\ : CascadeMux
    port map (
            O => \N__54922\,
            I => \N__54502\
        );

    \I__12870\ : CascadeMux
    port map (
            O => \N__54921\,
            I => \N__54498\
        );

    \I__12869\ : CascadeMux
    port map (
            O => \N__54920\,
            I => \N__54495\
        );

    \I__12868\ : InMux
    port map (
            O => \N__54917\,
            I => \N__54488\
        );

    \I__12867\ : InMux
    port map (
            O => \N__54914\,
            I => \N__54488\
        );

    \I__12866\ : InMux
    port map (
            O => \N__54911\,
            I => \N__54488\
        );

    \I__12865\ : InMux
    port map (
            O => \N__54908\,
            I => \N__54479\
        );

    \I__12864\ : InMux
    port map (
            O => \N__54905\,
            I => \N__54479\
        );

    \I__12863\ : InMux
    port map (
            O => \N__54902\,
            I => \N__54479\
        );

    \I__12862\ : InMux
    port map (
            O => \N__54899\,
            I => \N__54479\
        );

    \I__12861\ : InMux
    port map (
            O => \N__54896\,
            I => \N__54472\
        );

    \I__12860\ : InMux
    port map (
            O => \N__54893\,
            I => \N__54472\
        );

    \I__12859\ : InMux
    port map (
            O => \N__54890\,
            I => \N__54472\
        );

    \I__12858\ : CascadeMux
    port map (
            O => \N__54889\,
            I => \N__54468\
        );

    \I__12857\ : CascadeMux
    port map (
            O => \N__54888\,
            I => \N__54465\
        );

    \I__12856\ : CascadeMux
    port map (
            O => \N__54887\,
            I => \N__54462\
        );

    \I__12855\ : CascadeMux
    port map (
            O => \N__54886\,
            I => \N__54459\
        );

    \I__12854\ : CascadeMux
    port map (
            O => \N__54885\,
            I => \N__54456\
        );

    \I__12853\ : CascadeMux
    port map (
            O => \N__54884\,
            I => \N__54453\
        );

    \I__12852\ : CascadeMux
    port map (
            O => \N__54883\,
            I => \N__54450\
        );

    \I__12851\ : CascadeMux
    port map (
            O => \N__54882\,
            I => \N__54447\
        );

    \I__12850\ : CascadeMux
    port map (
            O => \N__54881\,
            I => \N__54444\
        );

    \I__12849\ : CascadeMux
    port map (
            O => \N__54880\,
            I => \N__54441\
        );

    \I__12848\ : CascadeMux
    port map (
            O => \N__54879\,
            I => \N__54438\
        );

    \I__12847\ : CascadeMux
    port map (
            O => \N__54878\,
            I => \N__54435\
        );

    \I__12846\ : CascadeMux
    port map (
            O => \N__54877\,
            I => \N__54432\
        );

    \I__12845\ : CascadeMux
    port map (
            O => \N__54876\,
            I => \N__54428\
        );

    \I__12844\ : CascadeMux
    port map (
            O => \N__54875\,
            I => \N__54425\
        );

    \I__12843\ : CascadeMux
    port map (
            O => \N__54874\,
            I => \N__54422\
        );

    \I__12842\ : CascadeMux
    port map (
            O => \N__54873\,
            I => \N__54419\
        );

    \I__12841\ : CascadeMux
    port map (
            O => \N__54872\,
            I => \N__54416\
        );

    \I__12840\ : CascadeMux
    port map (
            O => \N__54871\,
            I => \N__54413\
        );

    \I__12839\ : CascadeMux
    port map (
            O => \N__54870\,
            I => \N__54410\
        );

    \I__12838\ : CascadeMux
    port map (
            O => \N__54869\,
            I => \N__54407\
        );

    \I__12837\ : CascadeMux
    port map (
            O => \N__54868\,
            I => \N__54404\
        );

    \I__12836\ : CascadeMux
    port map (
            O => \N__54867\,
            I => \N__54400\
        );

    \I__12835\ : CascadeMux
    port map (
            O => \N__54866\,
            I => \N__54397\
        );

    \I__12834\ : CascadeMux
    port map (
            O => \N__54865\,
            I => \N__54394\
        );

    \I__12833\ : LocalMux
    port map (
            O => \N__54848\,
            I => \N__54389\
        );

    \I__12832\ : LocalMux
    port map (
            O => \N__54831\,
            I => \N__54389\
        );

    \I__12831\ : InMux
    port map (
            O => \N__54828\,
            I => \N__54374\
        );

    \I__12830\ : InMux
    port map (
            O => \N__54827\,
            I => \N__54374\
        );

    \I__12829\ : InMux
    port map (
            O => \N__54824\,
            I => \N__54374\
        );

    \I__12828\ : InMux
    port map (
            O => \N__54823\,
            I => \N__54374\
        );

    \I__12827\ : InMux
    port map (
            O => \N__54820\,
            I => \N__54374\
        );

    \I__12826\ : InMux
    port map (
            O => \N__54819\,
            I => \N__54374\
        );

    \I__12825\ : InMux
    port map (
            O => \N__54816\,
            I => \N__54374\
        );

    \I__12824\ : InMux
    port map (
            O => \N__54815\,
            I => \N__54367\
        );

    \I__12823\ : InMux
    port map (
            O => \N__54812\,
            I => \N__54367\
        );

    \I__12822\ : InMux
    port map (
            O => \N__54809\,
            I => \N__54367\
        );

    \I__12821\ : InMux
    port map (
            O => \N__54806\,
            I => \N__54358\
        );

    \I__12820\ : InMux
    port map (
            O => \N__54803\,
            I => \N__54358\
        );

    \I__12819\ : InMux
    port map (
            O => \N__54800\,
            I => \N__54358\
        );

    \I__12818\ : InMux
    port map (
            O => \N__54797\,
            I => \N__54358\
        );

    \I__12817\ : InMux
    port map (
            O => \N__54794\,
            I => \N__54347\
        );

    \I__12816\ : InMux
    port map (
            O => \N__54791\,
            I => \N__54347\
        );

    \I__12815\ : InMux
    port map (
            O => \N__54788\,
            I => \N__54347\
        );

    \I__12814\ : InMux
    port map (
            O => \N__54785\,
            I => \N__54347\
        );

    \I__12813\ : InMux
    port map (
            O => \N__54784\,
            I => \N__54347\
        );

    \I__12812\ : LocalMux
    port map (
            O => \N__54779\,
            I => \N__54331\
        );

    \I__12811\ : LocalMux
    port map (
            O => \N__54774\,
            I => \N__54331\
        );

    \I__12810\ : InMux
    port map (
            O => \N__54773\,
            I => \N__54324\
        );

    \I__12809\ : InMux
    port map (
            O => \N__54772\,
            I => \N__54324\
        );

    \I__12808\ : InMux
    port map (
            O => \N__54771\,
            I => \N__54324\
        );

    \I__12807\ : CascadeMux
    port map (
            O => \N__54770\,
            I => \N__54318\
        );

    \I__12806\ : CascadeMux
    port map (
            O => \N__54769\,
            I => \N__54315\
        );

    \I__12805\ : CascadeMux
    port map (
            O => \N__54768\,
            I => \N__54312\
        );

    \I__12804\ : CascadeMux
    port map (
            O => \N__54767\,
            I => \N__54309\
        );

    \I__12803\ : LocalMux
    port map (
            O => \N__54762\,
            I => \N__54299\
        );

    \I__12802\ : LocalMux
    port map (
            O => \N__54759\,
            I => \N__54299\
        );

    \I__12801\ : LocalMux
    port map (
            O => \N__54756\,
            I => \N__54299\
        );

    \I__12800\ : LocalMux
    port map (
            O => \N__54749\,
            I => \N__54299\
        );

    \I__12799\ : InMux
    port map (
            O => \N__54748\,
            I => \N__54292\
        );

    \I__12798\ : InMux
    port map (
            O => \N__54745\,
            I => \N__54292\
        );

    \I__12797\ : InMux
    port map (
            O => \N__54744\,
            I => \N__54292\
        );

    \I__12796\ : InMux
    port map (
            O => \N__54743\,
            I => \N__54287\
        );

    \I__12795\ : InMux
    port map (
            O => \N__54742\,
            I => \N__54287\
        );

    \I__12794\ : InMux
    port map (
            O => \N__54741\,
            I => \N__54284\
        );

    \I__12793\ : InMux
    port map (
            O => \N__54740\,
            I => \N__54277\
        );

    \I__12792\ : InMux
    port map (
            O => \N__54739\,
            I => \N__54277\
        );

    \I__12791\ : InMux
    port map (
            O => \N__54738\,
            I => \N__54277\
        );

    \I__12790\ : InMux
    port map (
            O => \N__54735\,
            I => \N__54272\
        );

    \I__12789\ : InMux
    port map (
            O => \N__54734\,
            I => \N__54272\
        );

    \I__12788\ : InMux
    port map (
            O => \N__54733\,
            I => \N__54267\
        );

    \I__12787\ : InMux
    port map (
            O => \N__54732\,
            I => \N__54267\
        );

    \I__12786\ : CascadeMux
    port map (
            O => \N__54731\,
            I => \N__54263\
        );

    \I__12785\ : CascadeMux
    port map (
            O => \N__54730\,
            I => \N__54260\
        );

    \I__12784\ : CascadeMux
    port map (
            O => \N__54729\,
            I => \N__54257\
        );

    \I__12783\ : CascadeMux
    port map (
            O => \N__54728\,
            I => \N__54245\
        );

    \I__12782\ : CascadeMux
    port map (
            O => \N__54727\,
            I => \N__54242\
        );

    \I__12781\ : LocalMux
    port map (
            O => \N__54724\,
            I => \N__54235\
        );

    \I__12780\ : Span4Mux_v
    port map (
            O => \N__54717\,
            I => \N__54235\
        );

    \I__12779\ : LocalMux
    port map (
            O => \N__54712\,
            I => \N__54230\
        );

    \I__12778\ : LocalMux
    port map (
            O => \N__54703\,
            I => \N__54230\
        );

    \I__12777\ : InMux
    port map (
            O => \N__54702\,
            I => \N__54227\
        );

    \I__12776\ : InMux
    port map (
            O => \N__54701\,
            I => \N__54220\
        );

    \I__12775\ : InMux
    port map (
            O => \N__54700\,
            I => \N__54220\
        );

    \I__12774\ : InMux
    port map (
            O => \N__54699\,
            I => \N__54220\
        );

    \I__12773\ : Span4Mux_v
    port map (
            O => \N__54694\,
            I => \N__54213\
        );

    \I__12772\ : Span4Mux_h
    port map (
            O => \N__54689\,
            I => \N__54213\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__54686\,
            I => \N__54213\
        );

    \I__12770\ : InMux
    port map (
            O => \N__54683\,
            I => \N__54204\
        );

    \I__12769\ : InMux
    port map (
            O => \N__54680\,
            I => \N__54204\
        );

    \I__12768\ : InMux
    port map (
            O => \N__54679\,
            I => \N__54204\
        );

    \I__12767\ : InMux
    port map (
            O => \N__54678\,
            I => \N__54204\
        );

    \I__12766\ : CascadeMux
    port map (
            O => \N__54677\,
            I => \N__54201\
        );

    \I__12765\ : CascadeMux
    port map (
            O => \N__54676\,
            I => \N__54198\
        );

    \I__12764\ : InMux
    port map (
            O => \N__54673\,
            I => \N__54191\
        );

    \I__12763\ : InMux
    port map (
            O => \N__54670\,
            I => \N__54191\
        );

    \I__12762\ : InMux
    port map (
            O => \N__54669\,
            I => \N__54191\
        );

    \I__12761\ : InMux
    port map (
            O => \N__54668\,
            I => \N__54186\
        );

    \I__12760\ : InMux
    port map (
            O => \N__54665\,
            I => \N__54186\
        );

    \I__12759\ : InMux
    port map (
            O => \N__54662\,
            I => \N__54183\
        );

    \I__12758\ : InMux
    port map (
            O => \N__54659\,
            I => \N__54172\
        );

    \I__12757\ : InMux
    port map (
            O => \N__54656\,
            I => \N__54172\
        );

    \I__12756\ : InMux
    port map (
            O => \N__54653\,
            I => \N__54172\
        );

    \I__12755\ : InMux
    port map (
            O => \N__54650\,
            I => \N__54172\
        );

    \I__12754\ : InMux
    port map (
            O => \N__54649\,
            I => \N__54172\
        );

    \I__12753\ : InMux
    port map (
            O => \N__54646\,
            I => \N__54163\
        );

    \I__12752\ : InMux
    port map (
            O => \N__54643\,
            I => \N__54163\
        );

    \I__12751\ : InMux
    port map (
            O => \N__54640\,
            I => \N__54163\
        );

    \I__12750\ : InMux
    port map (
            O => \N__54637\,
            I => \N__54163\
        );

    \I__12749\ : InMux
    port map (
            O => \N__54634\,
            I => \N__54154\
        );

    \I__12748\ : InMux
    port map (
            O => \N__54631\,
            I => \N__54154\
        );

    \I__12747\ : InMux
    port map (
            O => \N__54628\,
            I => \N__54154\
        );

    \I__12746\ : InMux
    port map (
            O => \N__54625\,
            I => \N__54154\
        );

    \I__12745\ : InMux
    port map (
            O => \N__54622\,
            I => \N__54143\
        );

    \I__12744\ : InMux
    port map (
            O => \N__54621\,
            I => \N__54143\
        );

    \I__12743\ : InMux
    port map (
            O => \N__54620\,
            I => \N__54143\
        );

    \I__12742\ : InMux
    port map (
            O => \N__54619\,
            I => \N__54143\
        );

    \I__12741\ : InMux
    port map (
            O => \N__54618\,
            I => \N__54143\
        );

    \I__12740\ : InMux
    port map (
            O => \N__54617\,
            I => \N__54134\
        );

    \I__12739\ : InMux
    port map (
            O => \N__54616\,
            I => \N__54134\
        );

    \I__12738\ : InMux
    port map (
            O => \N__54615\,
            I => \N__54134\
        );

    \I__12737\ : InMux
    port map (
            O => \N__54614\,
            I => \N__54134\
        );

    \I__12736\ : InMux
    port map (
            O => \N__54613\,
            I => \N__54131\
        );

    \I__12735\ : InMux
    port map (
            O => \N__54612\,
            I => \N__54124\
        );

    \I__12734\ : InMux
    port map (
            O => \N__54611\,
            I => \N__54124\
        );

    \I__12733\ : InMux
    port map (
            O => \N__54610\,
            I => \N__54124\
        );

    \I__12732\ : InMux
    port map (
            O => \N__54609\,
            I => \N__54119\
        );

    \I__12731\ : InMux
    port map (
            O => \N__54606\,
            I => \N__54119\
        );

    \I__12730\ : CascadeMux
    port map (
            O => \N__54605\,
            I => \N__54116\
        );

    \I__12729\ : CascadeMux
    port map (
            O => \N__54604\,
            I => \N__54112\
        );

    \I__12728\ : CascadeMux
    port map (
            O => \N__54603\,
            I => \N__54109\
        );

    \I__12727\ : InMux
    port map (
            O => \N__54600\,
            I => \N__54106\
        );

    \I__12726\ : InMux
    port map (
            O => \N__54599\,
            I => \N__54103\
        );

    \I__12725\ : InMux
    port map (
            O => \N__54598\,
            I => \N__54100\
        );

    \I__12724\ : InMux
    port map (
            O => \N__54597\,
            I => \N__54095\
        );

    \I__12723\ : InMux
    port map (
            O => \N__54596\,
            I => \N__54095\
        );

    \I__12722\ : InMux
    port map (
            O => \N__54595\,
            I => \N__54090\
        );

    \I__12721\ : InMux
    port map (
            O => \N__54594\,
            I => \N__54090\
        );

    \I__12720\ : InMux
    port map (
            O => \N__54593\,
            I => \N__54085\
        );

    \I__12719\ : InMux
    port map (
            O => \N__54590\,
            I => \N__54085\
        );

    \I__12718\ : CascadeMux
    port map (
            O => \N__54589\,
            I => \N__54079\
        );

    \I__12717\ : InMux
    port map (
            O => \N__54586\,
            I => \N__54070\
        );

    \I__12716\ : InMux
    port map (
            O => \N__54585\,
            I => \N__54070\
        );

    \I__12715\ : InMux
    port map (
            O => \N__54584\,
            I => \N__54070\
        );

    \I__12714\ : InMux
    port map (
            O => \N__54583\,
            I => \N__54063\
        );

    \I__12713\ : InMux
    port map (
            O => \N__54582\,
            I => \N__54063\
        );

    \I__12712\ : InMux
    port map (
            O => \N__54581\,
            I => \N__54063\
        );

    \I__12711\ : InMux
    port map (
            O => \N__54580\,
            I => \N__54060\
        );

    \I__12710\ : Span4Mux_v
    port map (
            O => \N__54573\,
            I => \N__54042\
        );

    \I__12709\ : LocalMux
    port map (
            O => \N__54570\,
            I => \N__54042\
        );

    \I__12708\ : LocalMux
    port map (
            O => \N__54567\,
            I => \N__54042\
        );

    \I__12707\ : LocalMux
    port map (
            O => \N__54560\,
            I => \N__54042\
        );

    \I__12706\ : LocalMux
    port map (
            O => \N__54549\,
            I => \N__54042\
        );

    \I__12705\ : LocalMux
    port map (
            O => \N__54546\,
            I => \N__54042\
        );

    \I__12704\ : LocalMux
    port map (
            O => \N__54539\,
            I => \N__54042\
        );

    \I__12703\ : InMux
    port map (
            O => \N__54536\,
            I => \N__54039\
        );

    \I__12702\ : InMux
    port map (
            O => \N__54535\,
            I => \N__54034\
        );

    \I__12701\ : InMux
    port map (
            O => \N__54532\,
            I => \N__54034\
        );

    \I__12700\ : InMux
    port map (
            O => \N__54531\,
            I => \N__54031\
        );

    \I__12699\ : LocalMux
    port map (
            O => \N__54522\,
            I => \N__54028\
        );

    \I__12698\ : InMux
    port map (
            O => \N__54521\,
            I => \N__54025\
        );

    \I__12697\ : InMux
    port map (
            O => \N__54520\,
            I => \N__54018\
        );

    \I__12696\ : InMux
    port map (
            O => \N__54519\,
            I => \N__54018\
        );

    \I__12695\ : InMux
    port map (
            O => \N__54518\,
            I => \N__54018\
        );

    \I__12694\ : InMux
    port map (
            O => \N__54517\,
            I => \N__54013\
        );

    \I__12693\ : InMux
    port map (
            O => \N__54514\,
            I => \N__54013\
        );

    \I__12692\ : InMux
    port map (
            O => \N__54511\,
            I => \N__53998\
        );

    \I__12691\ : InMux
    port map (
            O => \N__54510\,
            I => \N__53998\
        );

    \I__12690\ : InMux
    port map (
            O => \N__54509\,
            I => \N__53998\
        );

    \I__12689\ : InMux
    port map (
            O => \N__54506\,
            I => \N__53998\
        );

    \I__12688\ : InMux
    port map (
            O => \N__54505\,
            I => \N__53998\
        );

    \I__12687\ : InMux
    port map (
            O => \N__54502\,
            I => \N__53998\
        );

    \I__12686\ : InMux
    port map (
            O => \N__54501\,
            I => \N__53998\
        );

    \I__12685\ : InMux
    port map (
            O => \N__54498\,
            I => \N__53993\
        );

    \I__12684\ : InMux
    port map (
            O => \N__54495\,
            I => \N__53993\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__54488\,
            I => \N__53983\
        );

    \I__12682\ : LocalMux
    port map (
            O => \N__54479\,
            I => \N__53983\
        );

    \I__12681\ : LocalMux
    port map (
            O => \N__54472\,
            I => \N__53983\
        );

    \I__12680\ : InMux
    port map (
            O => \N__54471\,
            I => \N__53974\
        );

    \I__12679\ : InMux
    port map (
            O => \N__54468\,
            I => \N__53974\
        );

    \I__12678\ : InMux
    port map (
            O => \N__54465\,
            I => \N__53974\
        );

    \I__12677\ : InMux
    port map (
            O => \N__54462\,
            I => \N__53974\
        );

    \I__12676\ : InMux
    port map (
            O => \N__54459\,
            I => \N__53965\
        );

    \I__12675\ : InMux
    port map (
            O => \N__54456\,
            I => \N__53965\
        );

    \I__12674\ : InMux
    port map (
            O => \N__54453\,
            I => \N__53965\
        );

    \I__12673\ : InMux
    port map (
            O => \N__54450\,
            I => \N__53965\
        );

    \I__12672\ : InMux
    port map (
            O => \N__54447\,
            I => \N__53958\
        );

    \I__12671\ : InMux
    port map (
            O => \N__54444\,
            I => \N__53958\
        );

    \I__12670\ : InMux
    port map (
            O => \N__54441\,
            I => \N__53958\
        );

    \I__12669\ : InMux
    port map (
            O => \N__54438\,
            I => \N__53947\
        );

    \I__12668\ : InMux
    port map (
            O => \N__54435\,
            I => \N__53947\
        );

    \I__12667\ : InMux
    port map (
            O => \N__54432\,
            I => \N__53947\
        );

    \I__12666\ : InMux
    port map (
            O => \N__54431\,
            I => \N__53947\
        );

    \I__12665\ : InMux
    port map (
            O => \N__54428\,
            I => \N__53947\
        );

    \I__12664\ : InMux
    port map (
            O => \N__54425\,
            I => \N__53938\
        );

    \I__12663\ : InMux
    port map (
            O => \N__54422\,
            I => \N__53938\
        );

    \I__12662\ : InMux
    port map (
            O => \N__54419\,
            I => \N__53938\
        );

    \I__12661\ : InMux
    port map (
            O => \N__54416\,
            I => \N__53938\
        );

    \I__12660\ : InMux
    port map (
            O => \N__54413\,
            I => \N__53929\
        );

    \I__12659\ : InMux
    port map (
            O => \N__54410\,
            I => \N__53929\
        );

    \I__12658\ : InMux
    port map (
            O => \N__54407\,
            I => \N__53929\
        );

    \I__12657\ : InMux
    port map (
            O => \N__54404\,
            I => \N__53929\
        );

    \I__12656\ : InMux
    port map (
            O => \N__54403\,
            I => \N__53920\
        );

    \I__12655\ : InMux
    port map (
            O => \N__54400\,
            I => \N__53920\
        );

    \I__12654\ : InMux
    port map (
            O => \N__54397\,
            I => \N__53920\
        );

    \I__12653\ : InMux
    port map (
            O => \N__54394\,
            I => \N__53920\
        );

    \I__12652\ : Span4Mux_v
    port map (
            O => \N__54389\,
            I => \N__53909\
        );

    \I__12651\ : LocalMux
    port map (
            O => \N__54374\,
            I => \N__53909\
        );

    \I__12650\ : LocalMux
    port map (
            O => \N__54367\,
            I => \N__53909\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__54358\,
            I => \N__53909\
        );

    \I__12648\ : LocalMux
    port map (
            O => \N__54347\,
            I => \N__53909\
        );

    \I__12647\ : InMux
    port map (
            O => \N__54346\,
            I => \N__53906\
        );

    \I__12646\ : InMux
    port map (
            O => \N__54345\,
            I => \N__53899\
        );

    \I__12645\ : InMux
    port map (
            O => \N__54344\,
            I => \N__53899\
        );

    \I__12644\ : InMux
    port map (
            O => \N__54343\,
            I => \N__53899\
        );

    \I__12643\ : InMux
    port map (
            O => \N__54342\,
            I => \N__53892\
        );

    \I__12642\ : InMux
    port map (
            O => \N__54341\,
            I => \N__53892\
        );

    \I__12641\ : InMux
    port map (
            O => \N__54340\,
            I => \N__53892\
        );

    \I__12640\ : CascadeMux
    port map (
            O => \N__54339\,
            I => \N__53887\
        );

    \I__12639\ : CascadeMux
    port map (
            O => \N__54338\,
            I => \N__53884\
        );

    \I__12638\ : CascadeMux
    port map (
            O => \N__54337\,
            I => \N__53881\
        );

    \I__12637\ : CascadeMux
    port map (
            O => \N__54336\,
            I => \N__53878\
        );

    \I__12636\ : Span4Mux_h
    port map (
            O => \N__54331\,
            I => \N__53872\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__54324\,
            I => \N__53872\
        );

    \I__12634\ : CascadeMux
    port map (
            O => \N__54323\,
            I => \N__53866\
        );

    \I__12633\ : CascadeMux
    port map (
            O => \N__54322\,
            I => \N__53862\
        );

    \I__12632\ : CascadeMux
    port map (
            O => \N__54321\,
            I => \N__53855\
        );

    \I__12631\ : InMux
    port map (
            O => \N__54318\,
            I => \N__53852\
        );

    \I__12630\ : InMux
    port map (
            O => \N__54315\,
            I => \N__53845\
        );

    \I__12629\ : InMux
    port map (
            O => \N__54312\,
            I => \N__53845\
        );

    \I__12628\ : InMux
    port map (
            O => \N__54309\,
            I => \N__53845\
        );

    \I__12627\ : CascadeMux
    port map (
            O => \N__54308\,
            I => \N__53842\
        );

    \I__12626\ : Span4Mux_s3_v
    port map (
            O => \N__54299\,
            I => \N__53822\
        );

    \I__12625\ : LocalMux
    port map (
            O => \N__54292\,
            I => \N__53822\
        );

    \I__12624\ : LocalMux
    port map (
            O => \N__54287\,
            I => \N__53811\
        );

    \I__12623\ : LocalMux
    port map (
            O => \N__54284\,
            I => \N__53811\
        );

    \I__12622\ : LocalMux
    port map (
            O => \N__54277\,
            I => \N__53811\
        );

    \I__12621\ : LocalMux
    port map (
            O => \N__54272\,
            I => \N__53811\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__54267\,
            I => \N__53811\
        );

    \I__12619\ : InMux
    port map (
            O => \N__54266\,
            I => \N__53808\
        );

    \I__12618\ : InMux
    port map (
            O => \N__54263\,
            I => \N__53805\
        );

    \I__12617\ : InMux
    port map (
            O => \N__54260\,
            I => \N__53796\
        );

    \I__12616\ : InMux
    port map (
            O => \N__54257\,
            I => \N__53796\
        );

    \I__12615\ : InMux
    port map (
            O => \N__54256\,
            I => \N__53796\
        );

    \I__12614\ : InMux
    port map (
            O => \N__54255\,
            I => \N__53796\
        );

    \I__12613\ : InMux
    port map (
            O => \N__54254\,
            I => \N__53793\
        );

    \I__12612\ : CascadeMux
    port map (
            O => \N__54253\,
            I => \N__53786\
        );

    \I__12611\ : CascadeMux
    port map (
            O => \N__54252\,
            I => \N__53783\
        );

    \I__12610\ : CascadeMux
    port map (
            O => \N__54251\,
            I => \N__53780\
        );

    \I__12609\ : CascadeMux
    port map (
            O => \N__54250\,
            I => \N__53777\
        );

    \I__12608\ : CascadeMux
    port map (
            O => \N__54249\,
            I => \N__53774\
        );

    \I__12607\ : CascadeMux
    port map (
            O => \N__54248\,
            I => \N__53770\
        );

    \I__12606\ : InMux
    port map (
            O => \N__54245\,
            I => \N__53755\
        );

    \I__12605\ : InMux
    port map (
            O => \N__54242\,
            I => \N__53755\
        );

    \I__12604\ : InMux
    port map (
            O => \N__54241\,
            I => \N__53755\
        );

    \I__12603\ : InMux
    port map (
            O => \N__54240\,
            I => \N__53755\
        );

    \I__12602\ : Span4Mux_h
    port map (
            O => \N__54235\,
            I => \N__53742\
        );

    \I__12601\ : Span4Mux_v
    port map (
            O => \N__54230\,
            I => \N__53742\
        );

    \I__12600\ : LocalMux
    port map (
            O => \N__54227\,
            I => \N__53742\
        );

    \I__12599\ : LocalMux
    port map (
            O => \N__54220\,
            I => \N__53742\
        );

    \I__12598\ : Span4Mux_v
    port map (
            O => \N__54213\,
            I => \N__53742\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__54204\,
            I => \N__53742\
        );

    \I__12596\ : InMux
    port map (
            O => \N__54201\,
            I => \N__53737\
        );

    \I__12595\ : InMux
    port map (
            O => \N__54198\,
            I => \N__53737\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__54191\,
            I => \N__53719\
        );

    \I__12593\ : LocalMux
    port map (
            O => \N__54186\,
            I => \N__53719\
        );

    \I__12592\ : LocalMux
    port map (
            O => \N__54183\,
            I => \N__53719\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__54172\,
            I => \N__53719\
        );

    \I__12590\ : LocalMux
    port map (
            O => \N__54163\,
            I => \N__53719\
        );

    \I__12589\ : LocalMux
    port map (
            O => \N__54154\,
            I => \N__53719\
        );

    \I__12588\ : LocalMux
    port map (
            O => \N__54143\,
            I => \N__53719\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__54134\,
            I => \N__53719\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__54131\,
            I => \N__53714\
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__54124\,
            I => \N__53714\
        );

    \I__12584\ : LocalMux
    port map (
            O => \N__54119\,
            I => \N__53711\
        );

    \I__12583\ : InMux
    port map (
            O => \N__54116\,
            I => \N__53702\
        );

    \I__12582\ : InMux
    port map (
            O => \N__54115\,
            I => \N__53702\
        );

    \I__12581\ : InMux
    port map (
            O => \N__54112\,
            I => \N__53702\
        );

    \I__12580\ : InMux
    port map (
            O => \N__54109\,
            I => \N__53702\
        );

    \I__12579\ : LocalMux
    port map (
            O => \N__54106\,
            I => \N__53697\
        );

    \I__12578\ : LocalMux
    port map (
            O => \N__54103\,
            I => \N__53697\
        );

    \I__12577\ : LocalMux
    port map (
            O => \N__54100\,
            I => \N__53690\
        );

    \I__12576\ : LocalMux
    port map (
            O => \N__54095\,
            I => \N__53690\
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__54090\,
            I => \N__53690\
        );

    \I__12574\ : LocalMux
    port map (
            O => \N__54085\,
            I => \N__53687\
        );

    \I__12573\ : InMux
    port map (
            O => \N__54084\,
            I => \N__53682\
        );

    \I__12572\ : InMux
    port map (
            O => \N__54083\,
            I => \N__53682\
        );

    \I__12571\ : InMux
    port map (
            O => \N__54082\,
            I => \N__53677\
        );

    \I__12570\ : InMux
    port map (
            O => \N__54079\,
            I => \N__53677\
        );

    \I__12569\ : CascadeMux
    port map (
            O => \N__54078\,
            I => \N__53673\
        );

    \I__12568\ : CascadeMux
    port map (
            O => \N__54077\,
            I => \N__53669\
        );

    \I__12567\ : LocalMux
    port map (
            O => \N__54070\,
            I => \N__53659\
        );

    \I__12566\ : LocalMux
    port map (
            O => \N__54063\,
            I => \N__53654\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__54060\,
            I => \N__53654\
        );

    \I__12564\ : InMux
    port map (
            O => \N__54059\,
            I => \N__53647\
        );

    \I__12563\ : InMux
    port map (
            O => \N__54058\,
            I => \N__53647\
        );

    \I__12562\ : InMux
    port map (
            O => \N__54057\,
            I => \N__53647\
        );

    \I__12561\ : Span4Mux_v
    port map (
            O => \N__54042\,
            I => \N__53630\
        );

    \I__12560\ : LocalMux
    port map (
            O => \N__54039\,
            I => \N__53630\
        );

    \I__12559\ : LocalMux
    port map (
            O => \N__54034\,
            I => \N__53630\
        );

    \I__12558\ : LocalMux
    port map (
            O => \N__54031\,
            I => \N__53630\
        );

    \I__12557\ : Span4Mux_h
    port map (
            O => \N__54028\,
            I => \N__53630\
        );

    \I__12556\ : LocalMux
    port map (
            O => \N__54025\,
            I => \N__53630\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__54018\,
            I => \N__53630\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__54013\,
            I => \N__53630\
        );

    \I__12553\ : LocalMux
    port map (
            O => \N__53998\,
            I => \N__53625\
        );

    \I__12552\ : LocalMux
    port map (
            O => \N__53993\,
            I => \N__53625\
        );

    \I__12551\ : CascadeMux
    port map (
            O => \N__53992\,
            I => \N__53622\
        );

    \I__12550\ : CascadeMux
    port map (
            O => \N__53991\,
            I => \N__53617\
        );

    \I__12549\ : CascadeMux
    port map (
            O => \N__53990\,
            I => \N__53612\
        );

    \I__12548\ : Span4Mux_v
    port map (
            O => \N__53983\,
            I => \N__53608\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__53974\,
            I => \N__53593\
        );

    \I__12546\ : LocalMux
    port map (
            O => \N__53965\,
            I => \N__53593\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__53958\,
            I => \N__53593\
        );

    \I__12544\ : LocalMux
    port map (
            O => \N__53947\,
            I => \N__53593\
        );

    \I__12543\ : LocalMux
    port map (
            O => \N__53938\,
            I => \N__53593\
        );

    \I__12542\ : LocalMux
    port map (
            O => \N__53929\,
            I => \N__53593\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__53920\,
            I => \N__53593\
        );

    \I__12540\ : Span4Mux_v
    port map (
            O => \N__53909\,
            I => \N__53584\
        );

    \I__12539\ : LocalMux
    port map (
            O => \N__53906\,
            I => \N__53584\
        );

    \I__12538\ : LocalMux
    port map (
            O => \N__53899\,
            I => \N__53584\
        );

    \I__12537\ : LocalMux
    port map (
            O => \N__53892\,
            I => \N__53584\
        );

    \I__12536\ : InMux
    port map (
            O => \N__53891\,
            I => \N__53581\
        );

    \I__12535\ : InMux
    port map (
            O => \N__53890\,
            I => \N__53570\
        );

    \I__12534\ : InMux
    port map (
            O => \N__53887\,
            I => \N__53570\
        );

    \I__12533\ : InMux
    port map (
            O => \N__53884\,
            I => \N__53570\
        );

    \I__12532\ : InMux
    port map (
            O => \N__53881\,
            I => \N__53570\
        );

    \I__12531\ : InMux
    port map (
            O => \N__53878\,
            I => \N__53570\
        );

    \I__12530\ : CascadeMux
    port map (
            O => \N__53877\,
            I => \N__53566\
        );

    \I__12529\ : Span4Mux_v
    port map (
            O => \N__53872\,
            I => \N__53557\
        );

    \I__12528\ : CascadeMux
    port map (
            O => \N__53871\,
            I => \N__53554\
        );

    \I__12527\ : CascadeMux
    port map (
            O => \N__53870\,
            I => \N__53551\
        );

    \I__12526\ : CascadeMux
    port map (
            O => \N__53869\,
            I => \N__53547\
        );

    \I__12525\ : InMux
    port map (
            O => \N__53866\,
            I => \N__53536\
        );

    \I__12524\ : InMux
    port map (
            O => \N__53865\,
            I => \N__53536\
        );

    \I__12523\ : InMux
    port map (
            O => \N__53862\,
            I => \N__53536\
        );

    \I__12522\ : InMux
    port map (
            O => \N__53861\,
            I => \N__53536\
        );

    \I__12521\ : InMux
    port map (
            O => \N__53860\,
            I => \N__53536\
        );

    \I__12520\ : InMux
    port map (
            O => \N__53859\,
            I => \N__53529\
        );

    \I__12519\ : InMux
    port map (
            O => \N__53858\,
            I => \N__53529\
        );

    \I__12518\ : InMux
    port map (
            O => \N__53855\,
            I => \N__53529\
        );

    \I__12517\ : LocalMux
    port map (
            O => \N__53852\,
            I => \N__53524\
        );

    \I__12516\ : LocalMux
    port map (
            O => \N__53845\,
            I => \N__53524\
        );

    \I__12515\ : InMux
    port map (
            O => \N__53842\,
            I => \N__53514\
        );

    \I__12514\ : InMux
    port map (
            O => \N__53841\,
            I => \N__53514\
        );

    \I__12513\ : InMux
    port map (
            O => \N__53840\,
            I => \N__53514\
        );

    \I__12512\ : InMux
    port map (
            O => \N__53839\,
            I => \N__53514\
        );

    \I__12511\ : CascadeMux
    port map (
            O => \N__53838\,
            I => \N__53511\
        );

    \I__12510\ : CascadeMux
    port map (
            O => \N__53837\,
            I => \N__53507\
        );

    \I__12509\ : CascadeMux
    port map (
            O => \N__53836\,
            I => \N__53504\
        );

    \I__12508\ : CascadeMux
    port map (
            O => \N__53835\,
            I => \N__53501\
        );

    \I__12507\ : CascadeMux
    port map (
            O => \N__53834\,
            I => \N__53497\
        );

    \I__12506\ : CascadeMux
    port map (
            O => \N__53833\,
            I => \N__53493\
        );

    \I__12505\ : CascadeMux
    port map (
            O => \N__53832\,
            I => \N__53490\
        );

    \I__12504\ : CascadeMux
    port map (
            O => \N__53831\,
            I => \N__53486\
        );

    \I__12503\ : InMux
    port map (
            O => \N__53830\,
            I => \N__53479\
        );

    \I__12502\ : InMux
    port map (
            O => \N__53829\,
            I => \N__53472\
        );

    \I__12501\ : InMux
    port map (
            O => \N__53828\,
            I => \N__53472\
        );

    \I__12500\ : InMux
    port map (
            O => \N__53827\,
            I => \N__53472\
        );

    \I__12499\ : Span4Mux_v
    port map (
            O => \N__53822\,
            I => \N__53461\
        );

    \I__12498\ : Span4Mux_v
    port map (
            O => \N__53811\,
            I => \N__53461\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__53808\,
            I => \N__53461\
        );

    \I__12496\ : LocalMux
    port map (
            O => \N__53805\,
            I => \N__53461\
        );

    \I__12495\ : LocalMux
    port map (
            O => \N__53796\,
            I => \N__53461\
        );

    \I__12494\ : LocalMux
    port map (
            O => \N__53793\,
            I => \N__53458\
        );

    \I__12493\ : InMux
    port map (
            O => \N__53792\,
            I => \N__53451\
        );

    \I__12492\ : InMux
    port map (
            O => \N__53791\,
            I => \N__53451\
        );

    \I__12491\ : InMux
    port map (
            O => \N__53790\,
            I => \N__53451\
        );

    \I__12490\ : InMux
    port map (
            O => \N__53789\,
            I => \N__53444\
        );

    \I__12489\ : InMux
    port map (
            O => \N__53786\,
            I => \N__53444\
        );

    \I__12488\ : InMux
    port map (
            O => \N__53783\,
            I => \N__53444\
        );

    \I__12487\ : InMux
    port map (
            O => \N__53780\,
            I => \N__53437\
        );

    \I__12486\ : InMux
    port map (
            O => \N__53777\,
            I => \N__53437\
        );

    \I__12485\ : InMux
    port map (
            O => \N__53774\,
            I => \N__53437\
        );

    \I__12484\ : InMux
    port map (
            O => \N__53773\,
            I => \N__53426\
        );

    \I__12483\ : InMux
    port map (
            O => \N__53770\,
            I => \N__53426\
        );

    \I__12482\ : InMux
    port map (
            O => \N__53769\,
            I => \N__53426\
        );

    \I__12481\ : InMux
    port map (
            O => \N__53768\,
            I => \N__53426\
        );

    \I__12480\ : InMux
    port map (
            O => \N__53767\,
            I => \N__53426\
        );

    \I__12479\ : InMux
    port map (
            O => \N__53766\,
            I => \N__53419\
        );

    \I__12478\ : InMux
    port map (
            O => \N__53765\,
            I => \N__53419\
        );

    \I__12477\ : InMux
    port map (
            O => \N__53764\,
            I => \N__53419\
        );

    \I__12476\ : LocalMux
    port map (
            O => \N__53755\,
            I => \N__53408\
        );

    \I__12475\ : Span4Mux_h
    port map (
            O => \N__53742\,
            I => \N__53408\
        );

    \I__12474\ : LocalMux
    port map (
            O => \N__53737\,
            I => \N__53408\
        );

    \I__12473\ : InMux
    port map (
            O => \N__53736\,
            I => \N__53405\
        );

    \I__12472\ : Span4Mux_v
    port map (
            O => \N__53719\,
            I => \N__53400\
        );

    \I__12471\ : Span4Mux_h
    port map (
            O => \N__53714\,
            I => \N__53400\
        );

    \I__12470\ : Span4Mux_h
    port map (
            O => \N__53711\,
            I => \N__53395\
        );

    \I__12469\ : LocalMux
    port map (
            O => \N__53702\,
            I => \N__53395\
        );

    \I__12468\ : Span4Mux_h
    port map (
            O => \N__53697\,
            I => \N__53388\
        );

    \I__12467\ : Span4Mux_v
    port map (
            O => \N__53690\,
            I => \N__53388\
        );

    \I__12466\ : Span4Mux_h
    port map (
            O => \N__53687\,
            I => \N__53388\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__53682\,
            I => \N__53383\
        );

    \I__12464\ : LocalMux
    port map (
            O => \N__53677\,
            I => \N__53383\
        );

    \I__12463\ : InMux
    port map (
            O => \N__53676\,
            I => \N__53374\
        );

    \I__12462\ : InMux
    port map (
            O => \N__53673\,
            I => \N__53374\
        );

    \I__12461\ : InMux
    port map (
            O => \N__53672\,
            I => \N__53374\
        );

    \I__12460\ : InMux
    port map (
            O => \N__53669\,
            I => \N__53374\
        );

    \I__12459\ : CascadeMux
    port map (
            O => \N__53668\,
            I => \N__53370\
        );

    \I__12458\ : CascadeMux
    port map (
            O => \N__53667\,
            I => \N__53367\
        );

    \I__12457\ : CascadeMux
    port map (
            O => \N__53666\,
            I => \N__53363\
        );

    \I__12456\ : CascadeMux
    port map (
            O => \N__53665\,
            I => \N__53353\
        );

    \I__12455\ : CascadeMux
    port map (
            O => \N__53664\,
            I => \N__53344\
        );

    \I__12454\ : CascadeMux
    port map (
            O => \N__53663\,
            I => \N__53341\
        );

    \I__12453\ : CascadeMux
    port map (
            O => \N__53662\,
            I => \N__53337\
        );

    \I__12452\ : Span4Mux_v
    port map (
            O => \N__53659\,
            I => \N__53330\
        );

    \I__12451\ : Span4Mux_h
    port map (
            O => \N__53654\,
            I => \N__53330\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__53647\,
            I => \N__53330\
        );

    \I__12449\ : Span4Mux_v
    port map (
            O => \N__53630\,
            I => \N__53325\
        );

    \I__12448\ : Span4Mux_v
    port map (
            O => \N__53625\,
            I => \N__53325\
        );

    \I__12447\ : InMux
    port map (
            O => \N__53622\,
            I => \N__53318\
        );

    \I__12446\ : InMux
    port map (
            O => \N__53621\,
            I => \N__53318\
        );

    \I__12445\ : InMux
    port map (
            O => \N__53620\,
            I => \N__53318\
        );

    \I__12444\ : InMux
    port map (
            O => \N__53617\,
            I => \N__53307\
        );

    \I__12443\ : InMux
    port map (
            O => \N__53616\,
            I => \N__53307\
        );

    \I__12442\ : InMux
    port map (
            O => \N__53615\,
            I => \N__53307\
        );

    \I__12441\ : InMux
    port map (
            O => \N__53612\,
            I => \N__53307\
        );

    \I__12440\ : InMux
    port map (
            O => \N__53611\,
            I => \N__53307\
        );

    \I__12439\ : Span4Mux_h
    port map (
            O => \N__53608\,
            I => \N__53296\
        );

    \I__12438\ : Span4Mux_v
    port map (
            O => \N__53593\,
            I => \N__53296\
        );

    \I__12437\ : Span4Mux_h
    port map (
            O => \N__53584\,
            I => \N__53296\
        );

    \I__12436\ : LocalMux
    port map (
            O => \N__53581\,
            I => \N__53296\
        );

    \I__12435\ : LocalMux
    port map (
            O => \N__53570\,
            I => \N__53296\
        );

    \I__12434\ : InMux
    port map (
            O => \N__53569\,
            I => \N__53293\
        );

    \I__12433\ : InMux
    port map (
            O => \N__53566\,
            I => \N__53284\
        );

    \I__12432\ : InMux
    port map (
            O => \N__53565\,
            I => \N__53284\
        );

    \I__12431\ : InMux
    port map (
            O => \N__53564\,
            I => \N__53284\
        );

    \I__12430\ : InMux
    port map (
            O => \N__53563\,
            I => \N__53284\
        );

    \I__12429\ : InMux
    port map (
            O => \N__53562\,
            I => \N__53277\
        );

    \I__12428\ : InMux
    port map (
            O => \N__53561\,
            I => \N__53277\
        );

    \I__12427\ : InMux
    port map (
            O => \N__53560\,
            I => \N__53277\
        );

    \I__12426\ : Span4Mux_v
    port map (
            O => \N__53557\,
            I => \N__53274\
        );

    \I__12425\ : InMux
    port map (
            O => \N__53554\,
            I => \N__53265\
        );

    \I__12424\ : InMux
    port map (
            O => \N__53551\,
            I => \N__53265\
        );

    \I__12423\ : InMux
    port map (
            O => \N__53550\,
            I => \N__53265\
        );

    \I__12422\ : InMux
    port map (
            O => \N__53547\,
            I => \N__53265\
        );

    \I__12421\ : LocalMux
    port map (
            O => \N__53536\,
            I => \N__53258\
        );

    \I__12420\ : LocalMux
    port map (
            O => \N__53529\,
            I => \N__53258\
        );

    \I__12419\ : Span4Mux_v
    port map (
            O => \N__53524\,
            I => \N__53258\
        );

    \I__12418\ : InMux
    port map (
            O => \N__53523\,
            I => \N__53255\
        );

    \I__12417\ : LocalMux
    port map (
            O => \N__53514\,
            I => \N__53252\
        );

    \I__12416\ : InMux
    port map (
            O => \N__53511\,
            I => \N__53243\
        );

    \I__12415\ : InMux
    port map (
            O => \N__53510\,
            I => \N__53243\
        );

    \I__12414\ : InMux
    port map (
            O => \N__53507\,
            I => \N__53243\
        );

    \I__12413\ : InMux
    port map (
            O => \N__53504\,
            I => \N__53243\
        );

    \I__12412\ : InMux
    port map (
            O => \N__53501\,
            I => \N__53232\
        );

    \I__12411\ : InMux
    port map (
            O => \N__53500\,
            I => \N__53232\
        );

    \I__12410\ : InMux
    port map (
            O => \N__53497\,
            I => \N__53232\
        );

    \I__12409\ : InMux
    port map (
            O => \N__53496\,
            I => \N__53232\
        );

    \I__12408\ : InMux
    port map (
            O => \N__53493\,
            I => \N__53232\
        );

    \I__12407\ : InMux
    port map (
            O => \N__53490\,
            I => \N__53225\
        );

    \I__12406\ : InMux
    port map (
            O => \N__53489\,
            I => \N__53225\
        );

    \I__12405\ : InMux
    port map (
            O => \N__53486\,
            I => \N__53225\
        );

    \I__12404\ : InMux
    port map (
            O => \N__53485\,
            I => \N__53222\
        );

    \I__12403\ : InMux
    port map (
            O => \N__53484\,
            I => \N__53215\
        );

    \I__12402\ : InMux
    port map (
            O => \N__53483\,
            I => \N__53215\
        );

    \I__12401\ : InMux
    port map (
            O => \N__53482\,
            I => \N__53215\
        );

    \I__12400\ : LocalMux
    port map (
            O => \N__53479\,
            I => \N__53210\
        );

    \I__12399\ : LocalMux
    port map (
            O => \N__53472\,
            I => \N__53210\
        );

    \I__12398\ : Span4Mux_v
    port map (
            O => \N__53461\,
            I => \N__53195\
        );

    \I__12397\ : Span4Mux_s2_h
    port map (
            O => \N__53458\,
            I => \N__53195\
        );

    \I__12396\ : LocalMux
    port map (
            O => \N__53451\,
            I => \N__53195\
        );

    \I__12395\ : LocalMux
    port map (
            O => \N__53444\,
            I => \N__53195\
        );

    \I__12394\ : LocalMux
    port map (
            O => \N__53437\,
            I => \N__53195\
        );

    \I__12393\ : LocalMux
    port map (
            O => \N__53426\,
            I => \N__53195\
        );

    \I__12392\ : LocalMux
    port map (
            O => \N__53419\,
            I => \N__53195\
        );

    \I__12391\ : InMux
    port map (
            O => \N__53418\,
            I => \N__53192\
        );

    \I__12390\ : InMux
    port map (
            O => \N__53417\,
            I => \N__53185\
        );

    \I__12389\ : InMux
    port map (
            O => \N__53416\,
            I => \N__53185\
        );

    \I__12388\ : InMux
    port map (
            O => \N__53415\,
            I => \N__53185\
        );

    \I__12387\ : Span4Mux_v
    port map (
            O => \N__53408\,
            I => \N__53180\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__53405\,
            I => \N__53180\
        );

    \I__12385\ : Span4Mux_h
    port map (
            O => \N__53400\,
            I => \N__53172\
        );

    \I__12384\ : Span4Mux_v
    port map (
            O => \N__53395\,
            I => \N__53172\
        );

    \I__12383\ : Span4Mux_v
    port map (
            O => \N__53388\,
            I => \N__53165\
        );

    \I__12382\ : Span4Mux_h
    port map (
            O => \N__53383\,
            I => \N__53165\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__53374\,
            I => \N__53165\
        );

    \I__12380\ : InMux
    port map (
            O => \N__53373\,
            I => \N__53154\
        );

    \I__12379\ : InMux
    port map (
            O => \N__53370\,
            I => \N__53154\
        );

    \I__12378\ : InMux
    port map (
            O => \N__53367\,
            I => \N__53154\
        );

    \I__12377\ : InMux
    port map (
            O => \N__53366\,
            I => \N__53154\
        );

    \I__12376\ : InMux
    port map (
            O => \N__53363\,
            I => \N__53154\
        );

    \I__12375\ : InMux
    port map (
            O => \N__53362\,
            I => \N__53151\
        );

    \I__12374\ : InMux
    port map (
            O => \N__53361\,
            I => \N__53144\
        );

    \I__12373\ : InMux
    port map (
            O => \N__53360\,
            I => \N__53144\
        );

    \I__12372\ : InMux
    port map (
            O => \N__53359\,
            I => \N__53144\
        );

    \I__12371\ : InMux
    port map (
            O => \N__53358\,
            I => \N__53137\
        );

    \I__12370\ : InMux
    port map (
            O => \N__53357\,
            I => \N__53137\
        );

    \I__12369\ : InMux
    port map (
            O => \N__53356\,
            I => \N__53137\
        );

    \I__12368\ : InMux
    port map (
            O => \N__53353\,
            I => \N__53126\
        );

    \I__12367\ : InMux
    port map (
            O => \N__53352\,
            I => \N__53126\
        );

    \I__12366\ : InMux
    port map (
            O => \N__53351\,
            I => \N__53126\
        );

    \I__12365\ : InMux
    port map (
            O => \N__53350\,
            I => \N__53126\
        );

    \I__12364\ : InMux
    port map (
            O => \N__53349\,
            I => \N__53126\
        );

    \I__12363\ : CascadeMux
    port map (
            O => \N__53348\,
            I => \N__53121\
        );

    \I__12362\ : CascadeMux
    port map (
            O => \N__53347\,
            I => \N__53118\
        );

    \I__12361\ : InMux
    port map (
            O => \N__53344\,
            I => \N__53109\
        );

    \I__12360\ : InMux
    port map (
            O => \N__53341\,
            I => \N__53109\
        );

    \I__12359\ : InMux
    port map (
            O => \N__53340\,
            I => \N__53109\
        );

    \I__12358\ : InMux
    port map (
            O => \N__53337\,
            I => \N__53109\
        );

    \I__12357\ : Span4Mux_v
    port map (
            O => \N__53330\,
            I => \N__53105\
        );

    \I__12356\ : Span4Mux_v
    port map (
            O => \N__53325\,
            I => \N__53098\
        );

    \I__12355\ : LocalMux
    port map (
            O => \N__53318\,
            I => \N__53098\
        );

    \I__12354\ : LocalMux
    port map (
            O => \N__53307\,
            I => \N__53098\
        );

    \I__12353\ : Span4Mux_v
    port map (
            O => \N__53296\,
            I => \N__53093\
        );

    \I__12352\ : LocalMux
    port map (
            O => \N__53293\,
            I => \N__53093\
        );

    \I__12351\ : LocalMux
    port map (
            O => \N__53284\,
            I => \N__53088\
        );

    \I__12350\ : LocalMux
    port map (
            O => \N__53277\,
            I => \N__53088\
        );

    \I__12349\ : Span4Mux_h
    port map (
            O => \N__53274\,
            I => \N__53083\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__53265\,
            I => \N__53083\
        );

    \I__12347\ : Span4Mux_h
    port map (
            O => \N__53258\,
            I => \N__53066\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__53255\,
            I => \N__53066\
        );

    \I__12345\ : Span4Mux_h
    port map (
            O => \N__53252\,
            I => \N__53066\
        );

    \I__12344\ : LocalMux
    port map (
            O => \N__53243\,
            I => \N__53066\
        );

    \I__12343\ : LocalMux
    port map (
            O => \N__53232\,
            I => \N__53066\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__53225\,
            I => \N__53066\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__53222\,
            I => \N__53066\
        );

    \I__12340\ : LocalMux
    port map (
            O => \N__53215\,
            I => \N__53066\
        );

    \I__12339\ : Span4Mux_s2_h
    port map (
            O => \N__53210\,
            I => \N__53054\
        );

    \I__12338\ : Span4Mux_v
    port map (
            O => \N__53195\,
            I => \N__53054\
        );

    \I__12337\ : LocalMux
    port map (
            O => \N__53192\,
            I => \N__53054\
        );

    \I__12336\ : LocalMux
    port map (
            O => \N__53185\,
            I => \N__53054\
        );

    \I__12335\ : Span4Mux_v
    port map (
            O => \N__53180\,
            I => \N__53051\
        );

    \I__12334\ : InMux
    port map (
            O => \N__53179\,
            I => \N__53044\
        );

    \I__12333\ : InMux
    port map (
            O => \N__53178\,
            I => \N__53044\
        );

    \I__12332\ : InMux
    port map (
            O => \N__53177\,
            I => \N__53044\
        );

    \I__12331\ : Span4Mux_h
    port map (
            O => \N__53172\,
            I => \N__53029\
        );

    \I__12330\ : Span4Mux_v
    port map (
            O => \N__53165\,
            I => \N__53029\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__53154\,
            I => \N__53029\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__53151\,
            I => \N__53029\
        );

    \I__12327\ : LocalMux
    port map (
            O => \N__53144\,
            I => \N__53029\
        );

    \I__12326\ : LocalMux
    port map (
            O => \N__53137\,
            I => \N__53029\
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__53126\,
            I => \N__53029\
        );

    \I__12324\ : InMux
    port map (
            O => \N__53125\,
            I => \N__53020\
        );

    \I__12323\ : InMux
    port map (
            O => \N__53124\,
            I => \N__53020\
        );

    \I__12322\ : InMux
    port map (
            O => \N__53121\,
            I => \N__53020\
        );

    \I__12321\ : InMux
    port map (
            O => \N__53118\,
            I => \N__53020\
        );

    \I__12320\ : LocalMux
    port map (
            O => \N__53109\,
            I => \N__53017\
        );

    \I__12319\ : CascadeMux
    port map (
            O => \N__53108\,
            I => \N__53011\
        );

    \I__12318\ : Span4Mux_v
    port map (
            O => \N__53105\,
            I => \N__53002\
        );

    \I__12317\ : Span4Mux_h
    port map (
            O => \N__53098\,
            I => \N__53002\
        );

    \I__12316\ : Span4Mux_v
    port map (
            O => \N__53093\,
            I => \N__52999\
        );

    \I__12315\ : Span4Mux_v
    port map (
            O => \N__53088\,
            I => \N__52996\
        );

    \I__12314\ : Span4Mux_v
    port map (
            O => \N__53083\,
            I => \N__52991\
        );

    \I__12313\ : Span4Mux_v
    port map (
            O => \N__53066\,
            I => \N__52991\
        );

    \I__12312\ : InMux
    port map (
            O => \N__53065\,
            I => \N__52986\
        );

    \I__12311\ : InMux
    port map (
            O => \N__53064\,
            I => \N__52986\
        );

    \I__12310\ : CascadeMux
    port map (
            O => \N__53063\,
            I => \N__52982\
        );

    \I__12309\ : Span4Mux_h
    port map (
            O => \N__53054\,
            I => \N__52975\
        );

    \I__12308\ : Span4Mux_h
    port map (
            O => \N__53051\,
            I => \N__52975\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__53044\,
            I => \N__52975\
        );

    \I__12306\ : Span4Mux_v
    port map (
            O => \N__53029\,
            I => \N__52968\
        );

    \I__12305\ : LocalMux
    port map (
            O => \N__53020\,
            I => \N__52968\
        );

    \I__12304\ : Span4Mux_h
    port map (
            O => \N__53017\,
            I => \N__52968\
        );

    \I__12303\ : InMux
    port map (
            O => \N__53016\,
            I => \N__52961\
        );

    \I__12302\ : InMux
    port map (
            O => \N__53015\,
            I => \N__52961\
        );

    \I__12301\ : InMux
    port map (
            O => \N__53014\,
            I => \N__52961\
        );

    \I__12300\ : InMux
    port map (
            O => \N__53011\,
            I => \N__52950\
        );

    \I__12299\ : InMux
    port map (
            O => \N__53010\,
            I => \N__52950\
        );

    \I__12298\ : InMux
    port map (
            O => \N__53009\,
            I => \N__52950\
        );

    \I__12297\ : InMux
    port map (
            O => \N__53008\,
            I => \N__52950\
        );

    \I__12296\ : InMux
    port map (
            O => \N__53007\,
            I => \N__52950\
        );

    \I__12295\ : Span4Mux_v
    port map (
            O => \N__53002\,
            I => \N__52939\
        );

    \I__12294\ : Span4Mux_h
    port map (
            O => \N__52999\,
            I => \N__52939\
        );

    \I__12293\ : Span4Mux_h
    port map (
            O => \N__52996\,
            I => \N__52939\
        );

    \I__12292\ : Span4Mux_v
    port map (
            O => \N__52991\,
            I => \N__52939\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__52986\,
            I => \N__52939\
        );

    \I__12290\ : InMux
    port map (
            O => \N__52985\,
            I => \N__52934\
        );

    \I__12289\ : InMux
    port map (
            O => \N__52982\,
            I => \N__52934\
        );

    \I__12288\ : Odrv4
    port map (
            O => \N__52975\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12287\ : Odrv4
    port map (
            O => \N__52968\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__52961\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__52950\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12284\ : Odrv4
    port map (
            O => \N__52939\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12283\ : LocalMux
    port map (
            O => \N__52934\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12282\ : InMux
    port map (
            O => \N__52921\,
            I => n12685
        );

    \I__12281\ : InMux
    port map (
            O => \N__52918\,
            I => \N__52914\
        );

    \I__12280\ : InMux
    port map (
            O => \N__52917\,
            I => \N__52910\
        );

    \I__12279\ : LocalMux
    port map (
            O => \N__52914\,
            I => \N__52907\
        );

    \I__12278\ : InMux
    port map (
            O => \N__52913\,
            I => \N__52904\
        );

    \I__12277\ : LocalMux
    port map (
            O => \N__52910\,
            I => encoder0_position_target_23
        );

    \I__12276\ : Odrv4
    port map (
            O => \N__52907\,
            I => encoder0_position_target_23
        );

    \I__12275\ : LocalMux
    port map (
            O => \N__52904\,
            I => encoder0_position_target_23
        );

    \I__12274\ : CEMux
    port map (
            O => \N__52897\,
            I => \N__52893\
        );

    \I__12273\ : CEMux
    port map (
            O => \N__52896\,
            I => \N__52890\
        );

    \I__12272\ : LocalMux
    port map (
            O => \N__52893\,
            I => \N__52887\
        );

    \I__12271\ : LocalMux
    port map (
            O => \N__52890\,
            I => \N__52884\
        );

    \I__12270\ : Span4Mux_v
    port map (
            O => \N__52887\,
            I => \N__52876\
        );

    \I__12269\ : Span4Mux_h
    port map (
            O => \N__52884\,
            I => \N__52876\
        );

    \I__12268\ : SRMux
    port map (
            O => \N__52883\,
            I => \N__52873\
        );

    \I__12267\ : SRMux
    port map (
            O => \N__52882\,
            I => \N__52870\
        );

    \I__12266\ : CEMux
    port map (
            O => \N__52881\,
            I => \N__52866\
        );

    \I__12265\ : Span4Mux_v
    port map (
            O => \N__52876\,
            I => \N__52860\
        );

    \I__12264\ : LocalMux
    port map (
            O => \N__52873\,
            I => \N__52860\
        );

    \I__12263\ : LocalMux
    port map (
            O => \N__52870\,
            I => \N__52857\
        );

    \I__12262\ : SRMux
    port map (
            O => \N__52869\,
            I => \N__52854\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__52866\,
            I => \N__52851\
        );

    \I__12260\ : InMux
    port map (
            O => \N__52865\,
            I => \N__52848\
        );

    \I__12259\ : Span4Mux_v
    port map (
            O => \N__52860\,
            I => \N__52845\
        );

    \I__12258\ : Span4Mux_h
    port map (
            O => \N__52857\,
            I => \N__52840\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__52854\,
            I => \N__52840\
        );

    \I__12256\ : Span12Mux_h
    port map (
            O => \N__52851\,
            I => \N__52835\
        );

    \I__12255\ : LocalMux
    port map (
            O => \N__52848\,
            I => \N__52835\
        );

    \I__12254\ : Odrv4
    port map (
            O => \N__52845\,
            I => n4856
        );

    \I__12253\ : Odrv4
    port map (
            O => \N__52840\,
            I => n4856
        );

    \I__12252\ : Odrv12
    port map (
            O => \N__52835\,
            I => n4856
        );

    \I__12251\ : SRMux
    port map (
            O => \N__52828\,
            I => \N__52824\
        );

    \I__12250\ : SRMux
    port map (
            O => \N__52827\,
            I => \N__52820\
        );

    \I__12249\ : LocalMux
    port map (
            O => \N__52824\,
            I => \N__52817\
        );

    \I__12248\ : SRMux
    port map (
            O => \N__52823\,
            I => \N__52814\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__52820\,
            I => \N__52811\
        );

    \I__12246\ : Span4Mux_v
    port map (
            O => \N__52817\,
            I => \N__52806\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__52814\,
            I => \N__52806\
        );

    \I__12244\ : Odrv4
    port map (
            O => \N__52811\,
            I => n4890
        );

    \I__12243\ : Odrv4
    port map (
            O => \N__52806\,
            I => n4890
        );

    \I__12242\ : InMux
    port map (
            O => \N__52801\,
            I => \N__52798\
        );

    \I__12241\ : LocalMux
    port map (
            O => \N__52798\,
            I => \N__52795\
        );

    \I__12240\ : Odrv12
    port map (
            O => \N__52795\,
            I => \pwm_setpoint_23_N_171_9\
        );

    \I__12239\ : InMux
    port map (
            O => \N__52792\,
            I => \N__52789\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__52789\,
            I => \N__52785\
        );

    \I__12237\ : InMux
    port map (
            O => \N__52788\,
            I => \N__52782\
        );

    \I__12236\ : Span4Mux_h
    port map (
            O => \N__52785\,
            I => \N__52779\
        );

    \I__12235\ : LocalMux
    port map (
            O => \N__52782\,
            I => \N__52776\
        );

    \I__12234\ : Odrv4
    port map (
            O => \N__52779\,
            I => duty_9
        );

    \I__12233\ : Odrv12
    port map (
            O => \N__52776\,
            I => duty_9
        );

    \I__12232\ : InMux
    port map (
            O => \N__52771\,
            I => \N__52767\
        );

    \I__12231\ : InMux
    port map (
            O => \N__52770\,
            I => \N__52764\
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__52767\,
            I => \N__52760\
        );

    \I__12229\ : LocalMux
    port map (
            O => \N__52764\,
            I => \N__52757\
        );

    \I__12228\ : InMux
    port map (
            O => \N__52763\,
            I => \N__52754\
        );

    \I__12227\ : Span4Mux_h
    port map (
            O => \N__52760\,
            I => \N__52751\
        );

    \I__12226\ : Span4Mux_s3_v
    port map (
            O => \N__52757\,
            I => \N__52748\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__52754\,
            I => \N__52745\
        );

    \I__12224\ : Span4Mux_h
    port map (
            O => \N__52751\,
            I => \N__52742\
        );

    \I__12223\ : Sp12to4
    port map (
            O => \N__52748\,
            I => \N__52737\
        );

    \I__12222\ : Span12Mux_s3_v
    port map (
            O => \N__52745\,
            I => \N__52737\
        );

    \I__12221\ : Odrv4
    port map (
            O => \N__52742\,
            I => pwm_setpoint_9
        );

    \I__12220\ : Odrv12
    port map (
            O => \N__52737\,
            I => pwm_setpoint_9
        );

    \I__12219\ : InMux
    port map (
            O => \N__52732\,
            I => \N__52728\
        );

    \I__12218\ : InMux
    port map (
            O => \N__52731\,
            I => \N__52725\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__52728\,
            I => \N__52722\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__52725\,
            I => \N__52719\
        );

    \I__12215\ : Span4Mux_h
    port map (
            O => \N__52722\,
            I => \N__52714\
        );

    \I__12214\ : Span4Mux_h
    port map (
            O => \N__52719\,
            I => \N__52714\
        );

    \I__12213\ : Odrv4
    port map (
            O => \N__52714\,
            I => duty_8
        );

    \I__12212\ : InMux
    port map (
            O => \N__52711\,
            I => \N__52708\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__52708\,
            I => \N__52705\
        );

    \I__12210\ : Odrv4
    port map (
            O => \N__52705\,
            I => n17_adj_583
        );

    \I__12209\ : CascadeMux
    port map (
            O => \N__52702\,
            I => \N__52698\
        );

    \I__12208\ : InMux
    port map (
            O => \N__52701\,
            I => \N__52695\
        );

    \I__12207\ : InMux
    port map (
            O => \N__52698\,
            I => \N__52691\
        );

    \I__12206\ : LocalMux
    port map (
            O => \N__52695\,
            I => \N__52688\
        );

    \I__12205\ : InMux
    port map (
            O => \N__52694\,
            I => \N__52685\
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__52691\,
            I => encoder0_position_target_10
        );

    \I__12203\ : Odrv4
    port map (
            O => \N__52688\,
            I => encoder0_position_target_10
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__52685\,
            I => encoder0_position_target_10
        );

    \I__12201\ : InMux
    port map (
            O => \N__52678\,
            I => n12672
        );

    \I__12200\ : InMux
    port map (
            O => \N__52675\,
            I => \N__52671\
        );

    \I__12199\ : InMux
    port map (
            O => \N__52674\,
            I => \N__52667\
        );

    \I__12198\ : LocalMux
    port map (
            O => \N__52671\,
            I => \N__52664\
        );

    \I__12197\ : InMux
    port map (
            O => \N__52670\,
            I => \N__52661\
        );

    \I__12196\ : LocalMux
    port map (
            O => \N__52667\,
            I => encoder0_position_target_11
        );

    \I__12195\ : Odrv4
    port map (
            O => \N__52664\,
            I => encoder0_position_target_11
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__52661\,
            I => encoder0_position_target_11
        );

    \I__12193\ : InMux
    port map (
            O => \N__52654\,
            I => n12673
        );

    \I__12192\ : CascadeMux
    port map (
            O => \N__52651\,
            I => \N__52647\
        );

    \I__12191\ : CascadeMux
    port map (
            O => \N__52650\,
            I => \N__52644\
        );

    \I__12190\ : InMux
    port map (
            O => \N__52647\,
            I => \N__52641\
        );

    \I__12189\ : InMux
    port map (
            O => \N__52644\,
            I => \N__52637\
        );

    \I__12188\ : LocalMux
    port map (
            O => \N__52641\,
            I => \N__52634\
        );

    \I__12187\ : InMux
    port map (
            O => \N__52640\,
            I => \N__52631\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__52637\,
            I => encoder0_position_target_12
        );

    \I__12185\ : Odrv4
    port map (
            O => \N__52634\,
            I => encoder0_position_target_12
        );

    \I__12184\ : LocalMux
    port map (
            O => \N__52631\,
            I => encoder0_position_target_12
        );

    \I__12183\ : InMux
    port map (
            O => \N__52624\,
            I => n12674
        );

    \I__12182\ : CascadeMux
    port map (
            O => \N__52621\,
            I => \N__52618\
        );

    \I__12181\ : InMux
    port map (
            O => \N__52618\,
            I => \N__52613\
        );

    \I__12180\ : InMux
    port map (
            O => \N__52617\,
            I => \N__52610\
        );

    \I__12179\ : InMux
    port map (
            O => \N__52616\,
            I => \N__52607\
        );

    \I__12178\ : LocalMux
    port map (
            O => \N__52613\,
            I => \N__52604\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__52610\,
            I => \N__52601\
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__52607\,
            I => encoder0_position_target_13
        );

    \I__12175\ : Odrv4
    port map (
            O => \N__52604\,
            I => encoder0_position_target_13
        );

    \I__12174\ : Odrv4
    port map (
            O => \N__52601\,
            I => encoder0_position_target_13
        );

    \I__12173\ : InMux
    port map (
            O => \N__52594\,
            I => n12675
        );

    \I__12172\ : InMux
    port map (
            O => \N__52591\,
            I => \N__52587\
        );

    \I__12171\ : CascadeMux
    port map (
            O => \N__52590\,
            I => \N__52583\
        );

    \I__12170\ : LocalMux
    port map (
            O => \N__52587\,
            I => \N__52580\
        );

    \I__12169\ : CascadeMux
    port map (
            O => \N__52586\,
            I => \N__52577\
        );

    \I__12168\ : InMux
    port map (
            O => \N__52583\,
            I => \N__52574\
        );

    \I__12167\ : Span4Mux_h
    port map (
            O => \N__52580\,
            I => \N__52571\
        );

    \I__12166\ : InMux
    port map (
            O => \N__52577\,
            I => \N__52568\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__52574\,
            I => encoder0_position_target_14
        );

    \I__12164\ : Odrv4
    port map (
            O => \N__52571\,
            I => encoder0_position_target_14
        );

    \I__12163\ : LocalMux
    port map (
            O => \N__52568\,
            I => encoder0_position_target_14
        );

    \I__12162\ : InMux
    port map (
            O => \N__52561\,
            I => n12676
        );

    \I__12161\ : CascadeMux
    port map (
            O => \N__52558\,
            I => \N__52555\
        );

    \I__12160\ : InMux
    port map (
            O => \N__52555\,
            I => \N__52551\
        );

    \I__12159\ : InMux
    port map (
            O => \N__52554\,
            I => \N__52547\
        );

    \I__12158\ : LocalMux
    port map (
            O => \N__52551\,
            I => \N__52544\
        );

    \I__12157\ : InMux
    port map (
            O => \N__52550\,
            I => \N__52541\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__52547\,
            I => encoder0_position_target_15
        );

    \I__12155\ : Odrv12
    port map (
            O => \N__52544\,
            I => encoder0_position_target_15
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__52541\,
            I => encoder0_position_target_15
        );

    \I__12153\ : InMux
    port map (
            O => \N__52534\,
            I => n12677
        );

    \I__12152\ : InMux
    port map (
            O => \N__52531\,
            I => \N__52527\
        );

    \I__12151\ : InMux
    port map (
            O => \N__52530\,
            I => \N__52523\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__52527\,
            I => \N__52520\
        );

    \I__12149\ : InMux
    port map (
            O => \N__52526\,
            I => \N__52517\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__52523\,
            I => encoder0_position_target_16
        );

    \I__12147\ : Odrv4
    port map (
            O => \N__52520\,
            I => encoder0_position_target_16
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__52517\,
            I => encoder0_position_target_16
        );

    \I__12145\ : InMux
    port map (
            O => \N__52510\,
            I => \bfn_16_28_0_\
        );

    \I__12144\ : CascadeMux
    port map (
            O => \N__52507\,
            I => \N__52504\
        );

    \I__12143\ : InMux
    port map (
            O => \N__52504\,
            I => \N__52500\
        );

    \I__12142\ : CascadeMux
    port map (
            O => \N__52503\,
            I => \N__52497\
        );

    \I__12141\ : LocalMux
    port map (
            O => \N__52500\,
            I => \N__52494\
        );

    \I__12140\ : InMux
    port map (
            O => \N__52497\,
            I => \N__52490\
        );

    \I__12139\ : Span4Mux_h
    port map (
            O => \N__52494\,
            I => \N__52487\
        );

    \I__12138\ : InMux
    port map (
            O => \N__52493\,
            I => \N__52484\
        );

    \I__12137\ : LocalMux
    port map (
            O => \N__52490\,
            I => encoder0_position_target_17
        );

    \I__12136\ : Odrv4
    port map (
            O => \N__52487\,
            I => encoder0_position_target_17
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__52484\,
            I => encoder0_position_target_17
        );

    \I__12134\ : InMux
    port map (
            O => \N__52477\,
            I => n12679
        );

    \I__12133\ : InMux
    port map (
            O => \N__52474\,
            I => \N__52471\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__52471\,
            I => \N__52467\
        );

    \I__12131\ : InMux
    port map (
            O => \N__52470\,
            I => \N__52463\
        );

    \I__12130\ : Span4Mux_h
    port map (
            O => \N__52467\,
            I => \N__52460\
        );

    \I__12129\ : InMux
    port map (
            O => \N__52466\,
            I => \N__52457\
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__52463\,
            I => encoder0_position_target_1
        );

    \I__12127\ : Odrv4
    port map (
            O => \N__52460\,
            I => encoder0_position_target_1
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__52457\,
            I => encoder0_position_target_1
        );

    \I__12125\ : InMux
    port map (
            O => \N__52450\,
            I => n12663
        );

    \I__12124\ : CascadeMux
    port map (
            O => \N__52447\,
            I => \N__52444\
        );

    \I__12123\ : InMux
    port map (
            O => \N__52444\,
            I => \N__52440\
        );

    \I__12122\ : CascadeMux
    port map (
            O => \N__52443\,
            I => \N__52437\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__52440\,
            I => \N__52434\
        );

    \I__12120\ : InMux
    port map (
            O => \N__52437\,
            I => \N__52430\
        );

    \I__12119\ : Span4Mux_h
    port map (
            O => \N__52434\,
            I => \N__52427\
        );

    \I__12118\ : InMux
    port map (
            O => \N__52433\,
            I => \N__52424\
        );

    \I__12117\ : LocalMux
    port map (
            O => \N__52430\,
            I => encoder0_position_target_2
        );

    \I__12116\ : Odrv4
    port map (
            O => \N__52427\,
            I => encoder0_position_target_2
        );

    \I__12115\ : LocalMux
    port map (
            O => \N__52424\,
            I => encoder0_position_target_2
        );

    \I__12114\ : InMux
    port map (
            O => \N__52417\,
            I => n12664
        );

    \I__12113\ : InMux
    port map (
            O => \N__52414\,
            I => \N__52411\
        );

    \I__12112\ : LocalMux
    port map (
            O => \N__52411\,
            I => \N__52407\
        );

    \I__12111\ : InMux
    port map (
            O => \N__52410\,
            I => \N__52403\
        );

    \I__12110\ : Span4Mux_h
    port map (
            O => \N__52407\,
            I => \N__52400\
        );

    \I__12109\ : InMux
    port map (
            O => \N__52406\,
            I => \N__52397\
        );

    \I__12108\ : LocalMux
    port map (
            O => \N__52403\,
            I => encoder0_position_target_3
        );

    \I__12107\ : Odrv4
    port map (
            O => \N__52400\,
            I => encoder0_position_target_3
        );

    \I__12106\ : LocalMux
    port map (
            O => \N__52397\,
            I => encoder0_position_target_3
        );

    \I__12105\ : InMux
    port map (
            O => \N__52390\,
            I => n12665
        );

    \I__12104\ : InMux
    port map (
            O => \N__52387\,
            I => \N__52383\
        );

    \I__12103\ : CascadeMux
    port map (
            O => \N__52386\,
            I => \N__52380\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__52383\,
            I => \N__52377\
        );

    \I__12101\ : InMux
    port map (
            O => \N__52380\,
            I => \N__52373\
        );

    \I__12100\ : Span4Mux_h
    port map (
            O => \N__52377\,
            I => \N__52370\
        );

    \I__12099\ : InMux
    port map (
            O => \N__52376\,
            I => \N__52367\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__52373\,
            I => encoder0_position_target_4
        );

    \I__12097\ : Odrv4
    port map (
            O => \N__52370\,
            I => encoder0_position_target_4
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__52367\,
            I => encoder0_position_target_4
        );

    \I__12095\ : InMux
    port map (
            O => \N__52360\,
            I => n12666
        );

    \I__12094\ : InMux
    port map (
            O => \N__52357\,
            I => \N__52353\
        );

    \I__12093\ : InMux
    port map (
            O => \N__52356\,
            I => \N__52349\
        );

    \I__12092\ : LocalMux
    port map (
            O => \N__52353\,
            I => \N__52346\
        );

    \I__12091\ : InMux
    port map (
            O => \N__52352\,
            I => \N__52343\
        );

    \I__12090\ : LocalMux
    port map (
            O => \N__52349\,
            I => encoder0_position_target_5
        );

    \I__12089\ : Odrv4
    port map (
            O => \N__52346\,
            I => encoder0_position_target_5
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__52343\,
            I => encoder0_position_target_5
        );

    \I__12087\ : InMux
    port map (
            O => \N__52336\,
            I => n12667
        );

    \I__12086\ : CascadeMux
    port map (
            O => \N__52333\,
            I => \N__52329\
        );

    \I__12085\ : InMux
    port map (
            O => \N__52332\,
            I => \N__52326\
        );

    \I__12084\ : InMux
    port map (
            O => \N__52329\,
            I => \N__52322\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__52326\,
            I => \N__52319\
        );

    \I__12082\ : InMux
    port map (
            O => \N__52325\,
            I => \N__52316\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__52322\,
            I => encoder0_position_target_6
        );

    \I__12080\ : Odrv4
    port map (
            O => \N__52319\,
            I => encoder0_position_target_6
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__52316\,
            I => encoder0_position_target_6
        );

    \I__12078\ : InMux
    port map (
            O => \N__52309\,
            I => n12668
        );

    \I__12077\ : InMux
    port map (
            O => \N__52306\,
            I => \N__52302\
        );

    \I__12076\ : InMux
    port map (
            O => \N__52305\,
            I => \N__52298\
        );

    \I__12075\ : LocalMux
    port map (
            O => \N__52302\,
            I => \N__52295\
        );

    \I__12074\ : InMux
    port map (
            O => \N__52301\,
            I => \N__52292\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__52298\,
            I => encoder0_position_target_7
        );

    \I__12072\ : Odrv4
    port map (
            O => \N__52295\,
            I => encoder0_position_target_7
        );

    \I__12071\ : LocalMux
    port map (
            O => \N__52292\,
            I => encoder0_position_target_7
        );

    \I__12070\ : InMux
    port map (
            O => \N__52285\,
            I => n12669
        );

    \I__12069\ : CascadeMux
    port map (
            O => \N__52282\,
            I => \N__52277\
        );

    \I__12068\ : InMux
    port map (
            O => \N__52281\,
            I => \N__52274\
        );

    \I__12067\ : CascadeMux
    port map (
            O => \N__52280\,
            I => \N__52271\
        );

    \I__12066\ : InMux
    port map (
            O => \N__52277\,
            I => \N__52268\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__52274\,
            I => \N__52265\
        );

    \I__12064\ : InMux
    port map (
            O => \N__52271\,
            I => \N__52262\
        );

    \I__12063\ : LocalMux
    port map (
            O => \N__52268\,
            I => encoder0_position_target_8
        );

    \I__12062\ : Odrv4
    port map (
            O => \N__52265\,
            I => encoder0_position_target_8
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__52262\,
            I => encoder0_position_target_8
        );

    \I__12060\ : InMux
    port map (
            O => \N__52255\,
            I => \bfn_16_27_0_\
        );

    \I__12059\ : InMux
    port map (
            O => \N__52252\,
            I => \N__52249\
        );

    \I__12058\ : LocalMux
    port map (
            O => \N__52249\,
            I => \N__52245\
        );

    \I__12057\ : InMux
    port map (
            O => \N__52248\,
            I => \N__52241\
        );

    \I__12056\ : Span4Mux_h
    port map (
            O => \N__52245\,
            I => \N__52238\
        );

    \I__12055\ : InMux
    port map (
            O => \N__52244\,
            I => \N__52235\
        );

    \I__12054\ : LocalMux
    port map (
            O => \N__52241\,
            I => encoder0_position_target_9
        );

    \I__12053\ : Odrv4
    port map (
            O => \N__52238\,
            I => encoder0_position_target_9
        );

    \I__12052\ : LocalMux
    port map (
            O => \N__52235\,
            I => encoder0_position_target_9
        );

    \I__12051\ : InMux
    port map (
            O => \N__52228\,
            I => n12671
        );

    \I__12050\ : InMux
    port map (
            O => \N__52225\,
            I => \N__52221\
        );

    \I__12049\ : InMux
    port map (
            O => \N__52224\,
            I => \N__52218\
        );

    \I__12048\ : LocalMux
    port map (
            O => \N__52221\,
            I => \N__52215\
        );

    \I__12047\ : LocalMux
    port map (
            O => \N__52218\,
            I => \N__52211\
        );

    \I__12046\ : Span4Mux_v
    port map (
            O => \N__52215\,
            I => \N__52208\
        );

    \I__12045\ : InMux
    port map (
            O => \N__52214\,
            I => \N__52205\
        );

    \I__12044\ : Span4Mux_v
    port map (
            O => \N__52211\,
            I => \N__52202\
        );

    \I__12043\ : Span4Mux_h
    port map (
            O => \N__52208\,
            I => \N__52199\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__52205\,
            I => \N__52196\
        );

    \I__12041\ : Odrv4
    port map (
            O => \N__52202\,
            I => n3111
        );

    \I__12040\ : Odrv4
    port map (
            O => \N__52199\,
            I => n3111
        );

    \I__12039\ : Odrv12
    port map (
            O => \N__52196\,
            I => n3111
        );

    \I__12038\ : CascadeMux
    port map (
            O => \N__52189\,
            I => \N__52186\
        );

    \I__12037\ : InMux
    port map (
            O => \N__52186\,
            I => \N__52183\
        );

    \I__12036\ : LocalMux
    port map (
            O => \N__52183\,
            I => \N__52180\
        );

    \I__12035\ : Odrv12
    port map (
            O => \N__52180\,
            I => n3178
        );

    \I__12034\ : InMux
    port map (
            O => \N__52177\,
            I => n12514
        );

    \I__12033\ : InMux
    port map (
            O => \N__52174\,
            I => \N__52171\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__52171\,
            I => \N__52168\
        );

    \I__12031\ : Span4Mux_v
    port map (
            O => \N__52168\,
            I => \N__52164\
        );

    \I__12030\ : InMux
    port map (
            O => \N__52167\,
            I => \N__52161\
        );

    \I__12029\ : Span4Mux_h
    port map (
            O => \N__52164\,
            I => \N__52158\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__52161\,
            I => n3110
        );

    \I__12027\ : Odrv4
    port map (
            O => \N__52158\,
            I => n3110
        );

    \I__12026\ : InMux
    port map (
            O => \N__52153\,
            I => \N__52150\
        );

    \I__12025\ : LocalMux
    port map (
            O => \N__52150\,
            I => n3177
        );

    \I__12024\ : InMux
    port map (
            O => \N__52147\,
            I => \bfn_16_25_0_\
        );

    \I__12023\ : InMux
    port map (
            O => \N__52144\,
            I => \N__52141\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__52141\,
            I => \N__52137\
        );

    \I__12021\ : InMux
    port map (
            O => \N__52140\,
            I => \N__52134\
        );

    \I__12020\ : Span4Mux_v
    port map (
            O => \N__52137\,
            I => \N__52130\
        );

    \I__12019\ : LocalMux
    port map (
            O => \N__52134\,
            I => \N__52127\
        );

    \I__12018\ : InMux
    port map (
            O => \N__52133\,
            I => \N__52124\
        );

    \I__12017\ : Span4Mux_h
    port map (
            O => \N__52130\,
            I => \N__52119\
        );

    \I__12016\ : Span4Mux_v
    port map (
            O => \N__52127\,
            I => \N__52119\
        );

    \I__12015\ : LocalMux
    port map (
            O => \N__52124\,
            I => n3109
        );

    \I__12014\ : Odrv4
    port map (
            O => \N__52119\,
            I => n3109
        );

    \I__12013\ : CascadeMux
    port map (
            O => \N__52114\,
            I => \N__52111\
        );

    \I__12012\ : InMux
    port map (
            O => \N__52111\,
            I => \N__52108\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__52108\,
            I => \N__52105\
        );

    \I__12010\ : Span4Mux_v
    port map (
            O => \N__52105\,
            I => \N__52102\
        );

    \I__12009\ : Span4Mux_h
    port map (
            O => \N__52102\,
            I => \N__52099\
        );

    \I__12008\ : Odrv4
    port map (
            O => \N__52099\,
            I => n3176
        );

    \I__12007\ : InMux
    port map (
            O => \N__52096\,
            I => n12516
        );

    \I__12006\ : CascadeMux
    port map (
            O => \N__52093\,
            I => \N__52089\
        );

    \I__12005\ : InMux
    port map (
            O => \N__52092\,
            I => \N__52086\
        );

    \I__12004\ : InMux
    port map (
            O => \N__52089\,
            I => \N__52083\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__52086\,
            I => \N__52078\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__52083\,
            I => \N__52078\
        );

    \I__12001\ : Span4Mux_h
    port map (
            O => \N__52078\,
            I => \N__52074\
        );

    \I__12000\ : InMux
    port map (
            O => \N__52077\,
            I => \N__52071\
        );

    \I__11999\ : Span4Mux_h
    port map (
            O => \N__52074\,
            I => \N__52068\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__52071\,
            I => n3108
        );

    \I__11997\ : Odrv4
    port map (
            O => \N__52068\,
            I => n3108
        );

    \I__11996\ : InMux
    port map (
            O => \N__52063\,
            I => \N__52060\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__52060\,
            I => \N__52057\
        );

    \I__11994\ : Span4Mux_h
    port map (
            O => \N__52057\,
            I => \N__52054\
        );

    \I__11993\ : Span4Mux_h
    port map (
            O => \N__52054\,
            I => \N__52051\
        );

    \I__11992\ : Odrv4
    port map (
            O => \N__52051\,
            I => n3175
        );

    \I__11991\ : InMux
    port map (
            O => \N__52048\,
            I => n12517
        );

    \I__11990\ : InMux
    port map (
            O => \N__52045\,
            I => \N__52042\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__52042\,
            I => \N__52037\
        );

    \I__11988\ : InMux
    port map (
            O => \N__52041\,
            I => \N__52032\
        );

    \I__11987\ : InMux
    port map (
            O => \N__52040\,
            I => \N__52032\
        );

    \I__11986\ : Span4Mux_v
    port map (
            O => \N__52037\,
            I => \N__52029\
        );

    \I__11985\ : LocalMux
    port map (
            O => \N__52032\,
            I => \N__52026\
        );

    \I__11984\ : Span4Mux_h
    port map (
            O => \N__52029\,
            I => \N__52023\
        );

    \I__11983\ : Span4Mux_v
    port map (
            O => \N__52026\,
            I => \N__52020\
        );

    \I__11982\ : Odrv4
    port map (
            O => \N__52023\,
            I => n3107
        );

    \I__11981\ : Odrv4
    port map (
            O => \N__52020\,
            I => n3107
        );

    \I__11980\ : InMux
    port map (
            O => \N__52015\,
            I => \N__52012\
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__52012\,
            I => \N__52009\
        );

    \I__11978\ : Span12Mux_h
    port map (
            O => \N__52009\,
            I => \N__52006\
        );

    \I__11977\ : Odrv12
    port map (
            O => \N__52006\,
            I => n3174
        );

    \I__11976\ : InMux
    port map (
            O => \N__52003\,
            I => n12518
        );

    \I__11975\ : InMux
    port map (
            O => \N__52000\,
            I => \N__51997\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__51997\,
            I => \N__51993\
        );

    \I__11973\ : InMux
    port map (
            O => \N__51996\,
            I => \N__51989\
        );

    \I__11972\ : Span4Mux_h
    port map (
            O => \N__51993\,
            I => \N__51986\
        );

    \I__11971\ : InMux
    port map (
            O => \N__51992\,
            I => \N__51983\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__51989\,
            I => \N__51980\
        );

    \I__11969\ : Span4Mux_h
    port map (
            O => \N__51986\,
            I => \N__51975\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__51983\,
            I => \N__51975\
        );

    \I__11967\ : Odrv4
    port map (
            O => \N__51980\,
            I => n3106
        );

    \I__11966\ : Odrv4
    port map (
            O => \N__51975\,
            I => n3106
        );

    \I__11965\ : InMux
    port map (
            O => \N__51970\,
            I => \N__51967\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__51967\,
            I => \N__51964\
        );

    \I__11963\ : Span4Mux_h
    port map (
            O => \N__51964\,
            I => \N__51961\
        );

    \I__11962\ : Span4Mux_h
    port map (
            O => \N__51961\,
            I => \N__51958\
        );

    \I__11961\ : Odrv4
    port map (
            O => \N__51958\,
            I => n3173
        );

    \I__11960\ : InMux
    port map (
            O => \N__51955\,
            I => n12519
        );

    \I__11959\ : InMux
    port map (
            O => \N__51952\,
            I => \N__51948\
        );

    \I__11958\ : InMux
    port map (
            O => \N__51951\,
            I => \N__51945\
        );

    \I__11957\ : LocalMux
    port map (
            O => \N__51948\,
            I => \N__51942\
        );

    \I__11956\ : LocalMux
    port map (
            O => \N__51945\,
            I => n15158
        );

    \I__11955\ : Odrv12
    port map (
            O => \N__51942\,
            I => n15158
        );

    \I__11954\ : CascadeMux
    port map (
            O => \N__51937\,
            I => \N__51934\
        );

    \I__11953\ : InMux
    port map (
            O => \N__51934\,
            I => \N__51931\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__51931\,
            I => \N__51927\
        );

    \I__11951\ : InMux
    port map (
            O => \N__51930\,
            I => \N__51924\
        );

    \I__11950\ : Span4Mux_v
    port map (
            O => \N__51927\,
            I => \N__51921\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__51924\,
            I => \N__51918\
        );

    \I__11948\ : Odrv4
    port map (
            O => \N__51921\,
            I => n3105
        );

    \I__11947\ : Odrv12
    port map (
            O => \N__51918\,
            I => n3105
        );

    \I__11946\ : InMux
    port map (
            O => \N__51913\,
            I => n12520
        );

    \I__11945\ : CascadeMux
    port map (
            O => \N__51910\,
            I => \N__51906\
        );

    \I__11944\ : InMux
    port map (
            O => \N__51909\,
            I => \N__51903\
        );

    \I__11943\ : InMux
    port map (
            O => \N__51906\,
            I => \N__51900\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__51903\,
            I => \N__51897\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__51900\,
            I => \N__51894\
        );

    \I__11940\ : Span4Mux_h
    port map (
            O => \N__51897\,
            I => \N__51891\
        );

    \I__11939\ : Span4Mux_v
    port map (
            O => \N__51894\,
            I => \N__51888\
        );

    \I__11938\ : Span4Mux_h
    port map (
            O => \N__51891\,
            I => \N__51885\
        );

    \I__11937\ : Odrv4
    port map (
            O => \N__51888\,
            I => n3204
        );

    \I__11936\ : Odrv4
    port map (
            O => \N__51885\,
            I => n3204
        );

    \I__11935\ : InMux
    port map (
            O => \N__51880\,
            I => \N__51876\
        );

    \I__11934\ : InMux
    port map (
            O => \N__51879\,
            I => \N__51872\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__51876\,
            I => \N__51869\
        );

    \I__11932\ : InMux
    port map (
            O => \N__51875\,
            I => \N__51866\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__51872\,
            I => encoder0_position_target_0
        );

    \I__11930\ : Odrv4
    port map (
            O => \N__51869\,
            I => encoder0_position_target_0
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__51866\,
            I => encoder0_position_target_0
        );

    \I__11928\ : InMux
    port map (
            O => \N__51859\,
            I => \bfn_16_26_0_\
        );

    \I__11927\ : InMux
    port map (
            O => \N__51856\,
            I => \N__51853\
        );

    \I__11926\ : LocalMux
    port map (
            O => \N__51853\,
            I => \N__51849\
        );

    \I__11925\ : InMux
    port map (
            O => \N__51852\,
            I => \N__51846\
        );

    \I__11924\ : Span4Mux_h
    port map (
            O => \N__51849\,
            I => \N__51843\
        );

    \I__11923\ : LocalMux
    port map (
            O => \N__51846\,
            I => \N__51839\
        );

    \I__11922\ : Span4Mux_h
    port map (
            O => \N__51843\,
            I => \N__51836\
        );

    \I__11921\ : InMux
    port map (
            O => \N__51842\,
            I => \N__51833\
        );

    \I__11920\ : Odrv4
    port map (
            O => \N__51839\,
            I => n3118
        );

    \I__11919\ : Odrv4
    port map (
            O => \N__51836\,
            I => n3118
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__51833\,
            I => n3118
        );

    \I__11917\ : CascadeMux
    port map (
            O => \N__51826\,
            I => \N__51823\
        );

    \I__11916\ : InMux
    port map (
            O => \N__51823\,
            I => \N__51820\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__51820\,
            I => \N__51817\
        );

    \I__11914\ : Span4Mux_v
    port map (
            O => \N__51817\,
            I => \N__51814\
        );

    \I__11913\ : Span4Mux_h
    port map (
            O => \N__51814\,
            I => \N__51811\
        );

    \I__11912\ : Odrv4
    port map (
            O => \N__51811\,
            I => n3185
        );

    \I__11911\ : InMux
    port map (
            O => \N__51808\,
            I => \bfn_16_24_0_\
        );

    \I__11910\ : CascadeMux
    port map (
            O => \N__51805\,
            I => \N__51801\
        );

    \I__11909\ : InMux
    port map (
            O => \N__51804\,
            I => \N__51798\
        );

    \I__11908\ : InMux
    port map (
            O => \N__51801\,
            I => \N__51795\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__51798\,
            I => \N__51792\
        );

    \I__11906\ : LocalMux
    port map (
            O => \N__51795\,
            I => \N__51789\
        );

    \I__11905\ : Span4Mux_v
    port map (
            O => \N__51792\,
            I => \N__51786\
        );

    \I__11904\ : Span4Mux_v
    port map (
            O => \N__51789\,
            I => \N__51783\
        );

    \I__11903\ : Span4Mux_h
    port map (
            O => \N__51786\,
            I => \N__51780\
        );

    \I__11902\ : Odrv4
    port map (
            O => \N__51783\,
            I => n3117
        );

    \I__11901\ : Odrv4
    port map (
            O => \N__51780\,
            I => n3117
        );

    \I__11900\ : InMux
    port map (
            O => \N__51775\,
            I => \N__51772\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__51772\,
            I => \N__51769\
        );

    \I__11898\ : Span4Mux_v
    port map (
            O => \N__51769\,
            I => \N__51766\
        );

    \I__11897\ : Span4Mux_h
    port map (
            O => \N__51766\,
            I => \N__51763\
        );

    \I__11896\ : Odrv4
    port map (
            O => \N__51763\,
            I => n3184
        );

    \I__11895\ : InMux
    port map (
            O => \N__51760\,
            I => n12508
        );

    \I__11894\ : InMux
    port map (
            O => \N__51757\,
            I => \N__51754\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__51754\,
            I => \N__51751\
        );

    \I__11892\ : Span4Mux_h
    port map (
            O => \N__51751\,
            I => \N__51746\
        );

    \I__11891\ : InMux
    port map (
            O => \N__51750\,
            I => \N__51743\
        );

    \I__11890\ : InMux
    port map (
            O => \N__51749\,
            I => \N__51740\
        );

    \I__11889\ : Span4Mux_v
    port map (
            O => \N__51746\,
            I => \N__51735\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__51743\,
            I => \N__51735\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__51740\,
            I => n3116
        );

    \I__11886\ : Odrv4
    port map (
            O => \N__51735\,
            I => n3116
        );

    \I__11885\ : InMux
    port map (
            O => \N__51730\,
            I => \N__51727\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__51727\,
            I => \N__51724\
        );

    \I__11883\ : Span4Mux_h
    port map (
            O => \N__51724\,
            I => \N__51721\
        );

    \I__11882\ : Odrv4
    port map (
            O => \N__51721\,
            I => n3183
        );

    \I__11881\ : InMux
    port map (
            O => \N__51718\,
            I => n12509
        );

    \I__11880\ : CascadeMux
    port map (
            O => \N__51715\,
            I => \N__51712\
        );

    \I__11879\ : InMux
    port map (
            O => \N__51712\,
            I => \N__51708\
        );

    \I__11878\ : InMux
    port map (
            O => \N__51711\,
            I => \N__51705\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__51708\,
            I => \N__51702\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__51705\,
            I => \N__51699\
        );

    \I__11875\ : Span4Mux_v
    port map (
            O => \N__51702\,
            I => \N__51696\
        );

    \I__11874\ : Span4Mux_v
    port map (
            O => \N__51699\,
            I => \N__51693\
        );

    \I__11873\ : Span4Mux_v
    port map (
            O => \N__51696\,
            I => \N__51688\
        );

    \I__11872\ : Span4Mux_h
    port map (
            O => \N__51693\,
            I => \N__51688\
        );

    \I__11871\ : Odrv4
    port map (
            O => \N__51688\,
            I => n3115
        );

    \I__11870\ : InMux
    port map (
            O => \N__51685\,
            I => \N__51682\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__51682\,
            I => \N__51679\
        );

    \I__11868\ : Span4Mux_v
    port map (
            O => \N__51679\,
            I => \N__51676\
        );

    \I__11867\ : Odrv4
    port map (
            O => \N__51676\,
            I => n3182
        );

    \I__11866\ : InMux
    port map (
            O => \N__51673\,
            I => n12510
        );

    \I__11865\ : InMux
    port map (
            O => \N__51670\,
            I => \N__51667\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__51667\,
            I => \N__51664\
        );

    \I__11863\ : Span4Mux_h
    port map (
            O => \N__51664\,
            I => \N__51660\
        );

    \I__11862\ : InMux
    port map (
            O => \N__51663\,
            I => \N__51657\
        );

    \I__11861\ : Span4Mux_v
    port map (
            O => \N__51660\,
            I => \N__51654\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__51657\,
            I => n3114
        );

    \I__11859\ : Odrv4
    port map (
            O => \N__51654\,
            I => n3114
        );

    \I__11858\ : InMux
    port map (
            O => \N__51649\,
            I => \N__51646\
        );

    \I__11857\ : LocalMux
    port map (
            O => \N__51646\,
            I => n3181
        );

    \I__11856\ : InMux
    port map (
            O => \N__51643\,
            I => n12511
        );

    \I__11855\ : InMux
    port map (
            O => \N__51640\,
            I => \N__51636\
        );

    \I__11854\ : InMux
    port map (
            O => \N__51639\,
            I => \N__51633\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__51636\,
            I => \N__51629\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__51633\,
            I => \N__51626\
        );

    \I__11851\ : InMux
    port map (
            O => \N__51632\,
            I => \N__51623\
        );

    \I__11850\ : Span4Mux_v
    port map (
            O => \N__51629\,
            I => \N__51618\
        );

    \I__11849\ : Span4Mux_h
    port map (
            O => \N__51626\,
            I => \N__51618\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__51623\,
            I => n3113
        );

    \I__11847\ : Odrv4
    port map (
            O => \N__51618\,
            I => n3113
        );

    \I__11846\ : CascadeMux
    port map (
            O => \N__51613\,
            I => \N__51610\
        );

    \I__11845\ : InMux
    port map (
            O => \N__51610\,
            I => \N__51607\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__51607\,
            I => \N__51604\
        );

    \I__11843\ : Span4Mux_h
    port map (
            O => \N__51604\,
            I => \N__51601\
        );

    \I__11842\ : Span4Mux_h
    port map (
            O => \N__51601\,
            I => \N__51598\
        );

    \I__11841\ : Odrv4
    port map (
            O => \N__51598\,
            I => n3180
        );

    \I__11840\ : InMux
    port map (
            O => \N__51595\,
            I => n12512
        );

    \I__11839\ : InMux
    port map (
            O => \N__51592\,
            I => \N__51589\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__51589\,
            I => \N__51585\
        );

    \I__11837\ : InMux
    port map (
            O => \N__51588\,
            I => \N__51582\
        );

    \I__11836\ : Span4Mux_h
    port map (
            O => \N__51585\,
            I => \N__51579\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__51582\,
            I => \N__51576\
        );

    \I__11834\ : Odrv4
    port map (
            O => \N__51579\,
            I => n3112
        );

    \I__11833\ : Odrv4
    port map (
            O => \N__51576\,
            I => n3112
        );

    \I__11832\ : InMux
    port map (
            O => \N__51571\,
            I => \N__51568\
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__51568\,
            I => \N__51565\
        );

    \I__11830\ : Span4Mux_h
    port map (
            O => \N__51565\,
            I => \N__51562\
        );

    \I__11829\ : Odrv4
    port map (
            O => \N__51562\,
            I => n3179
        );

    \I__11828\ : InMux
    port map (
            O => \N__51559\,
            I => n12513
        );

    \I__11827\ : InMux
    port map (
            O => \N__51556\,
            I => \N__51552\
        );

    \I__11826\ : CascadeMux
    port map (
            O => \N__51555\,
            I => \N__51549\
        );

    \I__11825\ : LocalMux
    port map (
            O => \N__51552\,
            I => \N__51545\
        );

    \I__11824\ : InMux
    port map (
            O => \N__51549\,
            I => \N__51542\
        );

    \I__11823\ : InMux
    port map (
            O => \N__51548\,
            I => \N__51539\
        );

    \I__11822\ : Span4Mux_h
    port map (
            O => \N__51545\,
            I => \N__51536\
        );

    \I__11821\ : LocalMux
    port map (
            O => \N__51542\,
            I => \N__51533\
        );

    \I__11820\ : LocalMux
    port map (
            O => \N__51539\,
            I => \N__51530\
        );

    \I__11819\ : Span4Mux_v
    port map (
            O => \N__51536\,
            I => \N__51523\
        );

    \I__11818\ : Span4Mux_v
    port map (
            O => \N__51533\,
            I => \N__51523\
        );

    \I__11817\ : Span4Mux_h
    port map (
            O => \N__51530\,
            I => \N__51523\
        );

    \I__11816\ : Odrv4
    port map (
            O => \N__51523\,
            I => n3126
        );

    \I__11815\ : CascadeMux
    port map (
            O => \N__51520\,
            I => \N__51517\
        );

    \I__11814\ : InMux
    port map (
            O => \N__51517\,
            I => \N__51514\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__51514\,
            I => \N__51511\
        );

    \I__11812\ : Span4Mux_h
    port map (
            O => \N__51511\,
            I => \N__51508\
        );

    \I__11811\ : Span4Mux_h
    port map (
            O => \N__51508\,
            I => \N__51505\
        );

    \I__11810\ : Odrv4
    port map (
            O => \N__51505\,
            I => n3193
        );

    \I__11809\ : InMux
    port map (
            O => \N__51502\,
            I => \bfn_16_23_0_\
        );

    \I__11808\ : InMux
    port map (
            O => \N__51499\,
            I => \N__51494\
        );

    \I__11807\ : InMux
    port map (
            O => \N__51498\,
            I => \N__51491\
        );

    \I__11806\ : InMux
    port map (
            O => \N__51497\,
            I => \N__51488\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__51494\,
            I => \N__51485\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__51491\,
            I => \N__51482\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__51488\,
            I => \N__51479\
        );

    \I__11802\ : Span4Mux_h
    port map (
            O => \N__51485\,
            I => \N__51476\
        );

    \I__11801\ : Span4Mux_h
    port map (
            O => \N__51482\,
            I => \N__51473\
        );

    \I__11800\ : Odrv4
    port map (
            O => \N__51479\,
            I => n3125
        );

    \I__11799\ : Odrv4
    port map (
            O => \N__51476\,
            I => n3125
        );

    \I__11798\ : Odrv4
    port map (
            O => \N__51473\,
            I => n3125
        );

    \I__11797\ : CascadeMux
    port map (
            O => \N__51466\,
            I => \N__51463\
        );

    \I__11796\ : InMux
    port map (
            O => \N__51463\,
            I => \N__51460\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__51460\,
            I => \N__51457\
        );

    \I__11794\ : Span4Mux_v
    port map (
            O => \N__51457\,
            I => \N__51454\
        );

    \I__11793\ : Odrv4
    port map (
            O => \N__51454\,
            I => n3192
        );

    \I__11792\ : InMux
    port map (
            O => \N__51451\,
            I => n12500
        );

    \I__11791\ : InMux
    port map (
            O => \N__51448\,
            I => \N__51445\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__51445\,
            I => \N__51441\
        );

    \I__11789\ : InMux
    port map (
            O => \N__51444\,
            I => \N__51438\
        );

    \I__11788\ : Span4Mux_v
    port map (
            O => \N__51441\,
            I => \N__51435\
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__51438\,
            I => \N__51431\
        );

    \I__11786\ : Span4Mux_h
    port map (
            O => \N__51435\,
            I => \N__51428\
        );

    \I__11785\ : InMux
    port map (
            O => \N__51434\,
            I => \N__51425\
        );

    \I__11784\ : Odrv4
    port map (
            O => \N__51431\,
            I => n3124
        );

    \I__11783\ : Odrv4
    port map (
            O => \N__51428\,
            I => n3124
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__51425\,
            I => n3124
        );

    \I__11781\ : InMux
    port map (
            O => \N__51418\,
            I => \N__51415\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__51415\,
            I => \N__51412\
        );

    \I__11779\ : Odrv12
    port map (
            O => \N__51412\,
            I => n3191
        );

    \I__11778\ : InMux
    port map (
            O => \N__51409\,
            I => n12501
        );

    \I__11777\ : CascadeMux
    port map (
            O => \N__51406\,
            I => \N__51402\
        );

    \I__11776\ : InMux
    port map (
            O => \N__51405\,
            I => \N__51399\
        );

    \I__11775\ : InMux
    port map (
            O => \N__51402\,
            I => \N__51396\
        );

    \I__11774\ : LocalMux
    port map (
            O => \N__51399\,
            I => \N__51392\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__51396\,
            I => \N__51389\
        );

    \I__11772\ : InMux
    port map (
            O => \N__51395\,
            I => \N__51386\
        );

    \I__11771\ : Span4Mux_v
    port map (
            O => \N__51392\,
            I => \N__51383\
        );

    \I__11770\ : Span4Mux_h
    port map (
            O => \N__51389\,
            I => \N__51380\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__51386\,
            I => \N__51377\
        );

    \I__11768\ : Span4Mux_h
    port map (
            O => \N__51383\,
            I => \N__51372\
        );

    \I__11767\ : Span4Mux_v
    port map (
            O => \N__51380\,
            I => \N__51372\
        );

    \I__11766\ : Odrv4
    port map (
            O => \N__51377\,
            I => n3123
        );

    \I__11765\ : Odrv4
    port map (
            O => \N__51372\,
            I => n3123
        );

    \I__11764\ : CascadeMux
    port map (
            O => \N__51367\,
            I => \N__51364\
        );

    \I__11763\ : InMux
    port map (
            O => \N__51364\,
            I => \N__51361\
        );

    \I__11762\ : LocalMux
    port map (
            O => \N__51361\,
            I => \N__51358\
        );

    \I__11761\ : Span4Mux_v
    port map (
            O => \N__51358\,
            I => \N__51355\
        );

    \I__11760\ : Odrv4
    port map (
            O => \N__51355\,
            I => n3190
        );

    \I__11759\ : InMux
    port map (
            O => \N__51352\,
            I => n12502
        );

    \I__11758\ : InMux
    port map (
            O => \N__51349\,
            I => \N__51345\
        );

    \I__11757\ : CascadeMux
    port map (
            O => \N__51348\,
            I => \N__51342\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__51345\,
            I => \N__51339\
        );

    \I__11755\ : InMux
    port map (
            O => \N__51342\,
            I => \N__51336\
        );

    \I__11754\ : Span4Mux_h
    port map (
            O => \N__51339\,
            I => \N__51333\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__51336\,
            I => \N__51330\
        );

    \I__11752\ : Odrv4
    port map (
            O => \N__51333\,
            I => n3122
        );

    \I__11751\ : Odrv12
    port map (
            O => \N__51330\,
            I => n3122
        );

    \I__11750\ : InMux
    port map (
            O => \N__51325\,
            I => \N__51322\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__51322\,
            I => \N__51319\
        );

    \I__11748\ : Span4Mux_v
    port map (
            O => \N__51319\,
            I => \N__51316\
        );

    \I__11747\ : Odrv4
    port map (
            O => \N__51316\,
            I => n3189
        );

    \I__11746\ : InMux
    port map (
            O => \N__51313\,
            I => n12503
        );

    \I__11745\ : InMux
    port map (
            O => \N__51310\,
            I => \N__51306\
        );

    \I__11744\ : InMux
    port map (
            O => \N__51309\,
            I => \N__51303\
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__51306\,
            I => \N__51300\
        );

    \I__11742\ : LocalMux
    port map (
            O => \N__51303\,
            I => \N__51297\
        );

    \I__11741\ : Span4Mux_h
    port map (
            O => \N__51300\,
            I => \N__51294\
        );

    \I__11740\ : Odrv12
    port map (
            O => \N__51297\,
            I => n3121
        );

    \I__11739\ : Odrv4
    port map (
            O => \N__51294\,
            I => n3121
        );

    \I__11738\ : InMux
    port map (
            O => \N__51289\,
            I => \N__51286\
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__51286\,
            I => \N__51283\
        );

    \I__11736\ : Span4Mux_h
    port map (
            O => \N__51283\,
            I => \N__51280\
        );

    \I__11735\ : Odrv4
    port map (
            O => \N__51280\,
            I => n3188
        );

    \I__11734\ : InMux
    port map (
            O => \N__51277\,
            I => n12504
        );

    \I__11733\ : InMux
    port map (
            O => \N__51274\,
            I => \N__51269\
        );

    \I__11732\ : InMux
    port map (
            O => \N__51273\,
            I => \N__51266\
        );

    \I__11731\ : InMux
    port map (
            O => \N__51272\,
            I => \N__51263\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__51269\,
            I => \N__51260\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__51266\,
            I => \N__51257\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__51263\,
            I => \N__51254\
        );

    \I__11727\ : Span4Mux_h
    port map (
            O => \N__51260\,
            I => \N__51251\
        );

    \I__11726\ : Span4Mux_h
    port map (
            O => \N__51257\,
            I => \N__51248\
        );

    \I__11725\ : Odrv4
    port map (
            O => \N__51254\,
            I => n3120
        );

    \I__11724\ : Odrv4
    port map (
            O => \N__51251\,
            I => n3120
        );

    \I__11723\ : Odrv4
    port map (
            O => \N__51248\,
            I => n3120
        );

    \I__11722\ : CascadeMux
    port map (
            O => \N__51241\,
            I => \N__51238\
        );

    \I__11721\ : InMux
    port map (
            O => \N__51238\,
            I => \N__51235\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__51235\,
            I => \N__51232\
        );

    \I__11719\ : Span4Mux_h
    port map (
            O => \N__51232\,
            I => \N__51229\
        );

    \I__11718\ : Odrv4
    port map (
            O => \N__51229\,
            I => n3187
        );

    \I__11717\ : InMux
    port map (
            O => \N__51226\,
            I => n12505
        );

    \I__11716\ : InMux
    port map (
            O => \N__51223\,
            I => \N__51219\
        );

    \I__11715\ : InMux
    port map (
            O => \N__51222\,
            I => \N__51216\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__51219\,
            I => \N__51213\
        );

    \I__11713\ : LocalMux
    port map (
            O => \N__51216\,
            I => \N__51207\
        );

    \I__11712\ : Span12Mux_v
    port map (
            O => \N__51213\,
            I => \N__51207\
        );

    \I__11711\ : InMux
    port map (
            O => \N__51212\,
            I => \N__51204\
        );

    \I__11710\ : Odrv12
    port map (
            O => \N__51207\,
            I => n3119
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__51204\,
            I => n3119
        );

    \I__11708\ : CascadeMux
    port map (
            O => \N__51199\,
            I => \N__51196\
        );

    \I__11707\ : InMux
    port map (
            O => \N__51196\,
            I => \N__51193\
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__51193\,
            I => \N__51190\
        );

    \I__11705\ : Span4Mux_h
    port map (
            O => \N__51190\,
            I => \N__51187\
        );

    \I__11704\ : Odrv4
    port map (
            O => \N__51187\,
            I => n3186
        );

    \I__11703\ : InMux
    port map (
            O => \N__51184\,
            I => n12506
        );

    \I__11702\ : InMux
    port map (
            O => \N__51181\,
            I => \N__51177\
        );

    \I__11701\ : InMux
    port map (
            O => \N__51180\,
            I => \N__51173\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__51177\,
            I => \N__51170\
        );

    \I__11699\ : InMux
    port map (
            O => \N__51176\,
            I => \N__51167\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__51173\,
            I => \N__51164\
        );

    \I__11697\ : Span4Mux_v
    port map (
            O => \N__51170\,
            I => \N__51159\
        );

    \I__11696\ : LocalMux
    port map (
            O => \N__51167\,
            I => \N__51159\
        );

    \I__11695\ : Sp12to4
    port map (
            O => \N__51164\,
            I => \N__51156\
        );

    \I__11694\ : Span4Mux_h
    port map (
            O => \N__51159\,
            I => \N__51153\
        );

    \I__11693\ : Span12Mux_v
    port map (
            O => \N__51156\,
            I => \N__51150\
        );

    \I__11692\ : Span4Mux_v
    port map (
            O => \N__51153\,
            I => \N__51147\
        );

    \I__11691\ : Span12Mux_h
    port map (
            O => \N__51150\,
            I => \N__51144\
        );

    \I__11690\ : Odrv4
    port map (
            O => \N__51147\,
            I => n317
        );

    \I__11689\ : Odrv12
    port map (
            O => \N__51144\,
            I => n317
        );

    \I__11688\ : InMux
    port map (
            O => \N__51139\,
            I => \N__51136\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__51136\,
            I => \N__51133\
        );

    \I__11686\ : Span4Mux_h
    port map (
            O => \N__51133\,
            I => \N__51130\
        );

    \I__11685\ : Span4Mux_h
    port map (
            O => \N__51130\,
            I => \N__51127\
        );

    \I__11684\ : Span4Mux_h
    port map (
            O => \N__51127\,
            I => \N__51124\
        );

    \I__11683\ : Odrv4
    port map (
            O => \N__51124\,
            I => n3201
        );

    \I__11682\ : InMux
    port map (
            O => \N__51121\,
            I => \bfn_16_22_0_\
        );

    \I__11681\ : CascadeMux
    port map (
            O => \N__51118\,
            I => \N__51114\
        );

    \I__11680\ : CascadeMux
    port map (
            O => \N__51117\,
            I => \N__51111\
        );

    \I__11679\ : InMux
    port map (
            O => \N__51114\,
            I => \N__51107\
        );

    \I__11678\ : InMux
    port map (
            O => \N__51111\,
            I => \N__51102\
        );

    \I__11677\ : InMux
    port map (
            O => \N__51110\,
            I => \N__51102\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__51107\,
            I => \N__51099\
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__51102\,
            I => n3133
        );

    \I__11674\ : Odrv12
    port map (
            O => \N__51099\,
            I => n3133
        );

    \I__11673\ : InMux
    port map (
            O => \N__51094\,
            I => \N__51091\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__51091\,
            I => \N__51088\
        );

    \I__11671\ : Span4Mux_h
    port map (
            O => \N__51088\,
            I => \N__51085\
        );

    \I__11670\ : Span4Mux_h
    port map (
            O => \N__51085\,
            I => \N__51082\
        );

    \I__11669\ : Odrv4
    port map (
            O => \N__51082\,
            I => n3200
        );

    \I__11668\ : InMux
    port map (
            O => \N__51079\,
            I => n12492
        );

    \I__11667\ : CascadeMux
    port map (
            O => \N__51076\,
            I => \N__51073\
        );

    \I__11666\ : InMux
    port map (
            O => \N__51073\,
            I => \N__51070\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__51070\,
            I => \N__51065\
        );

    \I__11664\ : InMux
    port map (
            O => \N__51069\,
            I => \N__51062\
        );

    \I__11663\ : CascadeMux
    port map (
            O => \N__51068\,
            I => \N__51059\
        );

    \I__11662\ : Span4Mux_h
    port map (
            O => \N__51065\,
            I => \N__51056\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__51062\,
            I => \N__51053\
        );

    \I__11660\ : InMux
    port map (
            O => \N__51059\,
            I => \N__51050\
        );

    \I__11659\ : Span4Mux_h
    port map (
            O => \N__51056\,
            I => \N__51047\
        );

    \I__11658\ : Odrv4
    port map (
            O => \N__51053\,
            I => n3132
        );

    \I__11657\ : LocalMux
    port map (
            O => \N__51050\,
            I => n3132
        );

    \I__11656\ : Odrv4
    port map (
            O => \N__51047\,
            I => n3132
        );

    \I__11655\ : CascadeMux
    port map (
            O => \N__51040\,
            I => \N__51037\
        );

    \I__11654\ : InMux
    port map (
            O => \N__51037\,
            I => \N__51034\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__51034\,
            I => \N__51031\
        );

    \I__11652\ : Span4Mux_v
    port map (
            O => \N__51031\,
            I => \N__51028\
        );

    \I__11651\ : Span4Mux_h
    port map (
            O => \N__51028\,
            I => \N__51025\
        );

    \I__11650\ : Odrv4
    port map (
            O => \N__51025\,
            I => n3199
        );

    \I__11649\ : InMux
    port map (
            O => \N__51022\,
            I => n12493
        );

    \I__11648\ : CascadeMux
    port map (
            O => \N__51019\,
            I => \N__51016\
        );

    \I__11647\ : InMux
    port map (
            O => \N__51016\,
            I => \N__51013\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__51013\,
            I => \N__51008\
        );

    \I__11645\ : InMux
    port map (
            O => \N__51012\,
            I => \N__51003\
        );

    \I__11644\ : InMux
    port map (
            O => \N__51011\,
            I => \N__51003\
        );

    \I__11643\ : Odrv12
    port map (
            O => \N__51008\,
            I => n3131
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__51003\,
            I => n3131
        );

    \I__11641\ : InMux
    port map (
            O => \N__50998\,
            I => \N__50995\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__50995\,
            I => \N__50992\
        );

    \I__11639\ : Span12Mux_s10_v
    port map (
            O => \N__50992\,
            I => \N__50989\
        );

    \I__11638\ : Odrv12
    port map (
            O => \N__50989\,
            I => n3198
        );

    \I__11637\ : InMux
    port map (
            O => \N__50986\,
            I => n12494
        );

    \I__11636\ : CascadeMux
    port map (
            O => \N__50983\,
            I => \N__50979\
        );

    \I__11635\ : InMux
    port map (
            O => \N__50982\,
            I => \N__50975\
        );

    \I__11634\ : InMux
    port map (
            O => \N__50979\,
            I => \N__50972\
        );

    \I__11633\ : InMux
    port map (
            O => \N__50978\,
            I => \N__50969\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__50975\,
            I => \N__50966\
        );

    \I__11631\ : LocalMux
    port map (
            O => \N__50972\,
            I => \N__50963\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__50969\,
            I => \N__50960\
        );

    \I__11629\ : Span4Mux_v
    port map (
            O => \N__50966\,
            I => \N__50953\
        );

    \I__11628\ : Span4Mux_h
    port map (
            O => \N__50963\,
            I => \N__50953\
        );

    \I__11627\ : Span4Mux_v
    port map (
            O => \N__50960\,
            I => \N__50953\
        );

    \I__11626\ : Odrv4
    port map (
            O => \N__50953\,
            I => n3130
        );

    \I__11625\ : CascadeMux
    port map (
            O => \N__50950\,
            I => \N__50947\
        );

    \I__11624\ : InMux
    port map (
            O => \N__50947\,
            I => \N__50944\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__50944\,
            I => \N__50941\
        );

    \I__11622\ : Span4Mux_h
    port map (
            O => \N__50941\,
            I => \N__50938\
        );

    \I__11621\ : Span4Mux_h
    port map (
            O => \N__50938\,
            I => \N__50935\
        );

    \I__11620\ : Odrv4
    port map (
            O => \N__50935\,
            I => n3197
        );

    \I__11619\ : InMux
    port map (
            O => \N__50932\,
            I => n12495
        );

    \I__11618\ : InMux
    port map (
            O => \N__50929\,
            I => \N__50925\
        );

    \I__11617\ : InMux
    port map (
            O => \N__50928\,
            I => \N__50921\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__50925\,
            I => \N__50918\
        );

    \I__11615\ : InMux
    port map (
            O => \N__50924\,
            I => \N__50915\
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__50921\,
            I => \N__50912\
        );

    \I__11613\ : Span4Mux_h
    port map (
            O => \N__50918\,
            I => \N__50909\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__50915\,
            I => \N__50906\
        );

    \I__11611\ : Span4Mux_h
    port map (
            O => \N__50912\,
            I => \N__50903\
        );

    \I__11610\ : Odrv4
    port map (
            O => \N__50909\,
            I => n3129
        );

    \I__11609\ : Odrv12
    port map (
            O => \N__50906\,
            I => n3129
        );

    \I__11608\ : Odrv4
    port map (
            O => \N__50903\,
            I => n3129
        );

    \I__11607\ : CascadeMux
    port map (
            O => \N__50896\,
            I => \N__50893\
        );

    \I__11606\ : InMux
    port map (
            O => \N__50893\,
            I => \N__50890\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__50890\,
            I => \N__50887\
        );

    \I__11604\ : Span4Mux_h
    port map (
            O => \N__50887\,
            I => \N__50884\
        );

    \I__11603\ : Odrv4
    port map (
            O => \N__50884\,
            I => n3196
        );

    \I__11602\ : InMux
    port map (
            O => \N__50881\,
            I => n12496
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__50878\,
            I => \N__50874\
        );

    \I__11600\ : InMux
    port map (
            O => \N__50877\,
            I => \N__50871\
        );

    \I__11599\ : InMux
    port map (
            O => \N__50874\,
            I => \N__50868\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__50871\,
            I => \N__50865\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__50868\,
            I => \N__50862\
        );

    \I__11596\ : Span4Mux_v
    port map (
            O => \N__50865\,
            I => \N__50859\
        );

    \I__11595\ : Span4Mux_h
    port map (
            O => \N__50862\,
            I => \N__50856\
        );

    \I__11594\ : Span4Mux_v
    port map (
            O => \N__50859\,
            I => \N__50852\
        );

    \I__11593\ : Span4Mux_h
    port map (
            O => \N__50856\,
            I => \N__50849\
        );

    \I__11592\ : InMux
    port map (
            O => \N__50855\,
            I => \N__50846\
        );

    \I__11591\ : Odrv4
    port map (
            O => \N__50852\,
            I => n3128
        );

    \I__11590\ : Odrv4
    port map (
            O => \N__50849\,
            I => n3128
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__50846\,
            I => n3128
        );

    \I__11588\ : InMux
    port map (
            O => \N__50839\,
            I => \N__50836\
        );

    \I__11587\ : LocalMux
    port map (
            O => \N__50836\,
            I => \N__50833\
        );

    \I__11586\ : Span4Mux_v
    port map (
            O => \N__50833\,
            I => \N__50830\
        );

    \I__11585\ : Odrv4
    port map (
            O => \N__50830\,
            I => n3195
        );

    \I__11584\ : InMux
    port map (
            O => \N__50827\,
            I => n12497
        );

    \I__11583\ : CascadeMux
    port map (
            O => \N__50824\,
            I => \N__50821\
        );

    \I__11582\ : InMux
    port map (
            O => \N__50821\,
            I => \N__50817\
        );

    \I__11581\ : CascadeMux
    port map (
            O => \N__50820\,
            I => \N__50814\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__50817\,
            I => \N__50811\
        );

    \I__11579\ : InMux
    port map (
            O => \N__50814\,
            I => \N__50808\
        );

    \I__11578\ : Span4Mux_v
    port map (
            O => \N__50811\,
            I => \N__50803\
        );

    \I__11577\ : LocalMux
    port map (
            O => \N__50808\,
            I => \N__50803\
        );

    \I__11576\ : Span4Mux_v
    port map (
            O => \N__50803\,
            I => \N__50800\
        );

    \I__11575\ : Span4Mux_h
    port map (
            O => \N__50800\,
            I => \N__50796\
        );

    \I__11574\ : InMux
    port map (
            O => \N__50799\,
            I => \N__50793\
        );

    \I__11573\ : Odrv4
    port map (
            O => \N__50796\,
            I => n3127
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__50793\,
            I => n3127
        );

    \I__11571\ : InMux
    port map (
            O => \N__50788\,
            I => \N__50785\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__50785\,
            I => \N__50782\
        );

    \I__11569\ : Odrv4
    port map (
            O => \N__50782\,
            I => n3194
        );

    \I__11568\ : InMux
    port map (
            O => \N__50779\,
            I => n12498
        );

    \I__11567\ : InMux
    port map (
            O => \N__50776\,
            I => \N__50772\
        );

    \I__11566\ : InMux
    port map (
            O => \N__50775\,
            I => \N__50769\
        );

    \I__11565\ : LocalMux
    port map (
            O => \N__50772\,
            I => sweep_counter_10
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__50769\,
            I => sweep_counter_10
        );

    \I__11563\ : InMux
    port map (
            O => \N__50764\,
            I => n12615
        );

    \I__11562\ : InMux
    port map (
            O => \N__50761\,
            I => \N__50757\
        );

    \I__11561\ : InMux
    port map (
            O => \N__50760\,
            I => \N__50754\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__50757\,
            I => sweep_counter_11
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__50754\,
            I => sweep_counter_11
        );

    \I__11558\ : InMux
    port map (
            O => \N__50749\,
            I => n12616
        );

    \I__11557\ : InMux
    port map (
            O => \N__50746\,
            I => \N__50742\
        );

    \I__11556\ : InMux
    port map (
            O => \N__50745\,
            I => \N__50739\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__50742\,
            I => sweep_counter_12
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__50739\,
            I => sweep_counter_12
        );

    \I__11553\ : InMux
    port map (
            O => \N__50734\,
            I => n12617
        );

    \I__11552\ : InMux
    port map (
            O => \N__50731\,
            I => \N__50727\
        );

    \I__11551\ : InMux
    port map (
            O => \N__50730\,
            I => \N__50724\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__50727\,
            I => sweep_counter_13
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__50724\,
            I => sweep_counter_13
        );

    \I__11548\ : InMux
    port map (
            O => \N__50719\,
            I => n12618
        );

    \I__11547\ : CascadeMux
    port map (
            O => \N__50716\,
            I => \N__50712\
        );

    \I__11546\ : InMux
    port map (
            O => \N__50715\,
            I => \N__50709\
        );

    \I__11545\ : InMux
    port map (
            O => \N__50712\,
            I => \N__50706\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__50709\,
            I => sweep_counter_14
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__50706\,
            I => sweep_counter_14
        );

    \I__11542\ : InMux
    port map (
            O => \N__50701\,
            I => n12619
        );

    \I__11541\ : CascadeMux
    port map (
            O => \N__50698\,
            I => \N__50694\
        );

    \I__11540\ : InMux
    port map (
            O => \N__50697\,
            I => \N__50691\
        );

    \I__11539\ : InMux
    port map (
            O => \N__50694\,
            I => \N__50688\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__50691\,
            I => sweep_counter_15
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__50688\,
            I => sweep_counter_15
        );

    \I__11536\ : InMux
    port map (
            O => \N__50683\,
            I => n12620
        );

    \I__11535\ : InMux
    port map (
            O => \N__50680\,
            I => \N__50676\
        );

    \I__11534\ : InMux
    port map (
            O => \N__50679\,
            I => \N__50673\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__50676\,
            I => sweep_counter_16
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__50673\,
            I => sweep_counter_16
        );

    \I__11531\ : InMux
    port map (
            O => \N__50668\,
            I => \bfn_16_19_0_\
        );

    \I__11530\ : InMux
    port map (
            O => \N__50665\,
            I => n12622
        );

    \I__11529\ : InMux
    port map (
            O => \N__50662\,
            I => \N__50658\
        );

    \I__11528\ : InMux
    port map (
            O => \N__50661\,
            I => \N__50655\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__50658\,
            I => sweep_counter_17
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__50655\,
            I => sweep_counter_17
        );

    \I__11525\ : InMux
    port map (
            O => \N__50650\,
            I => \N__50646\
        );

    \I__11524\ : InMux
    port map (
            O => \N__50649\,
            I => \N__50643\
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__50646\,
            I => sweep_counter_1
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__50643\,
            I => sweep_counter_1
        );

    \I__11521\ : InMux
    port map (
            O => \N__50638\,
            I => n12606
        );

    \I__11520\ : CascadeMux
    port map (
            O => \N__50635\,
            I => \N__50631\
        );

    \I__11519\ : InMux
    port map (
            O => \N__50634\,
            I => \N__50628\
        );

    \I__11518\ : InMux
    port map (
            O => \N__50631\,
            I => \N__50625\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__50628\,
            I => sweep_counter_2
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__50625\,
            I => sweep_counter_2
        );

    \I__11515\ : InMux
    port map (
            O => \N__50620\,
            I => n12607
        );

    \I__11514\ : InMux
    port map (
            O => \N__50617\,
            I => \N__50613\
        );

    \I__11513\ : InMux
    port map (
            O => \N__50616\,
            I => \N__50610\
        );

    \I__11512\ : LocalMux
    port map (
            O => \N__50613\,
            I => sweep_counter_3
        );

    \I__11511\ : LocalMux
    port map (
            O => \N__50610\,
            I => sweep_counter_3
        );

    \I__11510\ : InMux
    port map (
            O => \N__50605\,
            I => n12608
        );

    \I__11509\ : InMux
    port map (
            O => \N__50602\,
            I => \N__50598\
        );

    \I__11508\ : InMux
    port map (
            O => \N__50601\,
            I => \N__50595\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__50598\,
            I => sweep_counter_4
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__50595\,
            I => sweep_counter_4
        );

    \I__11505\ : InMux
    port map (
            O => \N__50590\,
            I => n12609
        );

    \I__11504\ : InMux
    port map (
            O => \N__50587\,
            I => \N__50583\
        );

    \I__11503\ : InMux
    port map (
            O => \N__50586\,
            I => \N__50580\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__50583\,
            I => sweep_counter_5
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__50580\,
            I => sweep_counter_5
        );

    \I__11500\ : InMux
    port map (
            O => \N__50575\,
            I => n12610
        );

    \I__11499\ : CascadeMux
    port map (
            O => \N__50572\,
            I => \N__50568\
        );

    \I__11498\ : InMux
    port map (
            O => \N__50571\,
            I => \N__50565\
        );

    \I__11497\ : InMux
    port map (
            O => \N__50568\,
            I => \N__50562\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__50565\,
            I => \N__50557\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__50562\,
            I => \N__50557\
        );

    \I__11494\ : Odrv4
    port map (
            O => \N__50557\,
            I => sweep_counter_6
        );

    \I__11493\ : InMux
    port map (
            O => \N__50554\,
            I => n12611
        );

    \I__11492\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50547\
        );

    \I__11491\ : InMux
    port map (
            O => \N__50550\,
            I => \N__50544\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__50547\,
            I => sweep_counter_7
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__50544\,
            I => sweep_counter_7
        );

    \I__11488\ : InMux
    port map (
            O => \N__50539\,
            I => n12612
        );

    \I__11487\ : InMux
    port map (
            O => \N__50536\,
            I => \N__50532\
        );

    \I__11486\ : InMux
    port map (
            O => \N__50535\,
            I => \N__50529\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__50532\,
            I => sweep_counter_8
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__50529\,
            I => sweep_counter_8
        );

    \I__11483\ : InMux
    port map (
            O => \N__50524\,
            I => \bfn_16_18_0_\
        );

    \I__11482\ : InMux
    port map (
            O => \N__50521\,
            I => \N__50517\
        );

    \I__11481\ : InMux
    port map (
            O => \N__50520\,
            I => \N__50514\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__50517\,
            I => sweep_counter_9
        );

    \I__11479\ : LocalMux
    port map (
            O => \N__50514\,
            I => sweep_counter_9
        );

    \I__11478\ : InMux
    port map (
            O => \N__50509\,
            I => n12614
        );

    \I__11477\ : CascadeMux
    port map (
            O => \N__50506\,
            I => \quad_counter0.direction_N_534_cascade_\
        );

    \I__11476\ : InMux
    port map (
            O => \N__50503\,
            I => \N__50500\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__50500\,
            I => \quad_counter0.a_prev_N_537\
        );

    \I__11474\ : CascadeMux
    port map (
            O => \N__50497\,
            I => \N__50494\
        );

    \I__11473\ : InMux
    port map (
            O => \N__50494\,
            I => \N__50488\
        );

    \I__11472\ : InMux
    port map (
            O => \N__50493\,
            I => \N__50488\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__50488\,
            I => \quad_counter0.a_prev\
        );

    \I__11470\ : InMux
    port map (
            O => \N__50485\,
            I => \N__50473\
        );

    \I__11469\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50473\
        );

    \I__11468\ : InMux
    port map (
            O => \N__50483\,
            I => \N__50473\
        );

    \I__11467\ : InMux
    port map (
            O => \N__50482\,
            I => \N__50473\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__50473\,
            I => \quad_counter0.b_new_1\
        );

    \I__11465\ : CascadeMux
    port map (
            O => \N__50470\,
            I => \N__50466\
        );

    \I__11464\ : InMux
    port map (
            O => \N__50469\,
            I => \N__50462\
        );

    \I__11463\ : InMux
    port map (
            O => \N__50466\,
            I => \N__50457\
        );

    \I__11462\ : InMux
    port map (
            O => \N__50465\,
            I => \N__50457\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__50462\,
            I => \N__50452\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__50457\,
            I => \N__50452\
        );

    \I__11459\ : Odrv12
    port map (
            O => \N__50452\,
            I => \quad_counter0.b_new_0\
        );

    \I__11458\ : InMux
    port map (
            O => \N__50449\,
            I => \N__50440\
        );

    \I__11457\ : InMux
    port map (
            O => \N__50448\,
            I => \N__50440\
        );

    \I__11456\ : InMux
    port map (
            O => \N__50447\,
            I => \N__50440\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__50440\,
            I => \quad_counter0.debounce_cnt\
        );

    \I__11454\ : CEMux
    port map (
            O => \N__50437\,
            I => \N__50433\
        );

    \I__11453\ : CEMux
    port map (
            O => \N__50436\,
            I => \N__50428\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__50433\,
            I => \N__50425\
        );

    \I__11451\ : CEMux
    port map (
            O => \N__50432\,
            I => \N__50422\
        );

    \I__11450\ : CEMux
    port map (
            O => \N__50431\,
            I => \N__50419\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__50428\,
            I => \N__50416\
        );

    \I__11448\ : Span4Mux_v
    port map (
            O => \N__50425\,
            I => \N__50411\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__50422\,
            I => \N__50411\
        );

    \I__11446\ : LocalMux
    port map (
            O => \N__50419\,
            I => \N__50408\
        );

    \I__11445\ : Span4Mux_v
    port map (
            O => \N__50416\,
            I => \N__50403\
        );

    \I__11444\ : Span4Mux_h
    port map (
            O => \N__50411\,
            I => \N__50403\
        );

    \I__11443\ : Span4Mux_h
    port map (
            O => \N__50408\,
            I => \N__50400\
        );

    \I__11442\ : Span4Mux_h
    port map (
            O => \N__50403\,
            I => \N__50397\
        );

    \I__11441\ : Span4Mux_h
    port map (
            O => \N__50400\,
            I => \N__50394\
        );

    \I__11440\ : Span4Mux_h
    port map (
            O => \N__50397\,
            I => \N__50390\
        );

    \I__11439\ : Span4Mux_h
    port map (
            O => \N__50394\,
            I => \N__50387\
        );

    \I__11438\ : InMux
    port map (
            O => \N__50393\,
            I => \N__50384\
        );

    \I__11437\ : Odrv4
    port map (
            O => \N__50390\,
            I => \direction_N_531\
        );

    \I__11436\ : Odrv4
    port map (
            O => \N__50387\,
            I => \direction_N_531\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__50384\,
            I => \direction_N_531\
        );

    \I__11434\ : CascadeMux
    port map (
            O => \N__50377\,
            I => \N__50373\
        );

    \I__11433\ : InMux
    port map (
            O => \N__50376\,
            I => \N__50368\
        );

    \I__11432\ : InMux
    port map (
            O => \N__50373\,
            I => \N__50365\
        );

    \I__11431\ : InMux
    port map (
            O => \N__50372\,
            I => \N__50362\
        );

    \I__11430\ : InMux
    port map (
            O => \N__50371\,
            I => \N__50359\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__50368\,
            I => \N__50356\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__50365\,
            I => b_prev
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__50362\,
            I => b_prev
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__50359\,
            I => b_prev
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__50356\,
            I => b_prev
        );

    \I__11424\ : InMux
    port map (
            O => \N__50347\,
            I => \N__50344\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__50344\,
            I => n1185
        );

    \I__11422\ : InMux
    port map (
            O => \N__50341\,
            I => \N__50338\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__50338\,
            I => \N__50335\
        );

    \I__11420\ : Span4Mux_s3_v
    port map (
            O => \N__50335\,
            I => \N__50330\
        );

    \I__11419\ : InMux
    port map (
            O => \N__50334\,
            I => \N__50325\
        );

    \I__11418\ : InMux
    port map (
            O => \N__50333\,
            I => \N__50325\
        );

    \I__11417\ : Sp12to4
    port map (
            O => \N__50330\,
            I => \N__50320\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__50325\,
            I => \N__50320\
        );

    \I__11415\ : Odrv12
    port map (
            O => \N__50320\,
            I => \quad_counter0.a_new_0\
        );

    \I__11414\ : CascadeMux
    port map (
            O => \N__50317\,
            I => \N__50311\
        );

    \I__11413\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50306\
        );

    \I__11412\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50303\
        );

    \I__11411\ : InMux
    port map (
            O => \N__50314\,
            I => \N__50298\
        );

    \I__11410\ : InMux
    port map (
            O => \N__50311\,
            I => \N__50298\
        );

    \I__11409\ : InMux
    port map (
            O => \N__50310\,
            I => \N__50293\
        );

    \I__11408\ : InMux
    port map (
            O => \N__50309\,
            I => \N__50293\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__50306\,
            I => \N__50290\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__50303\,
            I => a_new_1
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__50298\,
            I => a_new_1
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__50293\,
            I => a_new_1
        );

    \I__11403\ : Odrv4
    port map (
            O => \N__50290\,
            I => a_new_1
        );

    \I__11402\ : InMux
    port map (
            O => \N__50281\,
            I => \N__50278\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__50278\,
            I => \N__50274\
        );

    \I__11400\ : InMux
    port map (
            O => \N__50277\,
            I => \N__50271\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__50274\,
            I => \N__50268\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__50271\,
            I => \N__50265\
        );

    \I__11397\ : Odrv4
    port map (
            O => \N__50268\,
            I => duty_19
        );

    \I__11396\ : Odrv4
    port map (
            O => \N__50265\,
            I => duty_19
        );

    \I__11395\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50257\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__50257\,
            I => \N__50254\
        );

    \I__11393\ : Odrv4
    port map (
            O => \N__50254\,
            I => n6_adj_572
        );

    \I__11392\ : InMux
    port map (
            O => \N__50251\,
            I => \N__50247\
        );

    \I__11391\ : InMux
    port map (
            O => \N__50250\,
            I => \N__50244\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__50247\,
            I => \N__50241\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__50244\,
            I => \N__50238\
        );

    \I__11388\ : Odrv4
    port map (
            O => \N__50241\,
            I => duty_18
        );

    \I__11387\ : Odrv4
    port map (
            O => \N__50238\,
            I => duty_18
        );

    \I__11386\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50230\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__50230\,
            I => \N__50227\
        );

    \I__11384\ : Span4Mux_h
    port map (
            O => \N__50227\,
            I => \N__50224\
        );

    \I__11383\ : Odrv4
    port map (
            O => \N__50224\,
            I => n7_adj_573
        );

    \I__11382\ : InMux
    port map (
            O => \N__50221\,
            I => \N__50217\
        );

    \I__11381\ : InMux
    port map (
            O => \N__50220\,
            I => \N__50214\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__50217\,
            I => sweep_counter_0
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__50214\,
            I => sweep_counter_0
        );

    \I__11378\ : InMux
    port map (
            O => \N__50209\,
            I => \bfn_16_17_0_\
        );

    \I__11377\ : InMux
    port map (
            O => \N__50206\,
            I => \N__50203\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__50203\,
            I => \N__50200\
        );

    \I__11375\ : Odrv4
    port map (
            O => \N__50200\,
            I => n24_adj_590
        );

    \I__11374\ : InMux
    port map (
            O => \N__50197\,
            I => \N__50194\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__50194\,
            I => \N__50191\
        );

    \I__11372\ : Span4Mux_v
    port map (
            O => \N__50191\,
            I => \N__50187\
        );

    \I__11371\ : InMux
    port map (
            O => \N__50190\,
            I => \N__50184\
        );

    \I__11370\ : Span4Mux_h
    port map (
            O => \N__50187\,
            I => \N__50181\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__50184\,
            I => \N__50178\
        );

    \I__11368\ : Odrv4
    port map (
            O => \N__50181\,
            I => duty_3
        );

    \I__11367\ : Odrv4
    port map (
            O => \N__50178\,
            I => duty_3
        );

    \I__11366\ : InMux
    port map (
            O => \N__50173\,
            I => \N__50170\
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__50170\,
            I => \N__50167\
        );

    \I__11364\ : Odrv4
    port map (
            O => \N__50167\,
            I => n22_adj_588
        );

    \I__11363\ : CascadeMux
    port map (
            O => \N__50164\,
            I => \n21_adj_700_cascade_\
        );

    \I__11362\ : InMux
    port map (
            O => \N__50161\,
            I => \N__50158\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__50158\,
            I => n22_adj_699
        );

    \I__11360\ : InMux
    port map (
            O => \N__50155\,
            I => \N__50151\
        );

    \I__11359\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50148\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__50151\,
            I => \N__50143\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__50148\,
            I => \N__50143\
        );

    \I__11356\ : Span4Mux_h
    port map (
            O => \N__50143\,
            I => \N__50140\
        );

    \I__11355\ : Odrv4
    port map (
            O => \N__50140\,
            I => duty_1
        );

    \I__11354\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50134\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__50134\,
            I => \N__50131\
        );

    \I__11352\ : Odrv4
    port map (
            O => \N__50131\,
            I => \pwm_setpoint_23_N_171_1\
        );

    \I__11351\ : InMux
    port map (
            O => \N__50128\,
            I => \N__50125\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__50125\,
            I => pwm_setpoint_1
        );

    \I__11349\ : CascadeMux
    port map (
            O => \N__50122\,
            I => \quad_counter0.a_prev_N_537_cascade_\
        );

    \I__11348\ : CascadeMux
    port map (
            O => \N__50119\,
            I => \N__50114\
        );

    \I__11347\ : CascadeMux
    port map (
            O => \N__50118\,
            I => \N__50110\
        );

    \I__11346\ : InMux
    port map (
            O => \N__50117\,
            I => \N__50098\
        );

    \I__11345\ : InMux
    port map (
            O => \N__50114\,
            I => \N__50098\
        );

    \I__11344\ : InMux
    port map (
            O => \N__50113\,
            I => \N__50098\
        );

    \I__11343\ : InMux
    port map (
            O => \N__50110\,
            I => \N__50090\
        );

    \I__11342\ : InMux
    port map (
            O => \N__50109\,
            I => \N__50090\
        );

    \I__11341\ : InMux
    port map (
            O => \N__50108\,
            I => \N__50087\
        );

    \I__11340\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50082\
        );

    \I__11339\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50079\
        );

    \I__11338\ : CascadeMux
    port map (
            O => \N__50105\,
            I => \N__50074\
        );

    \I__11337\ : LocalMux
    port map (
            O => \N__50098\,
            I => \N__50065\
        );

    \I__11336\ : InMux
    port map (
            O => \N__50097\,
            I => \N__50058\
        );

    \I__11335\ : InMux
    port map (
            O => \N__50096\,
            I => \N__50058\
        );

    \I__11334\ : InMux
    port map (
            O => \N__50095\,
            I => \N__50058\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__50090\,
            I => \N__50053\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__50087\,
            I => \N__50053\
        );

    \I__11331\ : InMux
    port map (
            O => \N__50086\,
            I => \N__50048\
        );

    \I__11330\ : InMux
    port map (
            O => \N__50085\,
            I => \N__50048\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__50082\,
            I => \N__50045\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__50079\,
            I => \N__50042\
        );

    \I__11327\ : InMux
    port map (
            O => \N__50078\,
            I => \N__50033\
        );

    \I__11326\ : InMux
    port map (
            O => \N__50077\,
            I => \N__50033\
        );

    \I__11325\ : InMux
    port map (
            O => \N__50074\,
            I => \N__50033\
        );

    \I__11324\ : InMux
    port map (
            O => \N__50073\,
            I => \N__50033\
        );

    \I__11323\ : CascadeMux
    port map (
            O => \N__50072\,
            I => \N__50029\
        );

    \I__11322\ : CascadeMux
    port map (
            O => \N__50071\,
            I => \N__50026\
        );

    \I__11321\ : CascadeMux
    port map (
            O => \N__50070\,
            I => \N__50020\
        );

    \I__11320\ : CascadeMux
    port map (
            O => \N__50069\,
            I => \N__50016\
        );

    \I__11319\ : InMux
    port map (
            O => \N__50068\,
            I => \N__50010\
        );

    \I__11318\ : Sp12to4
    port map (
            O => \N__50065\,
            I => \N__50005\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__50058\,
            I => \N__50005\
        );

    \I__11316\ : Span4Mux_h
    port map (
            O => \N__50053\,
            I => \N__50002\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__50048\,
            I => \N__49999\
        );

    \I__11314\ : Span4Mux_v
    port map (
            O => \N__50045\,
            I => \N__49992\
        );

    \I__11313\ : Span4Mux_v
    port map (
            O => \N__50042\,
            I => \N__49992\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__50033\,
            I => \N__49992\
        );

    \I__11311\ : InMux
    port map (
            O => \N__50032\,
            I => \N__49989\
        );

    \I__11310\ : InMux
    port map (
            O => \N__50029\,
            I => \N__49980\
        );

    \I__11309\ : InMux
    port map (
            O => \N__50026\,
            I => \N__49980\
        );

    \I__11308\ : InMux
    port map (
            O => \N__50025\,
            I => \N__49980\
        );

    \I__11307\ : InMux
    port map (
            O => \N__50024\,
            I => \N__49980\
        );

    \I__11306\ : InMux
    port map (
            O => \N__50023\,
            I => \N__49977\
        );

    \I__11305\ : InMux
    port map (
            O => \N__50020\,
            I => \N__49972\
        );

    \I__11304\ : InMux
    port map (
            O => \N__50019\,
            I => \N__49972\
        );

    \I__11303\ : InMux
    port map (
            O => \N__50016\,
            I => \N__49963\
        );

    \I__11302\ : InMux
    port map (
            O => \N__50015\,
            I => \N__49963\
        );

    \I__11301\ : InMux
    port map (
            O => \N__50014\,
            I => \N__49963\
        );

    \I__11300\ : InMux
    port map (
            O => \N__50013\,
            I => \N__49963\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__50010\,
            I => \N__49958\
        );

    \I__11298\ : Span12Mux_s8_v
    port map (
            O => \N__50005\,
            I => \N__49958\
        );

    \I__11297\ : Span4Mux_h
    port map (
            O => \N__50002\,
            I => \N__49955\
        );

    \I__11296\ : Span4Mux_h
    port map (
            O => \N__49999\,
            I => \N__49950\
        );

    \I__11295\ : Span4Mux_h
    port map (
            O => \N__49992\,
            I => \N__49950\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__49989\,
            I => n3138
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__49980\,
            I => n3138
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__49977\,
            I => n3138
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__49972\,
            I => n3138
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__49963\,
            I => n3138
        );

    \I__11289\ : Odrv12
    port map (
            O => \N__49958\,
            I => n3138
        );

    \I__11288\ : Odrv4
    port map (
            O => \N__49955\,
            I => n3138
        );

    \I__11287\ : Odrv4
    port map (
            O => \N__49950\,
            I => n3138
        );

    \I__11286\ : CascadeMux
    port map (
            O => \N__49933\,
            I => \n3114_cascade_\
        );

    \I__11285\ : InMux
    port map (
            O => \N__49930\,
            I => \N__49925\
        );

    \I__11284\ : InMux
    port map (
            O => \N__49929\,
            I => \N__49922\
        );

    \I__11283\ : InMux
    port map (
            O => \N__49928\,
            I => \N__49919\
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__49925\,
            I => \N__49916\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__49922\,
            I => \N__49913\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__49919\,
            I => \N__49910\
        );

    \I__11279\ : Span4Mux_h
    port map (
            O => \N__49916\,
            I => \N__49907\
        );

    \I__11278\ : Odrv4
    port map (
            O => \N__49913\,
            I => n3213
        );

    \I__11277\ : Odrv4
    port map (
            O => \N__49910\,
            I => n3213
        );

    \I__11276\ : Odrv4
    port map (
            O => \N__49907\,
            I => n3213
        );

    \I__11275\ : CascadeMux
    port map (
            O => \N__49900\,
            I => \n7_adj_712_cascade_\
        );

    \I__11274\ : InMux
    port map (
            O => \N__49897\,
            I => \N__49894\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__49894\,
            I => n8_adj_711
        );

    \I__11272\ : CascadeMux
    port map (
            O => \N__49891\,
            I => \N__49876\
        );

    \I__11271\ : CascadeMux
    port map (
            O => \N__49890\,
            I => \N__49872\
        );

    \I__11270\ : CascadeMux
    port map (
            O => \N__49889\,
            I => \N__49868\
        );

    \I__11269\ : CascadeMux
    port map (
            O => \N__49888\,
            I => \N__49864\
        );

    \I__11268\ : CascadeMux
    port map (
            O => \N__49887\,
            I => \N__49861\
        );

    \I__11267\ : CascadeMux
    port map (
            O => \N__49886\,
            I => \N__49857\
        );

    \I__11266\ : CascadeMux
    port map (
            O => \N__49885\,
            I => \N__49853\
        );

    \I__11265\ : CascadeMux
    port map (
            O => \N__49884\,
            I => \N__49849\
        );

    \I__11264\ : CascadeMux
    port map (
            O => \N__49883\,
            I => \N__49845\
        );

    \I__11263\ : CascadeMux
    port map (
            O => \N__49882\,
            I => \N__49841\
        );

    \I__11262\ : CascadeMux
    port map (
            O => \N__49881\,
            I => \N__49837\
        );

    \I__11261\ : CascadeMux
    port map (
            O => \N__49880\,
            I => \N__49833\
        );

    \I__11260\ : InMux
    port map (
            O => \N__49879\,
            I => \N__49812\
        );

    \I__11259\ : InMux
    port map (
            O => \N__49876\,
            I => \N__49812\
        );

    \I__11258\ : InMux
    port map (
            O => \N__49875\,
            I => \N__49812\
        );

    \I__11257\ : InMux
    port map (
            O => \N__49872\,
            I => \N__49812\
        );

    \I__11256\ : InMux
    port map (
            O => \N__49871\,
            I => \N__49812\
        );

    \I__11255\ : InMux
    port map (
            O => \N__49868\,
            I => \N__49812\
        );

    \I__11254\ : InMux
    port map (
            O => \N__49867\,
            I => \N__49812\
        );

    \I__11253\ : InMux
    port map (
            O => \N__49864\,
            I => \N__49812\
        );

    \I__11252\ : InMux
    port map (
            O => \N__49861\,
            I => \N__49795\
        );

    \I__11251\ : InMux
    port map (
            O => \N__49860\,
            I => \N__49795\
        );

    \I__11250\ : InMux
    port map (
            O => \N__49857\,
            I => \N__49795\
        );

    \I__11249\ : InMux
    port map (
            O => \N__49856\,
            I => \N__49795\
        );

    \I__11248\ : InMux
    port map (
            O => \N__49853\,
            I => \N__49795\
        );

    \I__11247\ : InMux
    port map (
            O => \N__49852\,
            I => \N__49795\
        );

    \I__11246\ : InMux
    port map (
            O => \N__49849\,
            I => \N__49795\
        );

    \I__11245\ : InMux
    port map (
            O => \N__49848\,
            I => \N__49795\
        );

    \I__11244\ : InMux
    port map (
            O => \N__49845\,
            I => \N__49778\
        );

    \I__11243\ : InMux
    port map (
            O => \N__49844\,
            I => \N__49778\
        );

    \I__11242\ : InMux
    port map (
            O => \N__49841\,
            I => \N__49778\
        );

    \I__11241\ : InMux
    port map (
            O => \N__49840\,
            I => \N__49778\
        );

    \I__11240\ : InMux
    port map (
            O => \N__49837\,
            I => \N__49778\
        );

    \I__11239\ : InMux
    port map (
            O => \N__49836\,
            I => \N__49778\
        );

    \I__11238\ : InMux
    port map (
            O => \N__49833\,
            I => \N__49778\
        );

    \I__11237\ : InMux
    port map (
            O => \N__49832\,
            I => \N__49778\
        );

    \I__11236\ : CascadeMux
    port map (
            O => \N__49831\,
            I => \N__49774\
        );

    \I__11235\ : CascadeMux
    port map (
            O => \N__49830\,
            I => \N__49770\
        );

    \I__11234\ : CascadeMux
    port map (
            O => \N__49829\,
            I => \N__49766\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__49812\,
            I => \N__49758\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__49795\,
            I => \N__49758\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__49778\,
            I => \N__49758\
        );

    \I__11230\ : InMux
    port map (
            O => \N__49777\,
            I => \N__49743\
        );

    \I__11229\ : InMux
    port map (
            O => \N__49774\,
            I => \N__49743\
        );

    \I__11228\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49743\
        );

    \I__11227\ : InMux
    port map (
            O => \N__49770\,
            I => \N__49743\
        );

    \I__11226\ : InMux
    port map (
            O => \N__49769\,
            I => \N__49743\
        );

    \I__11225\ : InMux
    port map (
            O => \N__49766\,
            I => \N__49743\
        );

    \I__11224\ : InMux
    port map (
            O => \N__49765\,
            I => \N__49743\
        );

    \I__11223\ : Span4Mux_v
    port map (
            O => \N__49758\,
            I => \N__49740\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__49743\,
            I => \N__49737\
        );

    \I__11221\ : Span4Mux_h
    port map (
            O => \N__49740\,
            I => \N__49732\
        );

    \I__11220\ : Span4Mux_h
    port map (
            O => \N__49737\,
            I => \N__49732\
        );

    \I__11219\ : Span4Mux_v
    port map (
            O => \N__49732\,
            I => \N__49729\
        );

    \I__11218\ : Span4Mux_h
    port map (
            O => \N__49729\,
            I => \N__49726\
        );

    \I__11217\ : Odrv4
    port map (
            O => \N__49726\,
            I => \quad_counter0.direction_N_530\
        );

    \I__11216\ : InMux
    port map (
            O => \N__49723\,
            I => \N__49720\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__49720\,
            I => n13676
        );

    \I__11214\ : CascadeMux
    port map (
            O => \N__49717\,
            I => \n10_adj_714_cascade_\
        );

    \I__11213\ : CascadeMux
    port map (
            O => \N__49714\,
            I => \n16_adj_702_cascade_\
        );

    \I__11212\ : InMux
    port map (
            O => \N__49711\,
            I => \N__49708\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__49708\,
            I => n19_adj_701
        );

    \I__11210\ : InMux
    port map (
            O => \N__49705\,
            I => \N__49702\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__49702\,
            I => \N__49699\
        );

    \I__11208\ : Span4Mux_v
    port map (
            O => \N__49699\,
            I => \N__49696\
        );

    \I__11207\ : Odrv4
    port map (
            O => \N__49696\,
            I => n3286
        );

    \I__11206\ : CascadeMux
    port map (
            O => \N__49693\,
            I => \n27_adj_709_cascade_\
        );

    \I__11205\ : InMux
    port map (
            O => \N__49690\,
            I => \N__49685\
        );

    \I__11204\ : InMux
    port map (
            O => \N__49689\,
            I => \N__49682\
        );

    \I__11203\ : InMux
    port map (
            O => \N__49688\,
            I => \N__49679\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__49685\,
            I => n3219
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__49682\,
            I => n3219
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__49679\,
            I => n3219
        );

    \I__11199\ : InMux
    port map (
            O => \N__49672\,
            I => \N__49669\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__49669\,
            I => n13830
        );

    \I__11197\ : InMux
    port map (
            O => \N__49666\,
            I => \N__49663\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__49663\,
            I => \N__49660\
        );

    \I__11195\ : Odrv4
    port map (
            O => \N__49660\,
            I => n3292
        );

    \I__11194\ : CascadeMux
    port map (
            O => \N__49657\,
            I => \N__49652\
        );

    \I__11193\ : InMux
    port map (
            O => \N__49656\,
            I => \N__49649\
        );

    \I__11192\ : InMux
    port map (
            O => \N__49655\,
            I => \N__49646\
        );

    \I__11191\ : InMux
    port map (
            O => \N__49652\,
            I => \N__49643\
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__49649\,
            I => \N__49640\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__49646\,
            I => \N__49637\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__49643\,
            I => \N__49634\
        );

    \I__11187\ : Span4Mux_v
    port map (
            O => \N__49640\,
            I => \N__49629\
        );

    \I__11186\ : Span4Mux_h
    port map (
            O => \N__49637\,
            I => \N__49629\
        );

    \I__11185\ : Span4Mux_h
    port map (
            O => \N__49634\,
            I => \N__49626\
        );

    \I__11184\ : Span4Mux_h
    port map (
            O => \N__49629\,
            I => \N__49623\
        );

    \I__11183\ : Odrv4
    port map (
            O => \N__49626\,
            I => n3225
        );

    \I__11182\ : Odrv4
    port map (
            O => \N__49623\,
            I => n3225
        );

    \I__11181\ : InMux
    port map (
            O => \N__49618\,
            I => \N__49609\
        );

    \I__11180\ : InMux
    port map (
            O => \N__49617\,
            I => \N__49593\
        );

    \I__11179\ : InMux
    port map (
            O => \N__49616\,
            I => \N__49593\
        );

    \I__11178\ : InMux
    port map (
            O => \N__49615\,
            I => \N__49593\
        );

    \I__11177\ : InMux
    port map (
            O => \N__49614\,
            I => \N__49593\
        );

    \I__11176\ : InMux
    port map (
            O => \N__49613\,
            I => \N__49593\
        );

    \I__11175\ : CascadeMux
    port map (
            O => \N__49612\,
            I => \N__49590\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__49609\,
            I => \N__49586\
        );

    \I__11173\ : CascadeMux
    port map (
            O => \N__49608\,
            I => \N__49578\
        );

    \I__11172\ : CascadeMux
    port map (
            O => \N__49607\,
            I => \N__49574\
        );

    \I__11171\ : CascadeMux
    port map (
            O => \N__49606\,
            I => \N__49570\
        );

    \I__11170\ : CascadeMux
    port map (
            O => \N__49605\,
            I => \N__49558\
        );

    \I__11169\ : CascadeMux
    port map (
            O => \N__49604\,
            I => \N__49555\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__49593\,
            I => \N__49551\
        );

    \I__11167\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49546\
        );

    \I__11166\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49546\
        );

    \I__11165\ : Span4Mux_v
    port map (
            O => \N__49586\,
            I => \N__49543\
        );

    \I__11164\ : InMux
    port map (
            O => \N__49585\,
            I => \N__49530\
        );

    \I__11163\ : InMux
    port map (
            O => \N__49584\,
            I => \N__49530\
        );

    \I__11162\ : InMux
    port map (
            O => \N__49583\,
            I => \N__49530\
        );

    \I__11161\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49530\
        );

    \I__11160\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49530\
        );

    \I__11159\ : InMux
    port map (
            O => \N__49578\,
            I => \N__49530\
        );

    \I__11158\ : InMux
    port map (
            O => \N__49577\,
            I => \N__49519\
        );

    \I__11157\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49519\
        );

    \I__11156\ : InMux
    port map (
            O => \N__49573\,
            I => \N__49519\
        );

    \I__11155\ : InMux
    port map (
            O => \N__49570\,
            I => \N__49519\
        );

    \I__11154\ : InMux
    port map (
            O => \N__49569\,
            I => \N__49519\
        );

    \I__11153\ : InMux
    port map (
            O => \N__49568\,
            I => \N__49506\
        );

    \I__11152\ : InMux
    port map (
            O => \N__49567\,
            I => \N__49506\
        );

    \I__11151\ : InMux
    port map (
            O => \N__49566\,
            I => \N__49506\
        );

    \I__11150\ : InMux
    port map (
            O => \N__49565\,
            I => \N__49506\
        );

    \I__11149\ : InMux
    port map (
            O => \N__49564\,
            I => \N__49506\
        );

    \I__11148\ : InMux
    port map (
            O => \N__49563\,
            I => \N__49506\
        );

    \I__11147\ : InMux
    port map (
            O => \N__49562\,
            I => \N__49495\
        );

    \I__11146\ : InMux
    port map (
            O => \N__49561\,
            I => \N__49495\
        );

    \I__11145\ : InMux
    port map (
            O => \N__49558\,
            I => \N__49495\
        );

    \I__11144\ : InMux
    port map (
            O => \N__49555\,
            I => \N__49495\
        );

    \I__11143\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49495\
        );

    \I__11142\ : Span4Mux_h
    port map (
            O => \N__49551\,
            I => \N__49490\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__49546\,
            I => \N__49490\
        );

    \I__11140\ : Odrv4
    port map (
            O => \N__49543\,
            I => n3237
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__49530\,
            I => n3237
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__49519\,
            I => n3237
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__49506\,
            I => n3237
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__49495\,
            I => n3237
        );

    \I__11135\ : Odrv4
    port map (
            O => \N__49490\,
            I => n3237
        );

    \I__11134\ : InMux
    port map (
            O => \N__49477\,
            I => \N__49474\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__49474\,
            I => n21_adj_706
        );

    \I__11132\ : InMux
    port map (
            O => \N__49471\,
            I => \N__49467\
        );

    \I__11131\ : InMux
    port map (
            O => \N__49470\,
            I => \N__49464\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__49467\,
            I => \N__49458\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__49464\,
            I => \N__49458\
        );

    \I__11128\ : InMux
    port map (
            O => \N__49463\,
            I => \N__49455\
        );

    \I__11127\ : Span4Mux_v
    port map (
            O => \N__49458\,
            I => \N__49450\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__49455\,
            I => \N__49450\
        );

    \I__11125\ : Odrv4
    port map (
            O => \N__49450\,
            I => n3011
        );

    \I__11124\ : CascadeMux
    port map (
            O => \N__49447\,
            I => \N__49444\
        );

    \I__11123\ : InMux
    port map (
            O => \N__49444\,
            I => \N__49441\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__49441\,
            I => \N__49438\
        );

    \I__11121\ : Span4Mux_h
    port map (
            O => \N__49438\,
            I => \N__49435\
        );

    \I__11120\ : Odrv4
    port map (
            O => \N__49435\,
            I => n3078
        );

    \I__11119\ : CascadeMux
    port map (
            O => \N__49432\,
            I => \n3110_cascade_\
        );

    \I__11118\ : InMux
    port map (
            O => \N__49429\,
            I => \N__49424\
        );

    \I__11117\ : InMux
    port map (
            O => \N__49428\,
            I => \N__49421\
        );

    \I__11116\ : InMux
    port map (
            O => \N__49427\,
            I => \N__49418\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__49424\,
            I => \N__49413\
        );

    \I__11114\ : LocalMux
    port map (
            O => \N__49421\,
            I => \N__49413\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__49418\,
            I => \N__49408\
        );

    \I__11112\ : Span4Mux_v
    port map (
            O => \N__49413\,
            I => \N__49408\
        );

    \I__11111\ : Span4Mux_h
    port map (
            O => \N__49408\,
            I => \N__49405\
        );

    \I__11110\ : Odrv4
    port map (
            O => \N__49405\,
            I => n3209
        );

    \I__11109\ : CascadeMux
    port map (
            O => \N__49402\,
            I => \N__49399\
        );

    \I__11108\ : InMux
    port map (
            O => \N__49399\,
            I => \N__49395\
        );

    \I__11107\ : InMux
    port map (
            O => \N__49398\,
            I => \N__49392\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__49395\,
            I => \N__49387\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__49392\,
            I => \N__49387\
        );

    \I__11104\ : Span4Mux_h
    port map (
            O => \N__49387\,
            I => \N__49383\
        );

    \I__11103\ : InMux
    port map (
            O => \N__49386\,
            I => \N__49380\
        );

    \I__11102\ : Odrv4
    port map (
            O => \N__49383\,
            I => n3226
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__49380\,
            I => n3226
        );

    \I__11100\ : CascadeMux
    port map (
            O => \N__49375\,
            I => \N__49368\
        );

    \I__11099\ : InMux
    port map (
            O => \N__49374\,
            I => \N__49363\
        );

    \I__11098\ : InMux
    port map (
            O => \N__49373\,
            I => \N__49360\
        );

    \I__11097\ : InMux
    port map (
            O => \N__49372\,
            I => \N__49355\
        );

    \I__11096\ : InMux
    port map (
            O => \N__49371\,
            I => \N__49350\
        );

    \I__11095\ : InMux
    port map (
            O => \N__49368\,
            I => \N__49347\
        );

    \I__11094\ : InMux
    port map (
            O => \N__49367\,
            I => \N__49344\
        );

    \I__11093\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49341\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__49363\,
            I => \N__49337\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__49360\,
            I => \N__49333\
        );

    \I__11090\ : InMux
    port map (
            O => \N__49359\,
            I => \N__49330\
        );

    \I__11089\ : CascadeMux
    port map (
            O => \N__49358\,
            I => \N__49327\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__49355\,
            I => \N__49321\
        );

    \I__11087\ : CascadeMux
    port map (
            O => \N__49354\,
            I => \N__49317\
        );

    \I__11086\ : CascadeMux
    port map (
            O => \N__49353\,
            I => \N__49313\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__49350\,
            I => \N__49303\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__49347\,
            I => \N__49303\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__49344\,
            I => \N__49303\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__49341\,
            I => \N__49303\
        );

    \I__11081\ : CascadeMux
    port map (
            O => \N__49340\,
            I => \N__49299\
        );

    \I__11080\ : Span4Mux_v
    port map (
            O => \N__49337\,
            I => \N__49289\
        );

    \I__11079\ : InMux
    port map (
            O => \N__49336\,
            I => \N__49286\
        );

    \I__11078\ : Span4Mux_h
    port map (
            O => \N__49333\,
            I => \N__49281\
        );

    \I__11077\ : LocalMux
    port map (
            O => \N__49330\,
            I => \N__49281\
        );

    \I__11076\ : InMux
    port map (
            O => \N__49327\,
            I => \N__49274\
        );

    \I__11075\ : InMux
    port map (
            O => \N__49326\,
            I => \N__49274\
        );

    \I__11074\ : InMux
    port map (
            O => \N__49325\,
            I => \N__49274\
        );

    \I__11073\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49270\
        );

    \I__11072\ : Span4Mux_v
    port map (
            O => \N__49321\,
            I => \N__49267\
        );

    \I__11071\ : InMux
    port map (
            O => \N__49320\,
            I => \N__49264\
        );

    \I__11070\ : InMux
    port map (
            O => \N__49317\,
            I => \N__49255\
        );

    \I__11069\ : InMux
    port map (
            O => \N__49316\,
            I => \N__49255\
        );

    \I__11068\ : InMux
    port map (
            O => \N__49313\,
            I => \N__49255\
        );

    \I__11067\ : InMux
    port map (
            O => \N__49312\,
            I => \N__49255\
        );

    \I__11066\ : Span4Mux_v
    port map (
            O => \N__49303\,
            I => \N__49252\
        );

    \I__11065\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49245\
        );

    \I__11064\ : InMux
    port map (
            O => \N__49299\,
            I => \N__49245\
        );

    \I__11063\ : InMux
    port map (
            O => \N__49298\,
            I => \N__49245\
        );

    \I__11062\ : InMux
    port map (
            O => \N__49297\,
            I => \N__49232\
        );

    \I__11061\ : InMux
    port map (
            O => \N__49296\,
            I => \N__49232\
        );

    \I__11060\ : InMux
    port map (
            O => \N__49295\,
            I => \N__49232\
        );

    \I__11059\ : InMux
    port map (
            O => \N__49294\,
            I => \N__49232\
        );

    \I__11058\ : InMux
    port map (
            O => \N__49293\,
            I => \N__49232\
        );

    \I__11057\ : InMux
    port map (
            O => \N__49292\,
            I => \N__49232\
        );

    \I__11056\ : Span4Mux_h
    port map (
            O => \N__49289\,
            I => \N__49223\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__49286\,
            I => \N__49223\
        );

    \I__11054\ : Span4Mux_v
    port map (
            O => \N__49281\,
            I => \N__49223\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__49274\,
            I => \N__49223\
        );

    \I__11052\ : InMux
    port map (
            O => \N__49273\,
            I => \N__49220\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__49270\,
            I => n2841
        );

    \I__11050\ : Odrv4
    port map (
            O => \N__49267\,
            I => n2841
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__49264\,
            I => n2841
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__49255\,
            I => n2841
        );

    \I__11047\ : Odrv4
    port map (
            O => \N__49252\,
            I => n2841
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__49245\,
            I => n2841
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__49232\,
            I => n2841
        );

    \I__11044\ : Odrv4
    port map (
            O => \N__49223\,
            I => n2841
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__49220\,
            I => n2841
        );

    \I__11042\ : InMux
    port map (
            O => \N__49201\,
            I => \N__49198\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__49198\,
            I => \N__49195\
        );

    \I__11040\ : Span4Mux_h
    port map (
            O => \N__49195\,
            I => \N__49192\
        );

    \I__11039\ : Odrv4
    port map (
            O => \N__49192\,
            I => n14921
        );

    \I__11038\ : InMux
    port map (
            O => \N__49189\,
            I => \N__49186\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__49186\,
            I => \N__49182\
        );

    \I__11036\ : InMux
    port map (
            O => \N__49185\,
            I => \N__49179\
        );

    \I__11035\ : Span4Mux_h
    port map (
            O => \N__49182\,
            I => \N__49174\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__49179\,
            I => \N__49174\
        );

    \I__11033\ : Span4Mux_v
    port map (
            O => \N__49174\,
            I => \N__49170\
        );

    \I__11032\ : InMux
    port map (
            O => \N__49173\,
            I => \N__49167\
        );

    \I__11031\ : Odrv4
    port map (
            O => \N__49170\,
            I => n3009
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__49167\,
            I => n3009
        );

    \I__11029\ : CascadeMux
    port map (
            O => \N__49162\,
            I => \N__49159\
        );

    \I__11028\ : InMux
    port map (
            O => \N__49159\,
            I => \N__49156\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__49156\,
            I => n3076
        );

    \I__11026\ : InMux
    port map (
            O => \N__49153\,
            I => \N__49150\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__49150\,
            I => \N__49147\
        );

    \I__11024\ : Span4Mux_v
    port map (
            O => \N__49147\,
            I => \N__49144\
        );

    \I__11023\ : Span4Mux_h
    port map (
            O => \N__49144\,
            I => \N__49141\
        );

    \I__11022\ : Span4Mux_h
    port map (
            O => \N__49141\,
            I => \N__49138\
        );

    \I__11021\ : Span4Mux_v
    port map (
            O => \N__49138\,
            I => \N__49135\
        );

    \I__11020\ : Sp12to4
    port map (
            O => \N__49135\,
            I => \N__49132\
        );

    \I__11019\ : Odrv12
    port map (
            O => \N__49132\,
            I => \ENCODER0_B_N\
        );

    \I__11018\ : InMux
    port map (
            O => \N__49129\,
            I => \N__49126\
        );

    \I__11017\ : LocalMux
    port map (
            O => \N__49126\,
            I => \N__49122\
        );

    \I__11016\ : InMux
    port map (
            O => \N__49125\,
            I => \N__49119\
        );

    \I__11015\ : Span4Mux_v
    port map (
            O => \N__49122\,
            I => \N__49115\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__49119\,
            I => \N__49112\
        );

    \I__11013\ : InMux
    port map (
            O => \N__49118\,
            I => \N__49109\
        );

    \I__11012\ : Span4Mux_h
    port map (
            O => \N__49115\,
            I => \N__49106\
        );

    \I__11011\ : Span4Mux_v
    port map (
            O => \N__49112\,
            I => \N__49101\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__49109\,
            I => \N__49101\
        );

    \I__11009\ : Odrv4
    port map (
            O => \N__49106\,
            I => n3015
        );

    \I__11008\ : Odrv4
    port map (
            O => \N__49101\,
            I => n3015
        );

    \I__11007\ : CascadeMux
    port map (
            O => \N__49096\,
            I => \N__49093\
        );

    \I__11006\ : InMux
    port map (
            O => \N__49093\,
            I => \N__49090\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__49090\,
            I => \N__49087\
        );

    \I__11004\ : Odrv4
    port map (
            O => \N__49087\,
            I => n3082
        );

    \I__11003\ : CascadeMux
    port map (
            O => \N__49084\,
            I => \N__49070\
        );

    \I__11002\ : CascadeMux
    port map (
            O => \N__49083\,
            I => \N__49066\
        );

    \I__11001\ : CascadeMux
    port map (
            O => \N__49082\,
            I => \N__49060\
        );

    \I__11000\ : CascadeMux
    port map (
            O => \N__49081\,
            I => \N__49057\
        );

    \I__10999\ : InMux
    port map (
            O => \N__49080\,
            I => \N__49054\
        );

    \I__10998\ : CascadeMux
    port map (
            O => \N__49079\,
            I => \N__49051\
        );

    \I__10997\ : InMux
    port map (
            O => \N__49078\,
            I => \N__49044\
        );

    \I__10996\ : InMux
    port map (
            O => \N__49077\,
            I => \N__49044\
        );

    \I__10995\ : InMux
    port map (
            O => \N__49076\,
            I => \N__49044\
        );

    \I__10994\ : InMux
    port map (
            O => \N__49075\,
            I => \N__49036\
        );

    \I__10993\ : InMux
    port map (
            O => \N__49074\,
            I => \N__49031\
        );

    \I__10992\ : InMux
    port map (
            O => \N__49073\,
            I => \N__49031\
        );

    \I__10991\ : InMux
    port map (
            O => \N__49070\,
            I => \N__49026\
        );

    \I__10990\ : InMux
    port map (
            O => \N__49069\,
            I => \N__49026\
        );

    \I__10989\ : InMux
    port map (
            O => \N__49066\,
            I => \N__49021\
        );

    \I__10988\ : InMux
    port map (
            O => \N__49065\,
            I => \N__49021\
        );

    \I__10987\ : InMux
    port map (
            O => \N__49064\,
            I => \N__49010\
        );

    \I__10986\ : InMux
    port map (
            O => \N__49063\,
            I => \N__49010\
        );

    \I__10985\ : InMux
    port map (
            O => \N__49060\,
            I => \N__49010\
        );

    \I__10984\ : InMux
    port map (
            O => \N__49057\,
            I => \N__49010\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__49054\,
            I => \N__49007\
        );

    \I__10982\ : InMux
    port map (
            O => \N__49051\,
            I => \N__49004\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__49044\,
            I => \N__49001\
        );

    \I__10980\ : CascadeMux
    port map (
            O => \N__49043\,
            I => \N__48996\
        );

    \I__10979\ : CascadeMux
    port map (
            O => \N__49042\,
            I => \N__48992\
        );

    \I__10978\ : CascadeMux
    port map (
            O => \N__49041\,
            I => \N__48989\
        );

    \I__10977\ : CascadeMux
    port map (
            O => \N__49040\,
            I => \N__48985\
        );

    \I__10976\ : CascadeMux
    port map (
            O => \N__49039\,
            I => \N__48982\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__49036\,
            I => \N__48973\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__49031\,
            I => \N__48973\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__49026\,
            I => \N__48973\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__49021\,
            I => \N__48970\
        );

    \I__10971\ : InMux
    port map (
            O => \N__49020\,
            I => \N__48967\
        );

    \I__10970\ : InMux
    port map (
            O => \N__49019\,
            I => \N__48964\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__49010\,
            I => \N__48961\
        );

    \I__10968\ : Span4Mux_h
    port map (
            O => \N__49007\,
            I => \N__48954\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__49004\,
            I => \N__48954\
        );

    \I__10966\ : Span4Mux_h
    port map (
            O => \N__49001\,
            I => \N__48954\
        );

    \I__10965\ : InMux
    port map (
            O => \N__49000\,
            I => \N__48945\
        );

    \I__10964\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48945\
        );

    \I__10963\ : InMux
    port map (
            O => \N__48996\,
            I => \N__48945\
        );

    \I__10962\ : InMux
    port map (
            O => \N__48995\,
            I => \N__48945\
        );

    \I__10961\ : InMux
    port map (
            O => \N__48992\,
            I => \N__48938\
        );

    \I__10960\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48938\
        );

    \I__10959\ : InMux
    port map (
            O => \N__48988\,
            I => \N__48938\
        );

    \I__10958\ : InMux
    port map (
            O => \N__48985\,
            I => \N__48929\
        );

    \I__10957\ : InMux
    port map (
            O => \N__48982\,
            I => \N__48929\
        );

    \I__10956\ : InMux
    port map (
            O => \N__48981\,
            I => \N__48929\
        );

    \I__10955\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48929\
        );

    \I__10954\ : Span4Mux_h
    port map (
            O => \N__48973\,
            I => \N__48924\
        );

    \I__10953\ : Span4Mux_h
    port map (
            O => \N__48970\,
            I => \N__48924\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__48967\,
            I => n3039
        );

    \I__10951\ : LocalMux
    port map (
            O => \N__48964\,
            I => n3039
        );

    \I__10950\ : Odrv4
    port map (
            O => \N__48961\,
            I => n3039
        );

    \I__10949\ : Odrv4
    port map (
            O => \N__48954\,
            I => n3039
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__48945\,
            I => n3039
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__48938\,
            I => n3039
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__48929\,
            I => n3039
        );

    \I__10945\ : Odrv4
    port map (
            O => \N__48924\,
            I => n3039
        );

    \I__10944\ : InMux
    port map (
            O => \N__48907\,
            I => \N__48903\
        );

    \I__10943\ : CascadeMux
    port map (
            O => \N__48906\,
            I => \N__48900\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__48903\,
            I => \N__48897\
        );

    \I__10941\ : InMux
    port map (
            O => \N__48900\,
            I => \N__48893\
        );

    \I__10940\ : Span4Mux_v
    port map (
            O => \N__48897\,
            I => \N__48890\
        );

    \I__10939\ : InMux
    port map (
            O => \N__48896\,
            I => \N__48887\
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__48893\,
            I => n2810
        );

    \I__10937\ : Odrv4
    port map (
            O => \N__48890\,
            I => n2810
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__48887\,
            I => n2810
        );

    \I__10935\ : InMux
    port map (
            O => \N__48880\,
            I => \N__48877\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__48877\,
            I => \N__48874\
        );

    \I__10933\ : Span4Mux_h
    port map (
            O => \N__48874\,
            I => \N__48871\
        );

    \I__10932\ : Odrv4
    port map (
            O => \N__48871\,
            I => n2877
        );

    \I__10931\ : InMux
    port map (
            O => \N__48868\,
            I => \bfn_15_23_0_\
        );

    \I__10930\ : InMux
    port map (
            O => \N__48865\,
            I => \N__48860\
        );

    \I__10929\ : InMux
    port map (
            O => \N__48864\,
            I => \N__48857\
        );

    \I__10928\ : CascadeMux
    port map (
            O => \N__48863\,
            I => \N__48854\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__48860\,
            I => \N__48851\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__48857\,
            I => \N__48848\
        );

    \I__10925\ : InMux
    port map (
            O => \N__48854\,
            I => \N__48845\
        );

    \I__10924\ : Span4Mux_h
    port map (
            O => \N__48851\,
            I => \N__48842\
        );

    \I__10923\ : Span4Mux_h
    port map (
            O => \N__48848\,
            I => \N__48839\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__48845\,
            I => \N__48836\
        );

    \I__10921\ : Span4Mux_h
    port map (
            O => \N__48842\,
            I => \N__48833\
        );

    \I__10920\ : Span4Mux_h
    port map (
            O => \N__48839\,
            I => \N__48830\
        );

    \I__10919\ : Odrv4
    port map (
            O => \N__48836\,
            I => n2809
        );

    \I__10918\ : Odrv4
    port map (
            O => \N__48833\,
            I => n2809
        );

    \I__10917\ : Odrv4
    port map (
            O => \N__48830\,
            I => n2809
        );

    \I__10916\ : InMux
    port map (
            O => \N__48823\,
            I => \N__48820\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__48820\,
            I => \N__48817\
        );

    \I__10914\ : Span4Mux_v
    port map (
            O => \N__48817\,
            I => \N__48814\
        );

    \I__10913\ : Odrv4
    port map (
            O => \N__48814\,
            I => n2876
        );

    \I__10912\ : InMux
    port map (
            O => \N__48811\,
            I => n12435
        );

    \I__10911\ : InMux
    port map (
            O => \N__48808\,
            I => n12436
        );

    \I__10910\ : CascadeMux
    port map (
            O => \N__48805\,
            I => \N__48801\
        );

    \I__10909\ : InMux
    port map (
            O => \N__48804\,
            I => \N__48795\
        );

    \I__10908\ : InMux
    port map (
            O => \N__48801\,
            I => \N__48795\
        );

    \I__10907\ : InMux
    port map (
            O => \N__48800\,
            I => \N__48792\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__48795\,
            I => \N__48789\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__48792\,
            I => \N__48786\
        );

    \I__10904\ : Span4Mux_v
    port map (
            O => \N__48789\,
            I => \N__48783\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__48786\,
            I => \N__48780\
        );

    \I__10902\ : Odrv4
    port map (
            O => \N__48783\,
            I => n2808
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__48780\,
            I => n2808
        );

    \I__10900\ : CascadeMux
    port map (
            O => \N__48775\,
            I => \N__48772\
        );

    \I__10899\ : InMux
    port map (
            O => \N__48772\,
            I => \N__48769\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__48769\,
            I => n2875
        );

    \I__10897\ : CascadeMux
    port map (
            O => \N__48766\,
            I => \N__48763\
        );

    \I__10896\ : InMux
    port map (
            O => \N__48763\,
            I => \N__48760\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__48760\,
            I => \N__48756\
        );

    \I__10894\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48753\
        );

    \I__10893\ : Span4Mux_v
    port map (
            O => \N__48756\,
            I => \N__48748\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__48753\,
            I => \N__48748\
        );

    \I__10891\ : Span4Mux_h
    port map (
            O => \N__48748\,
            I => \N__48745\
        );

    \I__10890\ : Odrv4
    port map (
            O => \N__48745\,
            I => n2907
        );

    \I__10889\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48738\
        );

    \I__10888\ : InMux
    port map (
            O => \N__48741\,
            I => \N__48735\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__48738\,
            I => \N__48729\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__48735\,
            I => \N__48729\
        );

    \I__10885\ : InMux
    port map (
            O => \N__48734\,
            I => \N__48726\
        );

    \I__10884\ : Span4Mux_v
    port map (
            O => \N__48729\,
            I => \N__48723\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__48726\,
            I => n3220
        );

    \I__10882\ : Odrv4
    port map (
            O => \N__48723\,
            I => n3220
        );

    \I__10881\ : CascadeMux
    port map (
            O => \N__48718\,
            I => \N__48715\
        );

    \I__10880\ : InMux
    port map (
            O => \N__48715\,
            I => \N__48712\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__48712\,
            I => \N__48709\
        );

    \I__10878\ : Odrv12
    port map (
            O => \N__48709\,
            I => n3287
        );

    \I__10877\ : InMux
    port map (
            O => \N__48706\,
            I => \N__48703\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__48703\,
            I => n17_adj_705
        );

    \I__10875\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48697\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__48697\,
            I => \N__48694\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__48694\,
            I => \N__48691\
        );

    \I__10872\ : Span4Mux_h
    port map (
            O => \N__48691\,
            I => \N__48688\
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__48688\,
            I => n3296
        );

    \I__10870\ : CascadeMux
    port map (
            O => \N__48685\,
            I => \n13822_cascade_\
        );

    \I__10869\ : InMux
    port map (
            O => \N__48682\,
            I => \N__48678\
        );

    \I__10868\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48675\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48672\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__48675\,
            I => \N__48669\
        );

    \I__10865\ : Span4Mux_h
    port map (
            O => \N__48672\,
            I => \N__48666\
        );

    \I__10864\ : Odrv12
    port map (
            O => \N__48669\,
            I => n3229
        );

    \I__10863\ : Odrv4
    port map (
            O => \N__48666\,
            I => n3229
        );

    \I__10862\ : InMux
    port map (
            O => \N__48661\,
            I => \N__48658\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__48658\,
            I => n15_adj_704
        );

    \I__10860\ : CascadeMux
    port map (
            O => \N__48655\,
            I => \n13834_cascade_\
        );

    \I__10859\ : InMux
    port map (
            O => \N__48652\,
            I => \N__48649\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__48649\,
            I => \N__48646\
        );

    \I__10857\ : Odrv4
    port map (
            O => \N__48646\,
            I => n13842
        );

    \I__10856\ : InMux
    port map (
            O => \N__48643\,
            I => \N__48640\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__48640\,
            I => \N__48636\
        );

    \I__10854\ : InMux
    port map (
            O => \N__48639\,
            I => \N__48632\
        );

    \I__10853\ : Span4Mux_h
    port map (
            O => \N__48636\,
            I => \N__48629\
        );

    \I__10852\ : InMux
    port map (
            O => \N__48635\,
            I => \N__48626\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__48632\,
            I => \N__48623\
        );

    \I__10850\ : Odrv4
    port map (
            O => \N__48629\,
            I => n3222
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__48626\,
            I => n3222
        );

    \I__10848\ : Odrv12
    port map (
            O => \N__48623\,
            I => n3222
        );

    \I__10847\ : CascadeMux
    port map (
            O => \N__48616\,
            I => \N__48613\
        );

    \I__10846\ : InMux
    port map (
            O => \N__48613\,
            I => \N__48610\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__48610\,
            I => \N__48607\
        );

    \I__10844\ : Odrv4
    port map (
            O => \N__48607\,
            I => n3289
        );

    \I__10843\ : InMux
    port map (
            O => \N__48604\,
            I => \N__48601\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__48601\,
            I => \N__48598\
        );

    \I__10841\ : Span4Mux_h
    port map (
            O => \N__48598\,
            I => \N__48595\
        );

    \I__10840\ : Odrv4
    port map (
            O => \N__48595\,
            I => n2885
        );

    \I__10839\ : InMux
    port map (
            O => \N__48592\,
            I => \bfn_15_22_0_\
        );

    \I__10838\ : InMux
    port map (
            O => \N__48589\,
            I => \N__48586\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__48586\,
            I => \N__48582\
        );

    \I__10836\ : InMux
    port map (
            O => \N__48585\,
            I => \N__48579\
        );

    \I__10835\ : Span4Mux_v
    port map (
            O => \N__48582\,
            I => \N__48574\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__48579\,
            I => \N__48574\
        );

    \I__10833\ : Span4Mux_h
    port map (
            O => \N__48574\,
            I => \N__48571\
        );

    \I__10832\ : Odrv4
    port map (
            O => \N__48571\,
            I => n2817
        );

    \I__10831\ : InMux
    port map (
            O => \N__48568\,
            I => \N__48565\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__48565\,
            I => \N__48562\
        );

    \I__10829\ : Span4Mux_h
    port map (
            O => \N__48562\,
            I => \N__48559\
        );

    \I__10828\ : Odrv4
    port map (
            O => \N__48559\,
            I => n2884
        );

    \I__10827\ : InMux
    port map (
            O => \N__48556\,
            I => n12427
        );

    \I__10826\ : InMux
    port map (
            O => \N__48553\,
            I => \N__48549\
        );

    \I__10825\ : InMux
    port map (
            O => \N__48552\,
            I => \N__48546\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__48549\,
            I => \N__48542\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__48546\,
            I => \N__48539\
        );

    \I__10822\ : InMux
    port map (
            O => \N__48545\,
            I => \N__48536\
        );

    \I__10821\ : Span4Mux_h
    port map (
            O => \N__48542\,
            I => \N__48533\
        );

    \I__10820\ : Span4Mux_v
    port map (
            O => \N__48539\,
            I => \N__48528\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__48536\,
            I => \N__48528\
        );

    \I__10818\ : Odrv4
    port map (
            O => \N__48533\,
            I => n2816
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__48528\,
            I => n2816
        );

    \I__10816\ : CascadeMux
    port map (
            O => \N__48523\,
            I => \N__48520\
        );

    \I__10815\ : InMux
    port map (
            O => \N__48520\,
            I => \N__48517\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__48517\,
            I => \N__48514\
        );

    \I__10813\ : Span4Mux_h
    port map (
            O => \N__48514\,
            I => \N__48511\
        );

    \I__10812\ : Odrv4
    port map (
            O => \N__48511\,
            I => n2883
        );

    \I__10811\ : InMux
    port map (
            O => \N__48508\,
            I => n12428
        );

    \I__10810\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48501\
        );

    \I__10809\ : InMux
    port map (
            O => \N__48504\,
            I => \N__48498\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__48501\,
            I => \N__48495\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__48498\,
            I => \N__48489\
        );

    \I__10806\ : Span4Mux_v
    port map (
            O => \N__48495\,
            I => \N__48489\
        );

    \I__10805\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48486\
        );

    \I__10804\ : Odrv4
    port map (
            O => \N__48489\,
            I => n2815
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__48486\,
            I => n2815
        );

    \I__10802\ : InMux
    port map (
            O => \N__48481\,
            I => \N__48478\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__48478\,
            I => \N__48475\
        );

    \I__10800\ : Odrv4
    port map (
            O => \N__48475\,
            I => n2882
        );

    \I__10799\ : InMux
    port map (
            O => \N__48472\,
            I => n12429
        );

    \I__10798\ : CascadeMux
    port map (
            O => \N__48469\,
            I => \N__48466\
        );

    \I__10797\ : InMux
    port map (
            O => \N__48466\,
            I => \N__48462\
        );

    \I__10796\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48459\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__48462\,
            I => \N__48456\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__48459\,
            I => \N__48453\
        );

    \I__10793\ : Span4Mux_v
    port map (
            O => \N__48456\,
            I => \N__48450\
        );

    \I__10792\ : Span4Mux_v
    port map (
            O => \N__48453\,
            I => \N__48447\
        );

    \I__10791\ : Odrv4
    port map (
            O => \N__48450\,
            I => n2814
        );

    \I__10790\ : Odrv4
    port map (
            O => \N__48447\,
            I => n2814
        );

    \I__10789\ : InMux
    port map (
            O => \N__48442\,
            I => \N__48439\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__48439\,
            I => \N__48436\
        );

    \I__10787\ : Odrv4
    port map (
            O => \N__48436\,
            I => n2881
        );

    \I__10786\ : InMux
    port map (
            O => \N__48433\,
            I => n12430
        );

    \I__10785\ : InMux
    port map (
            O => \N__48430\,
            I => \N__48426\
        );

    \I__10784\ : InMux
    port map (
            O => \N__48429\,
            I => \N__48422\
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__48426\,
            I => \N__48419\
        );

    \I__10782\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48416\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__48422\,
            I => \N__48413\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__48419\,
            I => \N__48410\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__48416\,
            I => \N__48407\
        );

    \I__10778\ : Span4Mux_v
    port map (
            O => \N__48413\,
            I => \N__48400\
        );

    \I__10777\ : Span4Mux_h
    port map (
            O => \N__48410\,
            I => \N__48400\
        );

    \I__10776\ : Span4Mux_h
    port map (
            O => \N__48407\,
            I => \N__48400\
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__48400\,
            I => n2813
        );

    \I__10774\ : InMux
    port map (
            O => \N__48397\,
            I => \N__48394\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__48394\,
            I => \N__48391\
        );

    \I__10772\ : Odrv12
    port map (
            O => \N__48391\,
            I => n2880
        );

    \I__10771\ : InMux
    port map (
            O => \N__48388\,
            I => n12431
        );

    \I__10770\ : InMux
    port map (
            O => \N__48385\,
            I => \N__48381\
        );

    \I__10769\ : InMux
    port map (
            O => \N__48384\,
            I => \N__48378\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__48381\,
            I => \N__48374\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__48378\,
            I => \N__48371\
        );

    \I__10766\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48368\
        );

    \I__10765\ : Span4Mux_h
    port map (
            O => \N__48374\,
            I => \N__48365\
        );

    \I__10764\ : Span4Mux_h
    port map (
            O => \N__48371\,
            I => \N__48362\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__48368\,
            I => n2812
        );

    \I__10762\ : Odrv4
    port map (
            O => \N__48365\,
            I => n2812
        );

    \I__10761\ : Odrv4
    port map (
            O => \N__48362\,
            I => n2812
        );

    \I__10760\ : CascadeMux
    port map (
            O => \N__48355\,
            I => \N__48352\
        );

    \I__10759\ : InMux
    port map (
            O => \N__48352\,
            I => \N__48349\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__48349\,
            I => \N__48346\
        );

    \I__10757\ : Span4Mux_h
    port map (
            O => \N__48346\,
            I => \N__48343\
        );

    \I__10756\ : Odrv4
    port map (
            O => \N__48343\,
            I => n2879
        );

    \I__10755\ : InMux
    port map (
            O => \N__48340\,
            I => n12432
        );

    \I__10754\ : InMux
    port map (
            O => \N__48337\,
            I => \N__48333\
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__48336\,
            I => \N__48330\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__48333\,
            I => \N__48327\
        );

    \I__10751\ : InMux
    port map (
            O => \N__48330\,
            I => \N__48324\
        );

    \I__10750\ : Span4Mux_v
    port map (
            O => \N__48327\,
            I => \N__48321\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__48324\,
            I => n2811
        );

    \I__10748\ : Odrv4
    port map (
            O => \N__48321\,
            I => n2811
        );

    \I__10747\ : InMux
    port map (
            O => \N__48316\,
            I => \N__48313\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__48313\,
            I => \N__48310\
        );

    \I__10745\ : Odrv12
    port map (
            O => \N__48310\,
            I => n2878
        );

    \I__10744\ : InMux
    port map (
            O => \N__48307\,
            I => n12433
        );

    \I__10743\ : CascadeMux
    port map (
            O => \N__48304\,
            I => \N__48300\
        );

    \I__10742\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48297\
        );

    \I__10741\ : InMux
    port map (
            O => \N__48300\,
            I => \N__48294\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__48297\,
            I => \N__48291\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__48294\,
            I => n2825
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__48291\,
            I => n2825
        );

    \I__10737\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48283\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__48283\,
            I => n2892
        );

    \I__10735\ : InMux
    port map (
            O => \N__48280\,
            I => n12419
        );

    \I__10734\ : CascadeMux
    port map (
            O => \N__48277\,
            I => \N__48274\
        );

    \I__10733\ : InMux
    port map (
            O => \N__48274\,
            I => \N__48270\
        );

    \I__10732\ : InMux
    port map (
            O => \N__48273\,
            I => \N__48267\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__48270\,
            I => \N__48264\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__48267\,
            I => \N__48260\
        );

    \I__10729\ : Span4Mux_v
    port map (
            O => \N__48264\,
            I => \N__48257\
        );

    \I__10728\ : InMux
    port map (
            O => \N__48263\,
            I => \N__48254\
        );

    \I__10727\ : Odrv4
    port map (
            O => \N__48260\,
            I => n2824
        );

    \I__10726\ : Odrv4
    port map (
            O => \N__48257\,
            I => n2824
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__48254\,
            I => n2824
        );

    \I__10724\ : InMux
    port map (
            O => \N__48247\,
            I => \N__48244\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__48244\,
            I => \N__48241\
        );

    \I__10722\ : Odrv4
    port map (
            O => \N__48241\,
            I => n2891
        );

    \I__10721\ : InMux
    port map (
            O => \N__48238\,
            I => n12420
        );

    \I__10720\ : CascadeMux
    port map (
            O => \N__48235\,
            I => \N__48231\
        );

    \I__10719\ : CascadeMux
    port map (
            O => \N__48234\,
            I => \N__48228\
        );

    \I__10718\ : InMux
    port map (
            O => \N__48231\,
            I => \N__48225\
        );

    \I__10717\ : InMux
    port map (
            O => \N__48228\,
            I => \N__48221\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__48225\,
            I => \N__48218\
        );

    \I__10715\ : CascadeMux
    port map (
            O => \N__48224\,
            I => \N__48215\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__48221\,
            I => \N__48210\
        );

    \I__10713\ : Span4Mux_h
    port map (
            O => \N__48218\,
            I => \N__48210\
        );

    \I__10712\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48207\
        );

    \I__10711\ : Odrv4
    port map (
            O => \N__48210\,
            I => n2823
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__48207\,
            I => n2823
        );

    \I__10709\ : InMux
    port map (
            O => \N__48202\,
            I => \N__48199\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__48199\,
            I => \N__48196\
        );

    \I__10707\ : Odrv4
    port map (
            O => \N__48196\,
            I => n2890
        );

    \I__10706\ : InMux
    port map (
            O => \N__48193\,
            I => n12421
        );

    \I__10705\ : CascadeMux
    port map (
            O => \N__48190\,
            I => \N__48187\
        );

    \I__10704\ : InMux
    port map (
            O => \N__48187\,
            I => \N__48183\
        );

    \I__10703\ : InMux
    port map (
            O => \N__48186\,
            I => \N__48180\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__48183\,
            I => \N__48177\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__48180\,
            I => \N__48173\
        );

    \I__10700\ : Span4Mux_v
    port map (
            O => \N__48177\,
            I => \N__48170\
        );

    \I__10699\ : InMux
    port map (
            O => \N__48176\,
            I => \N__48167\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__48173\,
            I => n2822
        );

    \I__10697\ : Odrv4
    port map (
            O => \N__48170\,
            I => n2822
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__48167\,
            I => n2822
        );

    \I__10695\ : CascadeMux
    port map (
            O => \N__48160\,
            I => \N__48157\
        );

    \I__10694\ : InMux
    port map (
            O => \N__48157\,
            I => \N__48154\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__48154\,
            I => \N__48151\
        );

    \I__10692\ : Span4Mux_h
    port map (
            O => \N__48151\,
            I => \N__48148\
        );

    \I__10691\ : Odrv4
    port map (
            O => \N__48148\,
            I => n2889
        );

    \I__10690\ : InMux
    port map (
            O => \N__48145\,
            I => n12422
        );

    \I__10689\ : CascadeMux
    port map (
            O => \N__48142\,
            I => \N__48139\
        );

    \I__10688\ : InMux
    port map (
            O => \N__48139\,
            I => \N__48135\
        );

    \I__10687\ : CascadeMux
    port map (
            O => \N__48138\,
            I => \N__48132\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__48135\,
            I => \N__48129\
        );

    \I__10685\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48125\
        );

    \I__10684\ : Span4Mux_h
    port map (
            O => \N__48129\,
            I => \N__48122\
        );

    \I__10683\ : InMux
    port map (
            O => \N__48128\,
            I => \N__48119\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__48125\,
            I => n2821
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__48122\,
            I => n2821
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__48119\,
            I => n2821
        );

    \I__10679\ : InMux
    port map (
            O => \N__48112\,
            I => \N__48109\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__48109\,
            I => \N__48106\
        );

    \I__10677\ : Odrv4
    port map (
            O => \N__48106\,
            I => n2888
        );

    \I__10676\ : InMux
    port map (
            O => \N__48103\,
            I => n12423
        );

    \I__10675\ : CascadeMux
    port map (
            O => \N__48100\,
            I => \N__48096\
        );

    \I__10674\ : CascadeMux
    port map (
            O => \N__48099\,
            I => \N__48093\
        );

    \I__10673\ : InMux
    port map (
            O => \N__48096\,
            I => \N__48090\
        );

    \I__10672\ : InMux
    port map (
            O => \N__48093\,
            I => \N__48087\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__48090\,
            I => \N__48084\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__48087\,
            I => \N__48081\
        );

    \I__10669\ : Span4Mux_v
    port map (
            O => \N__48084\,
            I => \N__48077\
        );

    \I__10668\ : Span4Mux_v
    port map (
            O => \N__48081\,
            I => \N__48074\
        );

    \I__10667\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48071\
        );

    \I__10666\ : Sp12to4
    port map (
            O => \N__48077\,
            I => \N__48064\
        );

    \I__10665\ : Sp12to4
    port map (
            O => \N__48074\,
            I => \N__48064\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__48071\,
            I => \N__48064\
        );

    \I__10663\ : Odrv12
    port map (
            O => \N__48064\,
            I => n2820
        );

    \I__10662\ : InMux
    port map (
            O => \N__48061\,
            I => \N__48058\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__48058\,
            I => \N__48055\
        );

    \I__10660\ : Odrv4
    port map (
            O => \N__48055\,
            I => n2887
        );

    \I__10659\ : InMux
    port map (
            O => \N__48052\,
            I => n12424
        );

    \I__10658\ : CascadeMux
    port map (
            O => \N__48049\,
            I => \N__48046\
        );

    \I__10657\ : InMux
    port map (
            O => \N__48046\,
            I => \N__48043\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__48043\,
            I => \N__48039\
        );

    \I__10655\ : InMux
    port map (
            O => \N__48042\,
            I => \N__48035\
        );

    \I__10654\ : Span4Mux_h
    port map (
            O => \N__48039\,
            I => \N__48032\
        );

    \I__10653\ : InMux
    port map (
            O => \N__48038\,
            I => \N__48029\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__48035\,
            I => n2819
        );

    \I__10651\ : Odrv4
    port map (
            O => \N__48032\,
            I => n2819
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__48029\,
            I => n2819
        );

    \I__10649\ : InMux
    port map (
            O => \N__48022\,
            I => \N__48019\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__48019\,
            I => \N__48016\
        );

    \I__10647\ : Span4Mux_h
    port map (
            O => \N__48016\,
            I => \N__48013\
        );

    \I__10646\ : Odrv4
    port map (
            O => \N__48013\,
            I => n2886
        );

    \I__10645\ : InMux
    port map (
            O => \N__48010\,
            I => n12425
        );

    \I__10644\ : InMux
    port map (
            O => \N__48007\,
            I => \N__48004\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__48004\,
            I => \N__48000\
        );

    \I__10642\ : InMux
    port map (
            O => \N__48003\,
            I => \N__47996\
        );

    \I__10641\ : Span4Mux_v
    port map (
            O => \N__48000\,
            I => \N__47993\
        );

    \I__10640\ : InMux
    port map (
            O => \N__47999\,
            I => \N__47990\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__47996\,
            I => n2818
        );

    \I__10638\ : Odrv4
    port map (
            O => \N__47993\,
            I => n2818
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__47990\,
            I => n2818
        );

    \I__10636\ : CascadeMux
    port map (
            O => \N__47983\,
            I => \N__47979\
        );

    \I__10635\ : InMux
    port map (
            O => \N__47982\,
            I => \N__47976\
        );

    \I__10634\ : InMux
    port map (
            O => \N__47979\,
            I => \N__47973\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__47976\,
            I => n2833
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__47973\,
            I => n2833
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__47968\,
            I => \N__47965\
        );

    \I__10630\ : InMux
    port map (
            O => \N__47965\,
            I => \N__47962\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__47962\,
            I => n2900
        );

    \I__10628\ : InMux
    port map (
            O => \N__47959\,
            I => n12411
        );

    \I__10627\ : CascadeMux
    port map (
            O => \N__47956\,
            I => \N__47953\
        );

    \I__10626\ : InMux
    port map (
            O => \N__47953\,
            I => \N__47948\
        );

    \I__10625\ : InMux
    port map (
            O => \N__47952\,
            I => \N__47943\
        );

    \I__10624\ : InMux
    port map (
            O => \N__47951\,
            I => \N__47943\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__47948\,
            I => \N__47940\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__47943\,
            I => n2832
        );

    \I__10621\ : Odrv4
    port map (
            O => \N__47940\,
            I => n2832
        );

    \I__10620\ : InMux
    port map (
            O => \N__47935\,
            I => \N__47932\
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__47932\,
            I => n2899
        );

    \I__10618\ : InMux
    port map (
            O => \N__47929\,
            I => n12412
        );

    \I__10617\ : CascadeMux
    port map (
            O => \N__47926\,
            I => \N__47923\
        );

    \I__10616\ : InMux
    port map (
            O => \N__47923\,
            I => \N__47918\
        );

    \I__10615\ : InMux
    port map (
            O => \N__47922\,
            I => \N__47913\
        );

    \I__10614\ : InMux
    port map (
            O => \N__47921\,
            I => \N__47913\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__47918\,
            I => \N__47910\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__47913\,
            I => n2831
        );

    \I__10611\ : Odrv4
    port map (
            O => \N__47910\,
            I => n2831
        );

    \I__10610\ : CascadeMux
    port map (
            O => \N__47905\,
            I => \N__47902\
        );

    \I__10609\ : InMux
    port map (
            O => \N__47902\,
            I => \N__47899\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__47899\,
            I => n2898
        );

    \I__10607\ : InMux
    port map (
            O => \N__47896\,
            I => n12413
        );

    \I__10606\ : CascadeMux
    port map (
            O => \N__47893\,
            I => \N__47890\
        );

    \I__10605\ : InMux
    port map (
            O => \N__47890\,
            I => \N__47886\
        );

    \I__10604\ : CascadeMux
    port map (
            O => \N__47889\,
            I => \N__47883\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__47886\,
            I => \N__47879\
        );

    \I__10602\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47874\
        );

    \I__10601\ : InMux
    port map (
            O => \N__47882\,
            I => \N__47874\
        );

    \I__10600\ : Span4Mux_h
    port map (
            O => \N__47879\,
            I => \N__47871\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__47874\,
            I => n2830
        );

    \I__10598\ : Odrv4
    port map (
            O => \N__47871\,
            I => n2830
        );

    \I__10597\ : InMux
    port map (
            O => \N__47866\,
            I => \N__47863\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__47863\,
            I => \N__47860\
        );

    \I__10595\ : Odrv4
    port map (
            O => \N__47860\,
            I => n2897
        );

    \I__10594\ : InMux
    port map (
            O => \N__47857\,
            I => n12414
        );

    \I__10593\ : CascadeMux
    port map (
            O => \N__47854\,
            I => \N__47851\
        );

    \I__10592\ : InMux
    port map (
            O => \N__47851\,
            I => \N__47847\
        );

    \I__10591\ : CascadeMux
    port map (
            O => \N__47850\,
            I => \N__47843\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__47847\,
            I => \N__47840\
        );

    \I__10589\ : InMux
    port map (
            O => \N__47846\,
            I => \N__47837\
        );

    \I__10588\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47834\
        );

    \I__10587\ : Span4Mux_h
    port map (
            O => \N__47840\,
            I => \N__47831\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__47837\,
            I => n2829
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__47834\,
            I => n2829
        );

    \I__10584\ : Odrv4
    port map (
            O => \N__47831\,
            I => n2829
        );

    \I__10583\ : InMux
    port map (
            O => \N__47824\,
            I => \N__47821\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__47821\,
            I => n2896
        );

    \I__10581\ : InMux
    port map (
            O => \N__47818\,
            I => n12415
        );

    \I__10580\ : CascadeMux
    port map (
            O => \N__47815\,
            I => \N__47811\
        );

    \I__10579\ : InMux
    port map (
            O => \N__47814\,
            I => \N__47807\
        );

    \I__10578\ : InMux
    port map (
            O => \N__47811\,
            I => \N__47804\
        );

    \I__10577\ : InMux
    port map (
            O => \N__47810\,
            I => \N__47801\
        );

    \I__10576\ : LocalMux
    port map (
            O => \N__47807\,
            I => \N__47796\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__47804\,
            I => \N__47796\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__47801\,
            I => n2828
        );

    \I__10573\ : Odrv4
    port map (
            O => \N__47796\,
            I => n2828
        );

    \I__10572\ : InMux
    port map (
            O => \N__47791\,
            I => \N__47788\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__47788\,
            I => n2895
        );

    \I__10570\ : InMux
    port map (
            O => \N__47785\,
            I => n12416
        );

    \I__10569\ : CascadeMux
    port map (
            O => \N__47782\,
            I => \N__47778\
        );

    \I__10568\ : CascadeMux
    port map (
            O => \N__47781\,
            I => \N__47775\
        );

    \I__10567\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47772\
        );

    \I__10566\ : InMux
    port map (
            O => \N__47775\,
            I => \N__47769\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__47772\,
            I => \N__47766\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__47769\,
            I => \N__47763\
        );

    \I__10563\ : Span4Mux_h
    port map (
            O => \N__47766\,
            I => \N__47759\
        );

    \I__10562\ : Span4Mux_h
    port map (
            O => \N__47763\,
            I => \N__47756\
        );

    \I__10561\ : InMux
    port map (
            O => \N__47762\,
            I => \N__47753\
        );

    \I__10560\ : Odrv4
    port map (
            O => \N__47759\,
            I => n2827
        );

    \I__10559\ : Odrv4
    port map (
            O => \N__47756\,
            I => n2827
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__47753\,
            I => n2827
        );

    \I__10557\ : InMux
    port map (
            O => \N__47746\,
            I => \N__47743\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__47743\,
            I => n2894
        );

    \I__10555\ : InMux
    port map (
            O => \N__47740\,
            I => n12417
        );

    \I__10554\ : CascadeMux
    port map (
            O => \N__47737\,
            I => \N__47733\
        );

    \I__10553\ : InMux
    port map (
            O => \N__47736\,
            I => \N__47730\
        );

    \I__10552\ : InMux
    port map (
            O => \N__47733\,
            I => \N__47727\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__47730\,
            I => \N__47721\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__47727\,
            I => \N__47721\
        );

    \I__10549\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47718\
        );

    \I__10548\ : Span4Mux_v
    port map (
            O => \N__47721\,
            I => \N__47715\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__47718\,
            I => \N__47712\
        );

    \I__10546\ : Odrv4
    port map (
            O => \N__47715\,
            I => n2826
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__47712\,
            I => n2826
        );

    \I__10544\ : CascadeMux
    port map (
            O => \N__47707\,
            I => \N__47704\
        );

    \I__10543\ : InMux
    port map (
            O => \N__47704\,
            I => \N__47701\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__47701\,
            I => n2893
        );

    \I__10541\ : InMux
    port map (
            O => \N__47698\,
            I => \bfn_15_21_0_\
        );

    \I__10540\ : InMux
    port map (
            O => \N__47695\,
            I => \N__47692\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__47692\,
            I => \N__47689\
        );

    \I__10538\ : Span4Mux_h
    port map (
            O => \N__47689\,
            I => \N__47686\
        );

    \I__10537\ : Odrv4
    port map (
            O => \N__47686\,
            I => n2801
        );

    \I__10536\ : InMux
    port map (
            O => \N__47683\,
            I => \N__47679\
        );

    \I__10535\ : InMux
    port map (
            O => \N__47682\,
            I => \N__47675\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__47679\,
            I => \N__47672\
        );

    \I__10533\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47669\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__47675\,
            I => \N__47666\
        );

    \I__10531\ : Span4Mux_v
    port map (
            O => \N__47672\,
            I => \N__47661\
        );

    \I__10530\ : LocalMux
    port map (
            O => \N__47669\,
            I => \N__47661\
        );

    \I__10529\ : Span4Mux_h
    port map (
            O => \N__47666\,
            I => \N__47658\
        );

    \I__10528\ : Span4Mux_h
    port map (
            O => \N__47661\,
            I => \N__47655\
        );

    \I__10527\ : Span4Mux_h
    port map (
            O => \N__47658\,
            I => \N__47652\
        );

    \I__10526\ : Span4Mux_v
    port map (
            O => \N__47655\,
            I => \N__47649\
        );

    \I__10525\ : Odrv4
    port map (
            O => \N__47652\,
            I => n313
        );

    \I__10524\ : Odrv4
    port map (
            O => \N__47649\,
            I => n313
        );

    \I__10523\ : CascadeMux
    port map (
            O => \N__47644\,
            I => \N__47641\
        );

    \I__10522\ : InMux
    port map (
            O => \N__47641\,
            I => \N__47638\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__47638\,
            I => \N__47634\
        );

    \I__10520\ : InMux
    port map (
            O => \N__47637\,
            I => \N__47631\
        );

    \I__10519\ : Span4Mux_v
    port map (
            O => \N__47634\,
            I => \N__47620\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__47631\,
            I => \N__47620\
        );

    \I__10517\ : InMux
    port map (
            O => \N__47630\,
            I => \N__47617\
        );

    \I__10516\ : InMux
    port map (
            O => \N__47629\,
            I => \N__47613\
        );

    \I__10515\ : InMux
    port map (
            O => \N__47628\,
            I => \N__47608\
        );

    \I__10514\ : InMux
    port map (
            O => \N__47627\,
            I => \N__47608\
        );

    \I__10513\ : CascadeMux
    port map (
            O => \N__47626\,
            I => \N__47599\
        );

    \I__10512\ : CascadeMux
    port map (
            O => \N__47625\,
            I => \N__47596\
        );

    \I__10511\ : Span4Mux_v
    port map (
            O => \N__47620\,
            I => \N__47589\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__47617\,
            I => \N__47589\
        );

    \I__10509\ : InMux
    port map (
            O => \N__47616\,
            I => \N__47586\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__47613\,
            I => \N__47581\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__47608\,
            I => \N__47581\
        );

    \I__10506\ : CascadeMux
    port map (
            O => \N__47607\,
            I => \N__47578\
        );

    \I__10505\ : CascadeMux
    port map (
            O => \N__47606\,
            I => \N__47574\
        );

    \I__10504\ : CascadeMux
    port map (
            O => \N__47605\,
            I => \N__47569\
        );

    \I__10503\ : CascadeMux
    port map (
            O => \N__47604\,
            I => \N__47564\
        );

    \I__10502\ : CascadeMux
    port map (
            O => \N__47603\,
            I => \N__47559\
        );

    \I__10501\ : CascadeMux
    port map (
            O => \N__47602\,
            I => \N__47555\
        );

    \I__10500\ : InMux
    port map (
            O => \N__47599\,
            I => \N__47549\
        );

    \I__10499\ : InMux
    port map (
            O => \N__47596\,
            I => \N__47549\
        );

    \I__10498\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47546\
        );

    \I__10497\ : InMux
    port map (
            O => \N__47594\,
            I => \N__47543\
        );

    \I__10496\ : Span4Mux_v
    port map (
            O => \N__47589\,
            I => \N__47540\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__47586\,
            I => \N__47537\
        );

    \I__10494\ : Span4Mux_v
    port map (
            O => \N__47581\,
            I => \N__47534\
        );

    \I__10493\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47523\
        );

    \I__10492\ : InMux
    port map (
            O => \N__47577\,
            I => \N__47523\
        );

    \I__10491\ : InMux
    port map (
            O => \N__47574\,
            I => \N__47523\
        );

    \I__10490\ : InMux
    port map (
            O => \N__47573\,
            I => \N__47523\
        );

    \I__10489\ : InMux
    port map (
            O => \N__47572\,
            I => \N__47523\
        );

    \I__10488\ : InMux
    port map (
            O => \N__47569\,
            I => \N__47516\
        );

    \I__10487\ : InMux
    port map (
            O => \N__47568\,
            I => \N__47516\
        );

    \I__10486\ : InMux
    port map (
            O => \N__47567\,
            I => \N__47516\
        );

    \I__10485\ : InMux
    port map (
            O => \N__47564\,
            I => \N__47511\
        );

    \I__10484\ : InMux
    port map (
            O => \N__47563\,
            I => \N__47511\
        );

    \I__10483\ : InMux
    port map (
            O => \N__47562\,
            I => \N__47500\
        );

    \I__10482\ : InMux
    port map (
            O => \N__47559\,
            I => \N__47500\
        );

    \I__10481\ : InMux
    port map (
            O => \N__47558\,
            I => \N__47500\
        );

    \I__10480\ : InMux
    port map (
            O => \N__47555\,
            I => \N__47500\
        );

    \I__10479\ : InMux
    port map (
            O => \N__47554\,
            I => \N__47500\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__47549\,
            I => \N__47495\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__47546\,
            I => \N__47495\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__47543\,
            I => \N__47488\
        );

    \I__10475\ : Span4Mux_h
    port map (
            O => \N__47540\,
            I => \N__47488\
        );

    \I__10474\ : Span4Mux_h
    port map (
            O => \N__47537\,
            I => \N__47488\
        );

    \I__10473\ : Odrv4
    port map (
            O => \N__47534\,
            I => n2742
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__47523\,
            I => n2742
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__47516\,
            I => n2742
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__47511\,
            I => n2742
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__47500\,
            I => n2742
        );

    \I__10468\ : Odrv4
    port map (
            O => \N__47495\,
            I => n2742
        );

    \I__10467\ : Odrv4
    port map (
            O => \N__47488\,
            I => n2742
        );

    \I__10466\ : CascadeMux
    port map (
            O => \N__47473\,
            I => \n2833_cascade_\
        );

    \I__10465\ : InMux
    port map (
            O => \N__47470\,
            I => \N__47467\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__47467\,
            I => n11756
        );

    \I__10463\ : CascadeMux
    port map (
            O => \N__47464\,
            I => \N__47461\
        );

    \I__10462\ : InMux
    port map (
            O => \N__47461\,
            I => \N__47457\
        );

    \I__10461\ : InMux
    port map (
            O => \N__47460\,
            I => \N__47454\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__47457\,
            I => \N__47451\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__47454\,
            I => \N__47448\
        );

    \I__10458\ : Span4Mux_v
    port map (
            O => \N__47451\,
            I => \N__47445\
        );

    \I__10457\ : Span4Mux_v
    port map (
            O => \N__47448\,
            I => \N__47442\
        );

    \I__10456\ : Span4Mux_h
    port map (
            O => \N__47445\,
            I => \N__47439\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__47442\,
            I => n2932
        );

    \I__10454\ : Odrv4
    port map (
            O => \N__47439\,
            I => n2932
        );

    \I__10453\ : InMux
    port map (
            O => \N__47434\,
            I => \N__47431\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__47431\,
            I => \N__47427\
        );

    \I__10451\ : CascadeMux
    port map (
            O => \N__47430\,
            I => \N__47424\
        );

    \I__10450\ : Span4Mux_v
    port map (
            O => \N__47427\,
            I => \N__47421\
        );

    \I__10449\ : InMux
    port map (
            O => \N__47424\,
            I => \N__47418\
        );

    \I__10448\ : Span4Mux_h
    port map (
            O => \N__47421\,
            I => \N__47415\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__47418\,
            I => n315
        );

    \I__10446\ : Odrv4
    port map (
            O => \N__47415\,
            I => n315
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__47410\,
            I => \n2932_cascade_\
        );

    \I__10444\ : CascadeMux
    port map (
            O => \N__47407\,
            I => \N__47403\
        );

    \I__10443\ : InMux
    port map (
            O => \N__47406\,
            I => \N__47400\
        );

    \I__10442\ : InMux
    port map (
            O => \N__47403\,
            I => \N__47397\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__47400\,
            I => \N__47391\
        );

    \I__10440\ : LocalMux
    port map (
            O => \N__47397\,
            I => \N__47391\
        );

    \I__10439\ : InMux
    port map (
            O => \N__47396\,
            I => \N__47388\
        );

    \I__10438\ : Span4Mux_v
    port map (
            O => \N__47391\,
            I => \N__47385\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__47388\,
            I => \N__47382\
        );

    \I__10436\ : Odrv4
    port map (
            O => \N__47385\,
            I => n2933
        );

    \I__10435\ : Odrv4
    port map (
            O => \N__47382\,
            I => n2933
        );

    \I__10434\ : CascadeMux
    port map (
            O => \N__47377\,
            I => \N__47373\
        );

    \I__10433\ : InMux
    port map (
            O => \N__47376\,
            I => \N__47370\
        );

    \I__10432\ : InMux
    port map (
            O => \N__47373\,
            I => \N__47367\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__47370\,
            I => \N__47364\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__47367\,
            I => \N__47361\
        );

    \I__10429\ : Span4Mux_v
    port map (
            O => \N__47364\,
            I => \N__47356\
        );

    \I__10428\ : Span4Mux_h
    port map (
            O => \N__47361\,
            I => \N__47356\
        );

    \I__10427\ : Span4Mux_h
    port map (
            O => \N__47356\,
            I => \N__47353\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__47353\,
            I => n2930
        );

    \I__10425\ : CascadeMux
    port map (
            O => \N__47350\,
            I => \N__47347\
        );

    \I__10424\ : InMux
    port map (
            O => \N__47347\,
            I => \N__47343\
        );

    \I__10423\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47340\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__47343\,
            I => \N__47337\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__47340\,
            I => \N__47334\
        );

    \I__10420\ : Span4Mux_v
    port map (
            O => \N__47337\,
            I => \N__47330\
        );

    \I__10419\ : Span4Mux_v
    port map (
            O => \N__47334\,
            I => \N__47327\
        );

    \I__10418\ : InMux
    port map (
            O => \N__47333\,
            I => \N__47324\
        );

    \I__10417\ : Span4Mux_h
    port map (
            O => \N__47330\,
            I => \N__47321\
        );

    \I__10416\ : Odrv4
    port map (
            O => \N__47327\,
            I => n2931
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__47324\,
            I => n2931
        );

    \I__10414\ : Odrv4
    port map (
            O => \N__47321\,
            I => n2931
        );

    \I__10413\ : CascadeMux
    port map (
            O => \N__47314\,
            I => \N__47310\
        );

    \I__10412\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47307\
        );

    \I__10411\ : InMux
    port map (
            O => \N__47310\,
            I => \N__47304\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__47307\,
            I => \N__47300\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__47304\,
            I => \N__47297\
        );

    \I__10408\ : InMux
    port map (
            O => \N__47303\,
            I => \N__47294\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__47300\,
            I => \N__47289\
        );

    \I__10406\ : Span4Mux_h
    port map (
            O => \N__47297\,
            I => \N__47289\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__47294\,
            I => n2929
        );

    \I__10404\ : Odrv4
    port map (
            O => \N__47289\,
            I => n2929
        );

    \I__10403\ : CascadeMux
    port map (
            O => \N__47284\,
            I => \n2930_cascade_\
        );

    \I__10402\ : InMux
    port map (
            O => \N__47281\,
            I => \N__47278\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__47278\,
            I => n11662
        );

    \I__10400\ : CascadeMux
    port map (
            O => \N__47275\,
            I => \N__47272\
        );

    \I__10399\ : InMux
    port map (
            O => \N__47272\,
            I => \N__47269\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__47269\,
            I => \N__47266\
        );

    \I__10397\ : Span4Mux_h
    port map (
            O => \N__47266\,
            I => \N__47263\
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__47263\,
            I => n13417
        );

    \I__10395\ : InMux
    port map (
            O => \N__47260\,
            I => \N__47257\
        );

    \I__10394\ : LocalMux
    port map (
            O => \N__47257\,
            I => \N__47253\
        );

    \I__10393\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47250\
        );

    \I__10392\ : Span4Mux_v
    port map (
            O => \N__47253\,
            I => \N__47244\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__47250\,
            I => \N__47244\
        );

    \I__10390\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47241\
        );

    \I__10389\ : Span4Mux_h
    port map (
            O => \N__47244\,
            I => \N__47236\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__47241\,
            I => \N__47236\
        );

    \I__10387\ : Span4Mux_v
    port map (
            O => \N__47236\,
            I => \N__47233\
        );

    \I__10386\ : Span4Mux_h
    port map (
            O => \N__47233\,
            I => \N__47230\
        );

    \I__10385\ : Odrv4
    port map (
            O => \N__47230\,
            I => n314
        );

    \I__10384\ : InMux
    port map (
            O => \N__47227\,
            I => \N__47224\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__47224\,
            I => \N__47221\
        );

    \I__10382\ : Span4Mux_h
    port map (
            O => \N__47221\,
            I => \N__47218\
        );

    \I__10381\ : Odrv4
    port map (
            O => \N__47218\,
            I => n2901
        );

    \I__10380\ : InMux
    port map (
            O => \N__47215\,
            I => \bfn_15_20_0_\
        );

    \I__10379\ : InMux
    port map (
            O => \N__47212\,
            I => \N__47207\
        );

    \I__10378\ : InMux
    port map (
            O => \N__47211\,
            I => \N__47204\
        );

    \I__10377\ : InMux
    port map (
            O => \N__47210\,
            I => \N__47201\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__47207\,
            I => n31_adj_624
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__47204\,
            I => n31_adj_624
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__47201\,
            I => n31_adj_624
        );

    \I__10373\ : InMux
    port map (
            O => \N__47194\,
            I => \N__47191\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__47191\,
            I => \N__47188\
        );

    \I__10371\ : Span4Mux_s2_v
    port map (
            O => \N__47188\,
            I => \N__47185\
        );

    \I__10370\ : Odrv4
    port map (
            O => \N__47185\,
            I => n14728
        );

    \I__10369\ : CascadeMux
    port map (
            O => \N__47182\,
            I => \n33_adj_625_cascade_\
        );

    \I__10368\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47175\
        );

    \I__10367\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47172\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__47175\,
            I => \N__47166\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__47172\,
            I => \N__47166\
        );

    \I__10364\ : InMux
    port map (
            O => \N__47171\,
            I => \N__47163\
        );

    \I__10363\ : Odrv4
    port map (
            O => \N__47166\,
            I => n29_adj_622
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__47163\,
            I => n29_adj_622
        );

    \I__10361\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47155\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__47155\,
            I => n14724
        );

    \I__10359\ : InMux
    port map (
            O => \N__47152\,
            I => \N__47149\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__47149\,
            I => \N__47145\
        );

    \I__10357\ : InMux
    port map (
            O => \N__47148\,
            I => \N__47142\
        );

    \I__10356\ : Sp12to4
    port map (
            O => \N__47145\,
            I => \N__47137\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__47142\,
            I => \N__47137\
        );

    \I__10354\ : Odrv12
    port map (
            O => \N__47137\,
            I => duty_17
        );

    \I__10353\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47131\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__47131\,
            I => \N__47128\
        );

    \I__10351\ : Odrv4
    port map (
            O => \N__47128\,
            I => n8_adj_574
        );

    \I__10350\ : InMux
    port map (
            O => \N__47125\,
            I => \N__47122\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__47122\,
            I => n28_adj_597
        );

    \I__10348\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47116\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__47116\,
            I => n31_adj_594
        );

    \I__10346\ : CascadeMux
    port map (
            O => \N__47113\,
            I => \n32_adj_593_cascade_\
        );

    \I__10345\ : InMux
    port map (
            O => \N__47110\,
            I => \N__47107\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__47107\,
            I => \N__47104\
        );

    \I__10343\ : Span4Mux_v
    port map (
            O => \N__47104\,
            I => \N__47099\
        );

    \I__10342\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47094\
        );

    \I__10341\ : InMux
    port map (
            O => \N__47102\,
            I => \N__47094\
        );

    \I__10340\ : Span4Mux_h
    port map (
            O => \N__47099\,
            I => \N__47091\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__47094\,
            I => \N__47088\
        );

    \I__10338\ : Span4Mux_v
    port map (
            O => \N__47091\,
            I => \N__47085\
        );

    \I__10337\ : Span4Mux_h
    port map (
            O => \N__47088\,
            I => \N__47082\
        );

    \I__10336\ : Odrv4
    port map (
            O => \N__47085\,
            I => n2910
        );

    \I__10335\ : Odrv4
    port map (
            O => \N__47082\,
            I => n2910
        );

    \I__10334\ : InMux
    port map (
            O => \N__47077\,
            I => \N__47074\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__47074\,
            I => n30_adj_595
        );

    \I__10332\ : InMux
    port map (
            O => \N__47071\,
            I => \N__47068\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__47068\,
            I => n29_adj_596
        );

    \I__10330\ : InMux
    port map (
            O => \N__47065\,
            I => \N__47062\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__47062\,
            I => \N__47058\
        );

    \I__10328\ : InMux
    port map (
            O => \N__47061\,
            I => \N__47055\
        );

    \I__10327\ : Span4Mux_h
    port map (
            O => \N__47058\,
            I => \N__47052\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__47055\,
            I => \N__47049\
        );

    \I__10325\ : Odrv4
    port map (
            O => \N__47052\,
            I => duty_20
        );

    \I__10324\ : Odrv4
    port map (
            O => \N__47049\,
            I => duty_20
        );

    \I__10323\ : InMux
    port map (
            O => \N__47044\,
            I => \N__47041\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__47041\,
            I => n5_adj_571
        );

    \I__10321\ : CascadeMux
    port map (
            O => \N__47038\,
            I => \N__47035\
        );

    \I__10320\ : InMux
    port map (
            O => \N__47035\,
            I => \N__47032\
        );

    \I__10319\ : LocalMux
    port map (
            O => \N__47032\,
            I => \N__47026\
        );

    \I__10318\ : InMux
    port map (
            O => \N__47031\,
            I => \N__47021\
        );

    \I__10317\ : InMux
    port map (
            O => \N__47030\,
            I => \N__47021\
        );

    \I__10316\ : InMux
    port map (
            O => \N__47029\,
            I => \N__47018\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__47026\,
            I => \N__47015\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__47021\,
            I => \N__47012\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__47018\,
            I => pwm_counter_7
        );

    \I__10312\ : Odrv4
    port map (
            O => \N__47015\,
            I => pwm_counter_7
        );

    \I__10311\ : Odrv4
    port map (
            O => \N__47012\,
            I => pwm_counter_7
        );

    \I__10310\ : InMux
    port map (
            O => \N__47005\,
            I => \N__47002\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__47002\,
            I => \N__46999\
        );

    \I__10308\ : Span4Mux_h
    port map (
            O => \N__46999\,
            I => \N__46996\
        );

    \I__10307\ : Odrv4
    port map (
            O => \N__46996\,
            I => n10_adj_609
        );

    \I__10306\ : CascadeMux
    port map (
            O => \N__46993\,
            I => \n14722_cascade_\
        );

    \I__10305\ : CascadeMux
    port map (
            O => \N__46990\,
            I => \n14876_cascade_\
        );

    \I__10304\ : InMux
    port map (
            O => \N__46987\,
            I => \N__46984\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__46984\,
            I => n14886
        );

    \I__10302\ : InMux
    port map (
            O => \N__46981\,
            I => \N__46977\
        );

    \I__10301\ : InMux
    port map (
            O => \N__46980\,
            I => \N__46974\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__46977\,
            I => pwm_setpoint_15
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__46974\,
            I => pwm_setpoint_15
        );

    \I__10298\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46966\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__46966\,
            I => n14841
        );

    \I__10296\ : InMux
    port map (
            O => \N__46963\,
            I => \N__46960\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__46960\,
            I => n14781
        );

    \I__10294\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46954\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__46954\,
            I => \N__46951\
        );

    \I__10292\ : Odrv4
    port map (
            O => \N__46951\,
            I => \pwm_setpoint_23_N_171_7\
        );

    \I__10291\ : InMux
    port map (
            O => \N__46948\,
            I => \N__46944\
        );

    \I__10290\ : InMux
    port map (
            O => \N__46947\,
            I => \N__46941\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__46944\,
            I => \N__46938\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__46941\,
            I => \N__46935\
        );

    \I__10287\ : Span4Mux_h
    port map (
            O => \N__46938\,
            I => \N__46932\
        );

    \I__10286\ : Odrv12
    port map (
            O => \N__46935\,
            I => duty_7
        );

    \I__10285\ : Odrv4
    port map (
            O => \N__46932\,
            I => duty_7
        );

    \I__10284\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46923\
        );

    \I__10283\ : InMux
    port map (
            O => \N__46926\,
            I => \N__46919\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__46923\,
            I => \N__46916\
        );

    \I__10281\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46913\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__46919\,
            I => pwm_setpoint_7
        );

    \I__10279\ : Odrv4
    port map (
            O => \N__46916\,
            I => pwm_setpoint_7
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__46913\,
            I => pwm_setpoint_7
        );

    \I__10277\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46902\
        );

    \I__10276\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46899\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__46902\,
            I => pwm_setpoint_17
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__46899\,
            I => pwm_setpoint_17
        );

    \I__10273\ : CascadeMux
    port map (
            O => \N__46894\,
            I => \n12_adj_611_cascade_\
        );

    \I__10272\ : CascadeMux
    port map (
            O => \N__46891\,
            I => \N__46888\
        );

    \I__10271\ : InMux
    port map (
            O => \N__46888\,
            I => \N__46882\
        );

    \I__10270\ : InMux
    port map (
            O => \N__46887\,
            I => \N__46877\
        );

    \I__10269\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46877\
        );

    \I__10268\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46874\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__46882\,
            I => n35
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__46877\,
            I => n35
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__46874\,
            I => n35
        );

    \I__10264\ : InMux
    port map (
            O => \N__46867\,
            I => \N__46864\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__46864\,
            I => n30_adj_623
        );

    \I__10262\ : InMux
    port map (
            O => \N__46861\,
            I => \N__46854\
        );

    \I__10261\ : InMux
    port map (
            O => \N__46860\,
            I => \N__46854\
        );

    \I__10260\ : InMux
    port map (
            O => \N__46859\,
            I => \N__46851\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__46854\,
            I => \N__46848\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__46851\,
            I => pwm_setpoint_16
        );

    \I__10257\ : Odrv4
    port map (
            O => \N__46848\,
            I => pwm_setpoint_16
        );

    \I__10256\ : CascadeMux
    port map (
            O => \N__46843\,
            I => \N__46837\
        );

    \I__10255\ : InMux
    port map (
            O => \N__46842\,
            I => \N__46834\
        );

    \I__10254\ : InMux
    port map (
            O => \N__46841\,
            I => \N__46829\
        );

    \I__10253\ : InMux
    port map (
            O => \N__46840\,
            I => \N__46829\
        );

    \I__10252\ : InMux
    port map (
            O => \N__46837\,
            I => \N__46825\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__46834\,
            I => \N__46822\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__46829\,
            I => \N__46819\
        );

    \I__10249\ : InMux
    port map (
            O => \N__46828\,
            I => \N__46816\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__46825\,
            I => \N__46809\
        );

    \I__10247\ : Span4Mux_h
    port map (
            O => \N__46822\,
            I => \N__46809\
        );

    \I__10246\ : Span4Mux_s1_v
    port map (
            O => \N__46819\,
            I => \N__46809\
        );

    \I__10245\ : LocalMux
    port map (
            O => \N__46816\,
            I => pwm_counter_16
        );

    \I__10244\ : Odrv4
    port map (
            O => \N__46809\,
            I => pwm_counter_16
        );

    \I__10243\ : InMux
    port map (
            O => \N__46804\,
            I => \N__46801\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__46801\,
            I => \N__46798\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__46798\,
            I => n33_adj_625
        );

    \I__10240\ : InMux
    port map (
            O => \N__46795\,
            I => \N__46792\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__46792\,
            I => \N__46788\
        );

    \I__10238\ : InMux
    port map (
            O => \N__46791\,
            I => \N__46785\
        );

    \I__10237\ : Span4Mux_h
    port map (
            O => \N__46788\,
            I => \N__46782\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__46785\,
            I => \N__46779\
        );

    \I__10235\ : Odrv4
    port map (
            O => \N__46782\,
            I => duty_12
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__46779\,
            I => duty_12
        );

    \I__10233\ : InMux
    port map (
            O => \N__46774\,
            I => \N__46771\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__46771\,
            I => n13_adj_579
        );

    \I__10231\ : InMux
    port map (
            O => \N__46768\,
            I => \N__46763\
        );

    \I__10230\ : InMux
    port map (
            O => \N__46767\,
            I => \N__46760\
        );

    \I__10229\ : InMux
    port map (
            O => \N__46766\,
            I => \N__46757\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__46763\,
            I => \N__46754\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__46760\,
            I => pwm_counter_14
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__46757\,
            I => pwm_counter_14
        );

    \I__10225\ : Odrv12
    port map (
            O => \N__46754\,
            I => pwm_counter_14
        );

    \I__10224\ : InMux
    port map (
            O => \N__46747\,
            I => \N__46744\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__46744\,
            I => \N__46739\
        );

    \I__10222\ : InMux
    port map (
            O => \N__46743\,
            I => \N__46736\
        );

    \I__10221\ : InMux
    port map (
            O => \N__46742\,
            I => \N__46733\
        );

    \I__10220\ : Span4Mux_s2_v
    port map (
            O => \N__46739\,
            I => \N__46730\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__46736\,
            I => \N__46727\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__46733\,
            I => pwm_counter_13
        );

    \I__10217\ : Odrv4
    port map (
            O => \N__46730\,
            I => pwm_counter_13
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__46727\,
            I => pwm_counter_13
        );

    \I__10215\ : CascadeMux
    port map (
            O => \N__46720\,
            I => \N__46717\
        );

    \I__10214\ : InMux
    port map (
            O => \N__46717\,
            I => \N__46714\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__46714\,
            I => \N__46710\
        );

    \I__10212\ : InMux
    port map (
            O => \N__46713\,
            I => \N__46707\
        );

    \I__10211\ : Span4Mux_s2_v
    port map (
            O => \N__46710\,
            I => \N__46704\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__46707\,
            I => \N__46701\
        );

    \I__10209\ : Odrv4
    port map (
            O => \N__46704\,
            I => n27_adj_621
        );

    \I__10208\ : Odrv4
    port map (
            O => \N__46701\,
            I => n27_adj_621
        );

    \I__10207\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46690\
        );

    \I__10206\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46690\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__46690\,
            I => pwm_setpoint_13
        );

    \I__10204\ : CascadeMux
    port map (
            O => \N__46687\,
            I => \n27_adj_621_cascade_\
        );

    \I__10203\ : InMux
    port map (
            O => \N__46684\,
            I => \N__46681\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__46681\,
            I => n4_adj_605
        );

    \I__10201\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46672\
        );

    \I__10200\ : InMux
    port map (
            O => \N__46677\,
            I => \N__46672\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__46672\,
            I => pwm_setpoint_14
        );

    \I__10198\ : CascadeMux
    port map (
            O => \N__46669\,
            I => \n14840_cascade_\
        );

    \I__10197\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46662\
        );

    \I__10196\ : InMux
    port map (
            O => \N__46665\,
            I => \N__46659\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__46662\,
            I => \N__46654\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__46659\,
            I => \N__46654\
        );

    \I__10193\ : Odrv4
    port map (
            O => \N__46654\,
            I => duty_22
        );

    \I__10192\ : InMux
    port map (
            O => \N__46651\,
            I => \N__46648\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__46648\,
            I => n3_adj_569
        );

    \I__10190\ : InMux
    port map (
            O => \N__46645\,
            I => \N__46642\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__46642\,
            I => n9_adj_575
        );

    \I__10188\ : InMux
    port map (
            O => \N__46639\,
            I => \N__46633\
        );

    \I__10187\ : InMux
    port map (
            O => \N__46638\,
            I => \N__46633\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__46633\,
            I => \N__46630\
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__46630\,
            I => duty_16
        );

    \I__10184\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46624\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__46624\,
            I => \pwm_setpoint_23_N_171_16\
        );

    \I__10182\ : InMux
    port map (
            O => \N__46621\,
            I => \N__46618\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__46618\,
            I => \N__46615\
        );

    \I__10180\ : Span4Mux_h
    port map (
            O => \N__46615\,
            I => \N__46612\
        );

    \I__10179\ : Odrv4
    port map (
            O => \N__46612\,
            I => n3
        );

    \I__10178\ : InMux
    port map (
            O => \N__46609\,
            I => n12094
        );

    \I__10177\ : InMux
    port map (
            O => \N__46606\,
            I => \N__46603\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__46603\,
            I => \N__46600\
        );

    \I__10175\ : Odrv12
    port map (
            O => \N__46600\,
            I => n2
        );

    \I__10174\ : InMux
    port map (
            O => \N__46597\,
            I => n12095
        );

    \I__10173\ : InMux
    port map (
            O => \N__46594\,
            I => \N__46591\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__46591\,
            I => \pwm_setpoint_23_N_171_13\
        );

    \I__10171\ : InMux
    port map (
            O => \N__46588\,
            I => \N__46585\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__46585\,
            I => \N__46581\
        );

    \I__10169\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46578\
        );

    \I__10168\ : Span4Mux_s2_v
    port map (
            O => \N__46581\,
            I => \N__46573\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__46578\,
            I => \N__46573\
        );

    \I__10166\ : Odrv4
    port map (
            O => \N__46573\,
            I => duty_15
        );

    \I__10165\ : InMux
    port map (
            O => \N__46570\,
            I => \N__46567\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__46567\,
            I => n10_adj_576
        );

    \I__10163\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46561\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__46561\,
            I => \N__46557\
        );

    \I__10161\ : InMux
    port map (
            O => \N__46560\,
            I => \N__46554\
        );

    \I__10160\ : Odrv4
    port map (
            O => \N__46557\,
            I => duty_14
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__46554\,
            I => duty_14
        );

    \I__10158\ : InMux
    port map (
            O => \N__46549\,
            I => \N__46546\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__46546\,
            I => \pwm_setpoint_23_N_171_14\
        );

    \I__10156\ : InMux
    port map (
            O => \N__46543\,
            I => \N__46539\
        );

    \I__10155\ : InMux
    port map (
            O => \N__46542\,
            I => \N__46536\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__46539\,
            I => \N__46533\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__46536\,
            I => pwm_counter_1
        );

    \I__10152\ : Odrv4
    port map (
            O => \N__46533\,
            I => pwm_counter_1
        );

    \I__10151\ : CascadeMux
    port map (
            O => \N__46528\,
            I => \N__46525\
        );

    \I__10150\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46521\
        );

    \I__10149\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46518\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__46521\,
            I => \N__46515\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__46518\,
            I => pwm_counter_0
        );

    \I__10146\ : Odrv4
    port map (
            O => \N__46515\,
            I => pwm_counter_0
        );

    \I__10145\ : InMux
    port map (
            O => \N__46510\,
            I => \N__46507\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__46507\,
            I => n16_adj_582
        );

    \I__10143\ : InMux
    port map (
            O => \N__46504\,
            I => \N__46500\
        );

    \I__10142\ : InMux
    port map (
            O => \N__46503\,
            I => \N__46497\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__46500\,
            I => \N__46492\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__46497\,
            I => \N__46492\
        );

    \I__10139\ : Odrv4
    port map (
            O => \N__46492\,
            I => duty_13
        );

    \I__10138\ : InMux
    port map (
            O => \N__46489\,
            I => \N__46486\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__46486\,
            I => n12_adj_578
        );

    \I__10136\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46480\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__46480\,
            I => \pwm_setpoint_23_N_171_0\
        );

    \I__10134\ : InMux
    port map (
            O => \N__46477\,
            I => \N__46474\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__46474\,
            I => \N__46470\
        );

    \I__10132\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46467\
        );

    \I__10131\ : Odrv12
    port map (
            O => \N__46470\,
            I => duty_0
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__46467\,
            I => duty_0
        );

    \I__10129\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46459\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__46459\,
            I => pwm_setpoint_0
        );

    \I__10127\ : CascadeMux
    port map (
            O => \N__46456\,
            I => \N__46453\
        );

    \I__10126\ : InMux
    port map (
            O => \N__46453\,
            I => \N__46450\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46447\
        );

    \I__10124\ : Odrv12
    port map (
            O => \N__46447\,
            I => n11_adj_559
        );

    \I__10123\ : InMux
    port map (
            O => \N__46444\,
            I => n12086
        );

    \I__10122\ : InMux
    port map (
            O => \N__46441\,
            I => \N__46438\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__46438\,
            I => \N__46435\
        );

    \I__10120\ : Span4Mux_h
    port map (
            O => \N__46435\,
            I => \N__46432\
        );

    \I__10119\ : Odrv4
    port map (
            O => \N__46432\,
            I => n10_adj_560
        );

    \I__10118\ : InMux
    port map (
            O => \N__46429\,
            I => n12087
        );

    \I__10117\ : CascadeMux
    port map (
            O => \N__46426\,
            I => \N__46423\
        );

    \I__10116\ : InMux
    port map (
            O => \N__46423\,
            I => \N__46420\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__46420\,
            I => \N__46417\
        );

    \I__10114\ : Odrv4
    port map (
            O => \N__46417\,
            I => n9_adj_561
        );

    \I__10113\ : InMux
    port map (
            O => \N__46414\,
            I => \bfn_14_28_0_\
        );

    \I__10112\ : InMux
    port map (
            O => \N__46411\,
            I => \N__46408\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__46408\,
            I => \N__46405\
        );

    \I__10110\ : Odrv12
    port map (
            O => \N__46405\,
            I => n8_adj_562
        );

    \I__10109\ : InMux
    port map (
            O => \N__46402\,
            I => n12089
        );

    \I__10108\ : InMux
    port map (
            O => \N__46399\,
            I => \N__46396\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__46396\,
            I => \N__46393\
        );

    \I__10106\ : Odrv12
    port map (
            O => \N__46393\,
            I => n7_adj_563
        );

    \I__10105\ : InMux
    port map (
            O => \N__46390\,
            I => n12090
        );

    \I__10104\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46384\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__46384\,
            I => \N__46381\
        );

    \I__10102\ : Span4Mux_v
    port map (
            O => \N__46381\,
            I => \N__46378\
        );

    \I__10101\ : Odrv4
    port map (
            O => \N__46378\,
            I => n6_adj_564
        );

    \I__10100\ : InMux
    port map (
            O => \N__46375\,
            I => n12091
        );

    \I__10099\ : InMux
    port map (
            O => \N__46372\,
            I => \N__46369\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__46369\,
            I => \N__46366\
        );

    \I__10097\ : Odrv12
    port map (
            O => \N__46366\,
            I => n5_adj_565
        );

    \I__10096\ : InMux
    port map (
            O => \N__46363\,
            I => n12092
        );

    \I__10095\ : InMux
    port map (
            O => \N__46360\,
            I => \N__46357\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__46357\,
            I => \N__46354\
        );

    \I__10093\ : Span4Mux_v
    port map (
            O => \N__46354\,
            I => \N__46351\
        );

    \I__10092\ : Odrv4
    port map (
            O => \N__46351\,
            I => n4_adj_566
        );

    \I__10091\ : InMux
    port map (
            O => \N__46348\,
            I => \N__46344\
        );

    \I__10090\ : InMux
    port map (
            O => \N__46347\,
            I => \N__46341\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__46344\,
            I => \N__46338\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__46341\,
            I => \N__46335\
        );

    \I__10087\ : Span4Mux_h
    port map (
            O => \N__46338\,
            I => \N__46332\
        );

    \I__10086\ : Span4Mux_h
    port map (
            O => \N__46335\,
            I => \N__46329\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__46332\,
            I => duty_21
        );

    \I__10084\ : Odrv4
    port map (
            O => \N__46329\,
            I => duty_21
        );

    \I__10083\ : InMux
    port map (
            O => \N__46324\,
            I => n12093
        );

    \I__10082\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46318\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__46318\,
            I => \N__46315\
        );

    \I__10080\ : Span4Mux_h
    port map (
            O => \N__46315\,
            I => \N__46311\
        );

    \I__10079\ : InMux
    port map (
            O => \N__46314\,
            I => \N__46308\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__46311\,
            I => duty_6
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__46308\,
            I => duty_6
        );

    \I__10076\ : InMux
    port map (
            O => \N__46303\,
            I => n12078
        );

    \I__10075\ : CascadeMux
    port map (
            O => \N__46300\,
            I => \N__46297\
        );

    \I__10074\ : InMux
    port map (
            O => \N__46297\,
            I => \N__46294\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__46294\,
            I => \N__46291\
        );

    \I__10072\ : Odrv12
    port map (
            O => \N__46291\,
            I => n18_adj_552
        );

    \I__10071\ : InMux
    port map (
            O => \N__46288\,
            I => n12079
        );

    \I__10070\ : CascadeMux
    port map (
            O => \N__46285\,
            I => \N__46282\
        );

    \I__10069\ : InMux
    port map (
            O => \N__46282\,
            I => \N__46279\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__46279\,
            I => \N__46276\
        );

    \I__10067\ : Span4Mux_h
    port map (
            O => \N__46276\,
            I => \N__46273\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__46273\,
            I => n17_adj_553
        );

    \I__10065\ : InMux
    port map (
            O => \N__46270\,
            I => \bfn_14_27_0_\
        );

    \I__10064\ : CascadeMux
    port map (
            O => \N__46267\,
            I => \N__46264\
        );

    \I__10063\ : InMux
    port map (
            O => \N__46264\,
            I => \N__46261\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__46261\,
            I => \N__46258\
        );

    \I__10061\ : Span4Mux_h
    port map (
            O => \N__46258\,
            I => \N__46255\
        );

    \I__10060\ : Odrv4
    port map (
            O => \N__46255\,
            I => n16_adj_554
        );

    \I__10059\ : InMux
    port map (
            O => \N__46252\,
            I => n12081
        );

    \I__10058\ : CascadeMux
    port map (
            O => \N__46249\,
            I => \N__46246\
        );

    \I__10057\ : InMux
    port map (
            O => \N__46246\,
            I => \N__46243\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__46243\,
            I => \N__46240\
        );

    \I__10055\ : Span4Mux_h
    port map (
            O => \N__46240\,
            I => \N__46237\
        );

    \I__10054\ : Odrv4
    port map (
            O => \N__46237\,
            I => n15_adj_555
        );

    \I__10053\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46231\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__46231\,
            I => \N__46228\
        );

    \I__10051\ : Span4Mux_v
    port map (
            O => \N__46228\,
            I => \N__46224\
        );

    \I__10050\ : InMux
    port map (
            O => \N__46227\,
            I => \N__46221\
        );

    \I__10049\ : Odrv4
    port map (
            O => \N__46224\,
            I => duty_10
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__46221\,
            I => duty_10
        );

    \I__10047\ : InMux
    port map (
            O => \N__46216\,
            I => n12082
        );

    \I__10046\ : CascadeMux
    port map (
            O => \N__46213\,
            I => \N__46210\
        );

    \I__10045\ : InMux
    port map (
            O => \N__46210\,
            I => \N__46207\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__46207\,
            I => \N__46204\
        );

    \I__10043\ : Span4Mux_v
    port map (
            O => \N__46204\,
            I => \N__46201\
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__46201\,
            I => n14_adj_556
        );

    \I__10041\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46194\
        );

    \I__10040\ : InMux
    port map (
            O => \N__46197\,
            I => \N__46191\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__46194\,
            I => \N__46188\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__46191\,
            I => \N__46185\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__46188\,
            I => \N__46182\
        );

    \I__10036\ : Span4Mux_h
    port map (
            O => \N__46185\,
            I => \N__46179\
        );

    \I__10035\ : Odrv4
    port map (
            O => \N__46182\,
            I => duty_11
        );

    \I__10034\ : Odrv4
    port map (
            O => \N__46179\,
            I => duty_11
        );

    \I__10033\ : InMux
    port map (
            O => \N__46174\,
            I => n12083
        );

    \I__10032\ : InMux
    port map (
            O => \N__46171\,
            I => \N__46168\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__46168\,
            I => \N__46165\
        );

    \I__10030\ : Span4Mux_h
    port map (
            O => \N__46165\,
            I => \N__46162\
        );

    \I__10029\ : Odrv4
    port map (
            O => \N__46162\,
            I => n13_adj_557
        );

    \I__10028\ : InMux
    port map (
            O => \N__46159\,
            I => n12084
        );

    \I__10027\ : CascadeMux
    port map (
            O => \N__46156\,
            I => \N__46153\
        );

    \I__10026\ : InMux
    port map (
            O => \N__46153\,
            I => \N__46150\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__46150\,
            I => \N__46147\
        );

    \I__10024\ : Odrv12
    port map (
            O => \N__46147\,
            I => n12_adj_558
        );

    \I__10023\ : InMux
    port map (
            O => \N__46144\,
            I => n12085
        );

    \I__10022\ : CascadeMux
    port map (
            O => \N__46141\,
            I => \N__46138\
        );

    \I__10021\ : InMux
    port map (
            O => \N__46138\,
            I => \N__46135\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__46135\,
            I => \N__46130\
        );

    \I__10019\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46127\
        );

    \I__10018\ : InMux
    port map (
            O => \N__46133\,
            I => \N__46124\
        );

    \I__10017\ : Span4Mux_h
    port map (
            O => \N__46130\,
            I => \N__46121\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__46127\,
            I => n3223
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__46124\,
            I => n3223
        );

    \I__10014\ : Odrv4
    port map (
            O => \N__46121\,
            I => n3223
        );

    \I__10013\ : InMux
    port map (
            O => \N__46114\,
            I => \N__46111\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__46111\,
            I => n14366
        );

    \I__10011\ : InMux
    port map (
            O => \N__46108\,
            I => \N__46103\
        );

    \I__10010\ : InMux
    port map (
            O => \N__46107\,
            I => \N__46100\
        );

    \I__10009\ : InMux
    port map (
            O => \N__46106\,
            I => \N__46097\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__46103\,
            I => n3227
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__46100\,
            I => n3227
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__46097\,
            I => n3227
        );

    \I__10005\ : CascadeMux
    port map (
            O => \N__46090\,
            I => \N__46087\
        );

    \I__10004\ : InMux
    port map (
            O => \N__46087\,
            I => \N__46084\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__46084\,
            I => \N__46081\
        );

    \I__10002\ : Odrv12
    port map (
            O => \N__46081\,
            I => n25_adj_545
        );

    \I__10001\ : InMux
    port map (
            O => \N__46078\,
            I => \bfn_14_26_0_\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__46075\,
            I => \N__46072\
        );

    \I__9999\ : InMux
    port map (
            O => \N__46072\,
            I => \N__46069\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__46069\,
            I => \N__46066\
        );

    \I__9997\ : Odrv12
    port map (
            O => \N__46066\,
            I => n24_adj_546
        );

    \I__9996\ : InMux
    port map (
            O => \N__46063\,
            I => n12073
        );

    \I__9995\ : InMux
    port map (
            O => \N__46060\,
            I => \N__46057\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__46057\,
            I => \N__46054\
        );

    \I__9993\ : Span4Mux_h
    port map (
            O => \N__46054\,
            I => \N__46051\
        );

    \I__9992\ : Odrv4
    port map (
            O => \N__46051\,
            I => n23_adj_547
        );

    \I__9991\ : InMux
    port map (
            O => \N__46048\,
            I => \N__46045\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__46045\,
            I => \N__46042\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__46042\,
            I => \N__46038\
        );

    \I__9988\ : InMux
    port map (
            O => \N__46041\,
            I => \N__46035\
        );

    \I__9987\ : Odrv4
    port map (
            O => \N__46038\,
            I => duty_2
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__46035\,
            I => duty_2
        );

    \I__9985\ : InMux
    port map (
            O => \N__46030\,
            I => n12074
        );

    \I__9984\ : CascadeMux
    port map (
            O => \N__46027\,
            I => \N__46024\
        );

    \I__9983\ : InMux
    port map (
            O => \N__46024\,
            I => \N__46021\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__46021\,
            I => n22_adj_548
        );

    \I__9981\ : InMux
    port map (
            O => \N__46018\,
            I => n12075
        );

    \I__9980\ : CascadeMux
    port map (
            O => \N__46015\,
            I => \N__46012\
        );

    \I__9979\ : InMux
    port map (
            O => \N__46012\,
            I => \N__46009\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__46009\,
            I => \N__46006\
        );

    \I__9977\ : Odrv12
    port map (
            O => \N__46006\,
            I => n21_adj_549
        );

    \I__9976\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45999\
        );

    \I__9975\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45996\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__45999\,
            I => \N__45993\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__45996\,
            I => \N__45990\
        );

    \I__9972\ : Span4Mux_h
    port map (
            O => \N__45993\,
            I => \N__45987\
        );

    \I__9971\ : Span4Mux_h
    port map (
            O => \N__45990\,
            I => \N__45984\
        );

    \I__9970\ : Odrv4
    port map (
            O => \N__45987\,
            I => duty_4
        );

    \I__9969\ : Odrv4
    port map (
            O => \N__45984\,
            I => duty_4
        );

    \I__9968\ : InMux
    port map (
            O => \N__45979\,
            I => n12076
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__45976\,
            I => \N__45973\
        );

    \I__9966\ : InMux
    port map (
            O => \N__45973\,
            I => \N__45970\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__45970\,
            I => \N__45967\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__45967\,
            I => \N__45964\
        );

    \I__9963\ : Odrv4
    port map (
            O => \N__45964\,
            I => n20_adj_550
        );

    \I__9962\ : InMux
    port map (
            O => \N__45961\,
            I => \N__45958\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__45958\,
            I => \N__45955\
        );

    \I__9960\ : Span4Mux_h
    port map (
            O => \N__45955\,
            I => \N__45951\
        );

    \I__9959\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45948\
        );

    \I__9958\ : Odrv4
    port map (
            O => \N__45951\,
            I => duty_5
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__45948\,
            I => duty_5
        );

    \I__9956\ : InMux
    port map (
            O => \N__45943\,
            I => n12077
        );

    \I__9955\ : CascadeMux
    port map (
            O => \N__45940\,
            I => \N__45936\
        );

    \I__9954\ : InMux
    port map (
            O => \N__45939\,
            I => \N__45933\
        );

    \I__9953\ : InMux
    port map (
            O => \N__45936\,
            I => \N__45930\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__45933\,
            I => \N__45927\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__45930\,
            I => \N__45924\
        );

    \I__9950\ : Span4Mux_h
    port map (
            O => \N__45927\,
            I => \N__45919\
        );

    \I__9949\ : Span4Mux_v
    port map (
            O => \N__45924\,
            I => \N__45919\
        );

    \I__9948\ : Odrv4
    port map (
            O => \N__45919\,
            I => n3006
        );

    \I__9947\ : CascadeMux
    port map (
            O => \N__45916\,
            I => \N__45912\
        );

    \I__9946\ : InMux
    port map (
            O => \N__45915\,
            I => \N__45909\
        );

    \I__9945\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45906\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__45909\,
            I => \N__45903\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__45906\,
            I => \N__45900\
        );

    \I__9942\ : Span4Mux_h
    port map (
            O => \N__45903\,
            I => \N__45897\
        );

    \I__9941\ : Span4Mux_h
    port map (
            O => \N__45900\,
            I => \N__45894\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__45897\,
            I => n15123
        );

    \I__9939\ : Odrv4
    port map (
            O => \N__45894\,
            I => n15123
        );

    \I__9938\ : InMux
    port map (
            O => \N__45889\,
            I => n12491
        );

    \I__9937\ : InMux
    port map (
            O => \N__45886\,
            I => \N__45883\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__45883\,
            I => n3295
        );

    \I__9935\ : CascadeMux
    port map (
            O => \N__45880\,
            I => \N__45877\
        );

    \I__9934\ : InMux
    port map (
            O => \N__45877\,
            I => \N__45874\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__45874\,
            I => n3294
        );

    \I__9932\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45867\
        );

    \I__9931\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45864\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__45867\,
            I => \N__45860\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__45864\,
            I => \N__45857\
        );

    \I__9928\ : InMux
    port map (
            O => \N__45863\,
            I => \N__45854\
        );

    \I__9927\ : Span4Mux_v
    port map (
            O => \N__45860\,
            I => \N__45851\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__45857\,
            I => \N__45848\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__45854\,
            I => \N__45845\
        );

    \I__9924\ : Odrv4
    port map (
            O => \N__45851\,
            I => n3221
        );

    \I__9923\ : Odrv4
    port map (
            O => \N__45848\,
            I => n3221
        );

    \I__9922\ : Odrv12
    port map (
            O => \N__45845\,
            I => n3221
        );

    \I__9921\ : CascadeMux
    port map (
            O => \N__45838\,
            I => \N__45834\
        );

    \I__9920\ : InMux
    port map (
            O => \N__45837\,
            I => \N__45830\
        );

    \I__9919\ : InMux
    port map (
            O => \N__45834\,
            I => \N__45827\
        );

    \I__9918\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45824\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45821\
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__45827\,
            I => \N__45816\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__45824\,
            I => \N__45816\
        );

    \I__9914\ : Span4Mux_v
    port map (
            O => \N__45821\,
            I => \N__45813\
        );

    \I__9913\ : Span4Mux_v
    port map (
            O => \N__45816\,
            I => \N__45810\
        );

    \I__9912\ : Odrv4
    port map (
            O => \N__45813\,
            I => n3218
        );

    \I__9911\ : Odrv4
    port map (
            O => \N__45810\,
            I => n3218
        );

    \I__9910\ : CascadeMux
    port map (
            O => \N__45805\,
            I => \n14368_cascade_\
        );

    \I__9909\ : CascadeMux
    port map (
            O => \N__45802\,
            I => \N__45799\
        );

    \I__9908\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45796\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__45796\,
            I => \N__45793\
        );

    \I__9906\ : Span4Mux_v
    port map (
            O => \N__45793\,
            I => \N__45790\
        );

    \I__9905\ : Odrv4
    port map (
            O => \N__45790\,
            I => n14374
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__45787\,
            I => \N__45784\
        );

    \I__9903\ : InMux
    port map (
            O => \N__45784\,
            I => \N__45780\
        );

    \I__9902\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45777\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__45780\,
            I => \N__45774\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__45777\,
            I => n3228
        );

    \I__9899\ : Odrv4
    port map (
            O => \N__45774\,
            I => n3228
        );

    \I__9898\ : CascadeMux
    port map (
            O => \N__45769\,
            I => \n3228_cascade_\
        );

    \I__9897\ : InMux
    port map (
            O => \N__45766\,
            I => \N__45762\
        );

    \I__9896\ : InMux
    port map (
            O => \N__45765\,
            I => \N__45759\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__45762\,
            I => \N__45753\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__45759\,
            I => \N__45753\
        );

    \I__9893\ : InMux
    port map (
            O => \N__45758\,
            I => \N__45750\
        );

    \I__9892\ : Odrv4
    port map (
            O => \N__45753\,
            I => n3224
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__45750\,
            I => n3224
        );

    \I__9890\ : CascadeMux
    port map (
            O => \N__45745\,
            I => \N__45742\
        );

    \I__9889\ : InMux
    port map (
            O => \N__45742\,
            I => \N__45739\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__45739\,
            I => n14362
        );

    \I__9887\ : CascadeMux
    port map (
            O => \N__45736\,
            I => \N__45733\
        );

    \I__9886\ : InMux
    port map (
            O => \N__45733\,
            I => \N__45729\
        );

    \I__9885\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45726\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__45729\,
            I => n3014
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__45726\,
            I => n3014
        );

    \I__9882\ : InMux
    port map (
            O => \N__45721\,
            I => \N__45718\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__45718\,
            I => \N__45715\
        );

    \I__9880\ : Odrv4
    port map (
            O => \N__45715\,
            I => n3081
        );

    \I__9879\ : InMux
    port map (
            O => \N__45712\,
            I => n12483
        );

    \I__9878\ : InMux
    port map (
            O => \N__45709\,
            I => \N__45706\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__45706\,
            I => \N__45701\
        );

    \I__9876\ : InMux
    port map (
            O => \N__45705\,
            I => \N__45698\
        );

    \I__9875\ : InMux
    port map (
            O => \N__45704\,
            I => \N__45695\
        );

    \I__9874\ : Span4Mux_h
    port map (
            O => \N__45701\,
            I => \N__45692\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__45698\,
            I => \N__45689\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__45695\,
            I => n3013
        );

    \I__9871\ : Odrv4
    port map (
            O => \N__45692\,
            I => n3013
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__45689\,
            I => n3013
        );

    \I__9869\ : InMux
    port map (
            O => \N__45682\,
            I => \N__45679\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__45679\,
            I => \N__45676\
        );

    \I__9867\ : Odrv4
    port map (
            O => \N__45676\,
            I => n3080
        );

    \I__9866\ : InMux
    port map (
            O => \N__45673\,
            I => n12484
        );

    \I__9865\ : InMux
    port map (
            O => \N__45670\,
            I => \N__45665\
        );

    \I__9864\ : InMux
    port map (
            O => \N__45669\,
            I => \N__45662\
        );

    \I__9863\ : CascadeMux
    port map (
            O => \N__45668\,
            I => \N__45659\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__45665\,
            I => \N__45654\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__45662\,
            I => \N__45654\
        );

    \I__9860\ : InMux
    port map (
            O => \N__45659\,
            I => \N__45651\
        );

    \I__9859\ : Odrv4
    port map (
            O => \N__45654\,
            I => n3012
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__45651\,
            I => n3012
        );

    \I__9857\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45643\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__45643\,
            I => \N__45640\
        );

    \I__9855\ : Odrv12
    port map (
            O => \N__45640\,
            I => n3079
        );

    \I__9854\ : InMux
    port map (
            O => \N__45637\,
            I => n12485
        );

    \I__9853\ : InMux
    port map (
            O => \N__45634\,
            I => n12486
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__45631\,
            I => \N__45628\
        );

    \I__9851\ : InMux
    port map (
            O => \N__45628\,
            I => \N__45625\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__45625\,
            I => \N__45622\
        );

    \I__9849\ : Span4Mux_v
    port map (
            O => \N__45622\,
            I => \N__45618\
        );

    \I__9848\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45615\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__45618\,
            I => n3010
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__45615\,
            I => n3010
        );

    \I__9845\ : InMux
    port map (
            O => \N__45610\,
            I => \N__45607\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__45607\,
            I => \N__45604\
        );

    \I__9843\ : Span4Mux_v
    port map (
            O => \N__45604\,
            I => \N__45601\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__45601\,
            I => \N__45598\
        );

    \I__9841\ : Odrv4
    port map (
            O => \N__45598\,
            I => n3077
        );

    \I__9840\ : InMux
    port map (
            O => \N__45595\,
            I => \bfn_14_24_0_\
        );

    \I__9839\ : InMux
    port map (
            O => \N__45592\,
            I => n12488
        );

    \I__9838\ : InMux
    port map (
            O => \N__45589\,
            I => \N__45585\
        );

    \I__9837\ : InMux
    port map (
            O => \N__45588\,
            I => \N__45582\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__45585\,
            I => \N__45579\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__45582\,
            I => \N__45575\
        );

    \I__9834\ : Span4Mux_v
    port map (
            O => \N__45579\,
            I => \N__45572\
        );

    \I__9833\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45569\
        );

    \I__9832\ : Odrv4
    port map (
            O => \N__45575\,
            I => n3008
        );

    \I__9831\ : Odrv4
    port map (
            O => \N__45572\,
            I => n3008
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__45569\,
            I => n3008
        );

    \I__9829\ : CascadeMux
    port map (
            O => \N__45562\,
            I => \N__45559\
        );

    \I__9828\ : InMux
    port map (
            O => \N__45559\,
            I => \N__45556\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__45556\,
            I => \N__45553\
        );

    \I__9826\ : Span4Mux_h
    port map (
            O => \N__45553\,
            I => \N__45550\
        );

    \I__9825\ : Odrv4
    port map (
            O => \N__45550\,
            I => n3075
        );

    \I__9824\ : InMux
    port map (
            O => \N__45547\,
            I => n12489
        );

    \I__9823\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45540\
        );

    \I__9822\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45537\
        );

    \I__9821\ : LocalMux
    port map (
            O => \N__45540\,
            I => \N__45534\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__45537\,
            I => \N__45530\
        );

    \I__9819\ : Span4Mux_h
    port map (
            O => \N__45534\,
            I => \N__45527\
        );

    \I__9818\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45524\
        );

    \I__9817\ : Odrv4
    port map (
            O => \N__45530\,
            I => n3007
        );

    \I__9816\ : Odrv4
    port map (
            O => \N__45527\,
            I => n3007
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__45524\,
            I => n3007
        );

    \I__9814\ : CascadeMux
    port map (
            O => \N__45517\,
            I => \N__45514\
        );

    \I__9813\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45511\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__45511\,
            I => \N__45508\
        );

    \I__9811\ : Span4Mux_v
    port map (
            O => \N__45508\,
            I => \N__45505\
        );

    \I__9810\ : Span4Mux_h
    port map (
            O => \N__45505\,
            I => \N__45502\
        );

    \I__9809\ : Odrv4
    port map (
            O => \N__45502\,
            I => n3074
        );

    \I__9808\ : InMux
    port map (
            O => \N__45499\,
            I => n12490
        );

    \I__9807\ : CascadeMux
    port map (
            O => \N__45496\,
            I => \N__45492\
        );

    \I__9806\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45488\
        );

    \I__9805\ : InMux
    port map (
            O => \N__45492\,
            I => \N__45485\
        );

    \I__9804\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45482\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__45488\,
            I => n3022
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__45485\,
            I => n3022
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__45482\,
            I => n3022
        );

    \I__9800\ : CascadeMux
    port map (
            O => \N__45475\,
            I => \N__45472\
        );

    \I__9799\ : InMux
    port map (
            O => \N__45472\,
            I => \N__45469\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__45469\,
            I => \N__45466\
        );

    \I__9797\ : Span4Mux_v
    port map (
            O => \N__45466\,
            I => \N__45463\
        );

    \I__9796\ : Odrv4
    port map (
            O => \N__45463\,
            I => n3089
        );

    \I__9795\ : InMux
    port map (
            O => \N__45460\,
            I => n12475
        );

    \I__9794\ : CascadeMux
    port map (
            O => \N__45457\,
            I => \N__45453\
        );

    \I__9793\ : CascadeMux
    port map (
            O => \N__45456\,
            I => \N__45450\
        );

    \I__9792\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45447\
        );

    \I__9791\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45444\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__45447\,
            I => n3021
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__45444\,
            I => n3021
        );

    \I__9788\ : InMux
    port map (
            O => \N__45439\,
            I => \N__45436\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__45436\,
            I => n3088
        );

    \I__9786\ : InMux
    port map (
            O => \N__45433\,
            I => n12476
        );

    \I__9785\ : CascadeMux
    port map (
            O => \N__45430\,
            I => \N__45427\
        );

    \I__9784\ : InMux
    port map (
            O => \N__45427\,
            I => \N__45424\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__45424\,
            I => \N__45419\
        );

    \I__9782\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45416\
        );

    \I__9781\ : InMux
    port map (
            O => \N__45422\,
            I => \N__45413\
        );

    \I__9780\ : Span4Mux_v
    port map (
            O => \N__45419\,
            I => \N__45408\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__45416\,
            I => \N__45408\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__45413\,
            I => n3020
        );

    \I__9777\ : Odrv4
    port map (
            O => \N__45408\,
            I => n3020
        );

    \I__9776\ : CascadeMux
    port map (
            O => \N__45403\,
            I => \N__45400\
        );

    \I__9775\ : InMux
    port map (
            O => \N__45400\,
            I => \N__45397\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__45397\,
            I => \N__45394\
        );

    \I__9773\ : Span4Mux_v
    port map (
            O => \N__45394\,
            I => \N__45391\
        );

    \I__9772\ : Span4Mux_h
    port map (
            O => \N__45391\,
            I => \N__45388\
        );

    \I__9771\ : Odrv4
    port map (
            O => \N__45388\,
            I => n3087
        );

    \I__9770\ : InMux
    port map (
            O => \N__45385\,
            I => n12477
        );

    \I__9769\ : InMux
    port map (
            O => \N__45382\,
            I => \N__45379\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__45379\,
            I => \N__45375\
        );

    \I__9767\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45372\
        );

    \I__9766\ : Span4Mux_v
    port map (
            O => \N__45375\,
            I => \N__45367\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__45372\,
            I => \N__45367\
        );

    \I__9764\ : Odrv4
    port map (
            O => \N__45367\,
            I => n3019
        );

    \I__9763\ : InMux
    port map (
            O => \N__45364\,
            I => \N__45361\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__45361\,
            I => \N__45358\
        );

    \I__9761\ : Span4Mux_v
    port map (
            O => \N__45358\,
            I => \N__45355\
        );

    \I__9760\ : Odrv4
    port map (
            O => \N__45355\,
            I => n3086
        );

    \I__9759\ : InMux
    port map (
            O => \N__45352\,
            I => n12478
        );

    \I__9758\ : CascadeMux
    port map (
            O => \N__45349\,
            I => \N__45346\
        );

    \I__9757\ : InMux
    port map (
            O => \N__45346\,
            I => \N__45342\
        );

    \I__9756\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45339\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__45342\,
            I => \N__45333\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__45339\,
            I => \N__45333\
        );

    \I__9753\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45330\
        );

    \I__9752\ : Span4Mux_v
    port map (
            O => \N__45333\,
            I => \N__45327\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__45330\,
            I => n3018
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__45327\,
            I => n3018
        );

    \I__9749\ : InMux
    port map (
            O => \N__45322\,
            I => \N__45319\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__45319\,
            I => \N__45316\
        );

    \I__9747\ : Span4Mux_h
    port map (
            O => \N__45316\,
            I => \N__45313\
        );

    \I__9746\ : Odrv4
    port map (
            O => \N__45313\,
            I => n3085
        );

    \I__9745\ : InMux
    port map (
            O => \N__45310\,
            I => \bfn_14_23_0_\
        );

    \I__9744\ : InMux
    port map (
            O => \N__45307\,
            I => \N__45304\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__45304\,
            I => \N__45300\
        );

    \I__9742\ : InMux
    port map (
            O => \N__45303\,
            I => \N__45297\
        );

    \I__9741\ : Span4Mux_h
    port map (
            O => \N__45300\,
            I => \N__45292\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__45297\,
            I => \N__45292\
        );

    \I__9739\ : Odrv4
    port map (
            O => \N__45292\,
            I => n3017
        );

    \I__9738\ : InMux
    port map (
            O => \N__45289\,
            I => \N__45286\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__45286\,
            I => \N__45283\
        );

    \I__9736\ : Span4Mux_h
    port map (
            O => \N__45283\,
            I => \N__45280\
        );

    \I__9735\ : Odrv4
    port map (
            O => \N__45280\,
            I => n3084
        );

    \I__9734\ : InMux
    port map (
            O => \N__45277\,
            I => n12480
        );

    \I__9733\ : InMux
    port map (
            O => \N__45274\,
            I => \N__45270\
        );

    \I__9732\ : CascadeMux
    port map (
            O => \N__45273\,
            I => \N__45266\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__45270\,
            I => \N__45263\
        );

    \I__9730\ : InMux
    port map (
            O => \N__45269\,
            I => \N__45260\
        );

    \I__9729\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45257\
        );

    \I__9728\ : Span4Mux_v
    port map (
            O => \N__45263\,
            I => \N__45252\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__45260\,
            I => \N__45252\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__45257\,
            I => n3016
        );

    \I__9725\ : Odrv4
    port map (
            O => \N__45252\,
            I => n3016
        );

    \I__9724\ : InMux
    port map (
            O => \N__45247\,
            I => \N__45244\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__45244\,
            I => \N__45241\
        );

    \I__9722\ : Span4Mux_v
    port map (
            O => \N__45241\,
            I => \N__45238\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__45238\,
            I => n3083
        );

    \I__9720\ : InMux
    port map (
            O => \N__45235\,
            I => n12481
        );

    \I__9719\ : InMux
    port map (
            O => \N__45232\,
            I => n12482
        );

    \I__9718\ : CascadeMux
    port map (
            O => \N__45229\,
            I => \N__45226\
        );

    \I__9717\ : InMux
    port map (
            O => \N__45226\,
            I => \N__45222\
        );

    \I__9716\ : InMux
    port map (
            O => \N__45225\,
            I => \N__45218\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__45222\,
            I => \N__45215\
        );

    \I__9714\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45212\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__45218\,
            I => n3030
        );

    \I__9712\ : Odrv4
    port map (
            O => \N__45215\,
            I => n3030
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__45212\,
            I => n3030
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__45205\,
            I => \N__45202\
        );

    \I__9709\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45199\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__45199\,
            I => \N__45196\
        );

    \I__9707\ : Span4Mux_v
    port map (
            O => \N__45196\,
            I => \N__45193\
        );

    \I__9706\ : Odrv4
    port map (
            O => \N__45193\,
            I => n3097
        );

    \I__9705\ : InMux
    port map (
            O => \N__45190\,
            I => n12467
        );

    \I__9704\ : InMux
    port map (
            O => \N__45187\,
            I => \N__45184\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__45184\,
            I => \N__45181\
        );

    \I__9702\ : Span4Mux_v
    port map (
            O => \N__45181\,
            I => \N__45177\
        );

    \I__9701\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45174\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__45177\,
            I => n3029
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__45174\,
            I => n3029
        );

    \I__9698\ : InMux
    port map (
            O => \N__45169\,
            I => \N__45166\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__45166\,
            I => \N__45163\
        );

    \I__9696\ : Span4Mux_h
    port map (
            O => \N__45163\,
            I => \N__45160\
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__45160\,
            I => n3096
        );

    \I__9694\ : InMux
    port map (
            O => \N__45157\,
            I => n12468
        );

    \I__9693\ : CascadeMux
    port map (
            O => \N__45154\,
            I => \N__45151\
        );

    \I__9692\ : InMux
    port map (
            O => \N__45151\,
            I => \N__45147\
        );

    \I__9691\ : InMux
    port map (
            O => \N__45150\,
            I => \N__45143\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__45147\,
            I => \N__45140\
        );

    \I__9689\ : InMux
    port map (
            O => \N__45146\,
            I => \N__45137\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__45143\,
            I => n3028
        );

    \I__9687\ : Odrv4
    port map (
            O => \N__45140\,
            I => n3028
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__45137\,
            I => n3028
        );

    \I__9685\ : InMux
    port map (
            O => \N__45130\,
            I => \N__45127\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__45127\,
            I => \N__45124\
        );

    \I__9683\ : Odrv12
    port map (
            O => \N__45124\,
            I => n3095
        );

    \I__9682\ : InMux
    port map (
            O => \N__45121\,
            I => n12469
        );

    \I__9681\ : CascadeMux
    port map (
            O => \N__45118\,
            I => \N__45114\
        );

    \I__9680\ : InMux
    port map (
            O => \N__45117\,
            I => \N__45110\
        );

    \I__9679\ : InMux
    port map (
            O => \N__45114\,
            I => \N__45107\
        );

    \I__9678\ : InMux
    port map (
            O => \N__45113\,
            I => \N__45104\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__45110\,
            I => n3027
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__45107\,
            I => n3027
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__45104\,
            I => n3027
        );

    \I__9674\ : InMux
    port map (
            O => \N__45097\,
            I => \N__45094\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__45094\,
            I => n3094
        );

    \I__9672\ : InMux
    port map (
            O => \N__45091\,
            I => n12470
        );

    \I__9671\ : CascadeMux
    port map (
            O => \N__45088\,
            I => \N__45084\
        );

    \I__9670\ : InMux
    port map (
            O => \N__45087\,
            I => \N__45080\
        );

    \I__9669\ : InMux
    port map (
            O => \N__45084\,
            I => \N__45077\
        );

    \I__9668\ : InMux
    port map (
            O => \N__45083\,
            I => \N__45074\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__45080\,
            I => n3026
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__45077\,
            I => n3026
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__45074\,
            I => n3026
        );

    \I__9664\ : InMux
    port map (
            O => \N__45067\,
            I => \N__45064\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__45064\,
            I => n3093
        );

    \I__9662\ : InMux
    port map (
            O => \N__45061\,
            I => \bfn_14_22_0_\
        );

    \I__9661\ : CascadeMux
    port map (
            O => \N__45058\,
            I => \N__45055\
        );

    \I__9660\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45051\
        );

    \I__9659\ : CascadeMux
    port map (
            O => \N__45054\,
            I => \N__45048\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__45051\,
            I => \N__45045\
        );

    \I__9657\ : InMux
    port map (
            O => \N__45048\,
            I => \N__45041\
        );

    \I__9656\ : Span4Mux_h
    port map (
            O => \N__45045\,
            I => \N__45038\
        );

    \I__9655\ : InMux
    port map (
            O => \N__45044\,
            I => \N__45035\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__45041\,
            I => n3025
        );

    \I__9653\ : Odrv4
    port map (
            O => \N__45038\,
            I => n3025
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__45035\,
            I => n3025
        );

    \I__9651\ : InMux
    port map (
            O => \N__45028\,
            I => \N__45025\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__45025\,
            I => \N__45022\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__45022\,
            I => \N__45019\
        );

    \I__9648\ : Odrv4
    port map (
            O => \N__45019\,
            I => n3092
        );

    \I__9647\ : InMux
    port map (
            O => \N__45016\,
            I => n12472
        );

    \I__9646\ : CascadeMux
    port map (
            O => \N__45013\,
            I => \N__45009\
        );

    \I__9645\ : InMux
    port map (
            O => \N__45012\,
            I => \N__45005\
        );

    \I__9644\ : InMux
    port map (
            O => \N__45009\,
            I => \N__45002\
        );

    \I__9643\ : InMux
    port map (
            O => \N__45008\,
            I => \N__44999\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__45005\,
            I => n3024
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__45002\,
            I => n3024
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__44999\,
            I => n3024
        );

    \I__9639\ : InMux
    port map (
            O => \N__44992\,
            I => \N__44989\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__44989\,
            I => \N__44986\
        );

    \I__9637\ : Odrv4
    port map (
            O => \N__44986\,
            I => n3091
        );

    \I__9636\ : InMux
    port map (
            O => \N__44983\,
            I => n12473
        );

    \I__9635\ : CascadeMux
    port map (
            O => \N__44980\,
            I => \N__44976\
        );

    \I__9634\ : InMux
    port map (
            O => \N__44979\,
            I => \N__44973\
        );

    \I__9633\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44970\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__44973\,
            I => n3023
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__44970\,
            I => n3023
        );

    \I__9630\ : CascadeMux
    port map (
            O => \N__44965\,
            I => \N__44962\
        );

    \I__9629\ : InMux
    port map (
            O => \N__44962\,
            I => \N__44959\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__44959\,
            I => \N__44956\
        );

    \I__9627\ : Odrv4
    port map (
            O => \N__44956\,
            I => n3090
        );

    \I__9626\ : InMux
    port map (
            O => \N__44953\,
            I => n12474
        );

    \I__9625\ : CascadeMux
    port map (
            O => \N__44950\,
            I => \N__44947\
        );

    \I__9624\ : InMux
    port map (
            O => \N__44947\,
            I => \N__44944\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__44944\,
            I => \N__44940\
        );

    \I__9622\ : InMux
    port map (
            O => \N__44943\,
            I => \N__44936\
        );

    \I__9621\ : Span4Mux_v
    port map (
            O => \N__44940\,
            I => \N__44933\
        );

    \I__9620\ : InMux
    port map (
            O => \N__44939\,
            I => \N__44930\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__44936\,
            I => n2925
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__44933\,
            I => n2925
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__44930\,
            I => n2925
        );

    \I__9616\ : CascadeMux
    port map (
            O => \N__44923\,
            I => \n3122_cascade_\
        );

    \I__9615\ : InMux
    port map (
            O => \N__44920\,
            I => \N__44916\
        );

    \I__9614\ : InMux
    port map (
            O => \N__44919\,
            I => \N__44913\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__44916\,
            I => \N__44907\
        );

    \I__9612\ : LocalMux
    port map (
            O => \N__44913\,
            I => \N__44907\
        );

    \I__9611\ : InMux
    port map (
            O => \N__44912\,
            I => \N__44904\
        );

    \I__9610\ : Span4Mux_v
    port map (
            O => \N__44907\,
            I => \N__44899\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__44904\,
            I => \N__44899\
        );

    \I__9608\ : Span4Mux_h
    port map (
            O => \N__44899\,
            I => \N__44896\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__44896\,
            I => n2914
        );

    \I__9606\ : InMux
    port map (
            O => \N__44893\,
            I => \N__44889\
        );

    \I__9605\ : InMux
    port map (
            O => \N__44892\,
            I => \N__44885\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__44889\,
            I => \N__44882\
        );

    \I__9603\ : InMux
    port map (
            O => \N__44888\,
            I => \N__44879\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__44885\,
            I => \N__44876\
        );

    \I__9601\ : Span4Mux_h
    port map (
            O => \N__44882\,
            I => \N__44873\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__44879\,
            I => \N__44870\
        );

    \I__9599\ : Span4Mux_h
    port map (
            O => \N__44876\,
            I => \N__44867\
        );

    \I__9598\ : Span4Mux_h
    port map (
            O => \N__44873\,
            I => \N__44864\
        );

    \I__9597\ : Span4Mux_h
    port map (
            O => \N__44870\,
            I => \N__44861\
        );

    \I__9596\ : Odrv4
    port map (
            O => \N__44867\,
            I => n316
        );

    \I__9595\ : Odrv4
    port map (
            O => \N__44864\,
            I => n316
        );

    \I__9594\ : Odrv4
    port map (
            O => \N__44861\,
            I => n316
        );

    \I__9593\ : InMux
    port map (
            O => \N__44854\,
            I => \N__44851\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__44851\,
            I => \N__44848\
        );

    \I__9591\ : Span4Mux_h
    port map (
            O => \N__44848\,
            I => \N__44845\
        );

    \I__9590\ : Span4Mux_h
    port map (
            O => \N__44845\,
            I => \N__44842\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__44842\,
            I => n3101
        );

    \I__9588\ : InMux
    port map (
            O => \N__44839\,
            I => \bfn_14_21_0_\
        );

    \I__9587\ : CascadeMux
    port map (
            O => \N__44836\,
            I => \N__44832\
        );

    \I__9586\ : InMux
    port map (
            O => \N__44835\,
            I => \N__44829\
        );

    \I__9585\ : InMux
    port map (
            O => \N__44832\,
            I => \N__44826\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__44829\,
            I => \N__44823\
        );

    \I__9583\ : LocalMux
    port map (
            O => \N__44826\,
            I => \N__44820\
        );

    \I__9582\ : Span4Mux_h
    port map (
            O => \N__44823\,
            I => \N__44816\
        );

    \I__9581\ : Span4Mux_h
    port map (
            O => \N__44820\,
            I => \N__44813\
        );

    \I__9580\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44810\
        );

    \I__9579\ : Odrv4
    port map (
            O => \N__44816\,
            I => n3033
        );

    \I__9578\ : Odrv4
    port map (
            O => \N__44813\,
            I => n3033
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__44810\,
            I => n3033
        );

    \I__9576\ : InMux
    port map (
            O => \N__44803\,
            I => \N__44800\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__44800\,
            I => \N__44797\
        );

    \I__9574\ : Span12Mux_s11_v
    port map (
            O => \N__44797\,
            I => \N__44794\
        );

    \I__9573\ : Odrv12
    port map (
            O => \N__44794\,
            I => n3100
        );

    \I__9572\ : InMux
    port map (
            O => \N__44791\,
            I => n12464
        );

    \I__9571\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44784\
        );

    \I__9570\ : InMux
    port map (
            O => \N__44787\,
            I => \N__44781\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__44784\,
            I => \N__44778\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__44781\,
            I => \N__44775\
        );

    \I__9567\ : Span4Mux_h
    port map (
            O => \N__44778\,
            I => \N__44772\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__44775\,
            I => \N__44769\
        );

    \I__9565\ : Odrv4
    port map (
            O => \N__44772\,
            I => n3032
        );

    \I__9564\ : Odrv4
    port map (
            O => \N__44769\,
            I => n3032
        );

    \I__9563\ : CascadeMux
    port map (
            O => \N__44764\,
            I => \N__44761\
        );

    \I__9562\ : InMux
    port map (
            O => \N__44761\,
            I => \N__44758\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__44758\,
            I => \N__44755\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__44755\,
            I => \N__44752\
        );

    \I__9559\ : Span4Mux_h
    port map (
            O => \N__44752\,
            I => \N__44749\
        );

    \I__9558\ : Odrv4
    port map (
            O => \N__44749\,
            I => n3099
        );

    \I__9557\ : InMux
    port map (
            O => \N__44746\,
            I => n12465
        );

    \I__9556\ : CascadeMux
    port map (
            O => \N__44743\,
            I => \N__44739\
        );

    \I__9555\ : InMux
    port map (
            O => \N__44742\,
            I => \N__44736\
        );

    \I__9554\ : InMux
    port map (
            O => \N__44739\,
            I => \N__44733\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__44736\,
            I => \N__44729\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__44733\,
            I => \N__44726\
        );

    \I__9551\ : InMux
    port map (
            O => \N__44732\,
            I => \N__44723\
        );

    \I__9550\ : Odrv4
    port map (
            O => \N__44729\,
            I => n3031
        );

    \I__9549\ : Odrv4
    port map (
            O => \N__44726\,
            I => n3031
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__44723\,
            I => n3031
        );

    \I__9547\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44713\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__44713\,
            I => n3098
        );

    \I__9545\ : InMux
    port map (
            O => \N__44710\,
            I => n12466
        );

    \I__9544\ : CascadeMux
    port map (
            O => \N__44707\,
            I => \n13932_cascade_\
        );

    \I__9543\ : InMux
    port map (
            O => \N__44704\,
            I => \N__44701\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__44701\,
            I => n13936
        );

    \I__9541\ : InMux
    port map (
            O => \N__44698\,
            I => \N__44694\
        );

    \I__9540\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44691\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__44694\,
            I => \N__44688\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__44691\,
            I => \N__44685\
        );

    \I__9537\ : Span4Mux_v
    port map (
            O => \N__44688\,
            I => \N__44681\
        );

    \I__9536\ : Span4Mux_h
    port map (
            O => \N__44685\,
            I => \N__44678\
        );

    \I__9535\ : InMux
    port map (
            O => \N__44684\,
            I => \N__44675\
        );

    \I__9534\ : Odrv4
    port map (
            O => \N__44681\,
            I => n2926
        );

    \I__9533\ : Odrv4
    port map (
            O => \N__44678\,
            I => n2926
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__44675\,
            I => n2926
        );

    \I__9531\ : CascadeMux
    port map (
            O => \N__44668\,
            I => \N__44664\
        );

    \I__9530\ : CascadeMux
    port map (
            O => \N__44667\,
            I => \N__44661\
        );

    \I__9529\ : InMux
    port map (
            O => \N__44664\,
            I => \N__44658\
        );

    \I__9528\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44655\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__44658\,
            I => \N__44651\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__44655\,
            I => \N__44648\
        );

    \I__9525\ : CascadeMux
    port map (
            O => \N__44654\,
            I => \N__44645\
        );

    \I__9524\ : Span4Mux_v
    port map (
            O => \N__44651\,
            I => \N__44642\
        );

    \I__9523\ : Span4Mux_h
    port map (
            O => \N__44648\,
            I => \N__44639\
        );

    \I__9522\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44636\
        );

    \I__9521\ : Odrv4
    port map (
            O => \N__44642\,
            I => n2920
        );

    \I__9520\ : Odrv4
    port map (
            O => \N__44639\,
            I => n2920
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__44636\,
            I => n2920
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__44629\,
            I => \N__44626\
        );

    \I__9517\ : InMux
    port map (
            O => \N__44626\,
            I => \N__44622\
        );

    \I__9516\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44619\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__44622\,
            I => \N__44616\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__44619\,
            I => \N__44610\
        );

    \I__9513\ : Span4Mux_h
    port map (
            O => \N__44616\,
            I => \N__44610\
        );

    \I__9512\ : InMux
    port map (
            O => \N__44615\,
            I => \N__44607\
        );

    \I__9511\ : Odrv4
    port map (
            O => \N__44610\,
            I => n2927
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__44607\,
            I => n2927
        );

    \I__9509\ : InMux
    port map (
            O => \N__44602\,
            I => \N__44598\
        );

    \I__9508\ : InMux
    port map (
            O => \N__44601\,
            I => \N__44595\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__44598\,
            I => \N__44592\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__44595\,
            I => \N__44589\
        );

    \I__9505\ : Span4Mux_v
    port map (
            O => \N__44592\,
            I => \N__44585\
        );

    \I__9504\ : Span4Mux_h
    port map (
            O => \N__44589\,
            I => \N__44582\
        );

    \I__9503\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44579\
        );

    \I__9502\ : Odrv4
    port map (
            O => \N__44585\,
            I => n2919
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__44582\,
            I => n2919
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__44579\,
            I => n2919
        );

    \I__9499\ : CascadeMux
    port map (
            O => \N__44572\,
            I => \N__44568\
        );

    \I__9498\ : InMux
    port map (
            O => \N__44571\,
            I => \N__44565\
        );

    \I__9497\ : InMux
    port map (
            O => \N__44568\,
            I => \N__44562\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__44565\,
            I => \N__44557\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__44562\,
            I => \N__44557\
        );

    \I__9494\ : Span4Mux_h
    port map (
            O => \N__44557\,
            I => \N__44553\
        );

    \I__9493\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44550\
        );

    \I__9492\ : Odrv4
    port map (
            O => \N__44553\,
            I => n2928
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__44550\,
            I => n2928
        );

    \I__9490\ : CascadeMux
    port map (
            O => \N__44545\,
            I => \N__44541\
        );

    \I__9489\ : CascadeMux
    port map (
            O => \N__44544\,
            I => \N__44538\
        );

    \I__9488\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44535\
        );

    \I__9487\ : InMux
    port map (
            O => \N__44538\,
            I => \N__44532\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__44535\,
            I => \N__44529\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__44532\,
            I => \N__44523\
        );

    \I__9484\ : Span4Mux_h
    port map (
            O => \N__44529\,
            I => \N__44523\
        );

    \I__9483\ : InMux
    port map (
            O => \N__44528\,
            I => \N__44520\
        );

    \I__9482\ : Odrv4
    port map (
            O => \N__44523\,
            I => n2922
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__44520\,
            I => n2922
        );

    \I__9480\ : InMux
    port map (
            O => \N__44515\,
            I => \N__44512\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__44512\,
            I => \N__44509\
        );

    \I__9478\ : Span4Mux_h
    port map (
            O => \N__44509\,
            I => \N__44506\
        );

    \I__9477\ : Odrv4
    port map (
            O => \N__44506\,
            I => n2793
        );

    \I__9476\ : CascadeMux
    port map (
            O => \N__44503\,
            I => \N__44500\
        );

    \I__9475\ : InMux
    port map (
            O => \N__44500\,
            I => \N__44496\
        );

    \I__9474\ : CascadeMux
    port map (
            O => \N__44499\,
            I => \N__44493\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__44496\,
            I => \N__44490\
        );

    \I__9472\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44487\
        );

    \I__9471\ : Span4Mux_h
    port map (
            O => \N__44490\,
            I => \N__44483\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__44487\,
            I => \N__44480\
        );

    \I__9469\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44477\
        );

    \I__9468\ : Odrv4
    port map (
            O => \N__44483\,
            I => n2726
        );

    \I__9467\ : Odrv4
    port map (
            O => \N__44480\,
            I => n2726
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__44477\,
            I => n2726
        );

    \I__9465\ : CascadeMux
    port map (
            O => \N__44470\,
            I => \n2825_cascade_\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__44467\,
            I => \N__44464\
        );

    \I__9463\ : InMux
    port map (
            O => \N__44464\,
            I => \N__44461\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__44461\,
            I => \N__44457\
        );

    \I__9461\ : InMux
    port map (
            O => \N__44460\,
            I => \N__44453\
        );

    \I__9460\ : Span4Mux_v
    port map (
            O => \N__44457\,
            I => \N__44450\
        );

    \I__9459\ : InMux
    port map (
            O => \N__44456\,
            I => \N__44447\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__44453\,
            I => n2924
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__44450\,
            I => n2924
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__44447\,
            I => n2924
        );

    \I__9455\ : InMux
    port map (
            O => \N__44440\,
            I => \N__44437\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__44437\,
            I => \N__44434\
        );

    \I__9453\ : Odrv4
    port map (
            O => \N__44434\,
            I => n2796
        );

    \I__9452\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44427\
        );

    \I__9451\ : CascadeMux
    port map (
            O => \N__44430\,
            I => \N__44424\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__44427\,
            I => \N__44420\
        );

    \I__9449\ : InMux
    port map (
            O => \N__44424\,
            I => \N__44417\
        );

    \I__9448\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44414\
        );

    \I__9447\ : Span4Mux_h
    port map (
            O => \N__44420\,
            I => \N__44409\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__44417\,
            I => \N__44409\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__44414\,
            I => n2729
        );

    \I__9444\ : Odrv4
    port map (
            O => \N__44409\,
            I => n2729
        );

    \I__9443\ : InMux
    port map (
            O => \N__44404\,
            I => \N__44401\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__44401\,
            I => \N__44398\
        );

    \I__9441\ : Span4Mux_h
    port map (
            O => \N__44398\,
            I => \N__44395\
        );

    \I__9440\ : Odrv4
    port map (
            O => \N__44395\,
            I => n2800
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__44392\,
            I => \N__44389\
        );

    \I__9438\ : InMux
    port map (
            O => \N__44389\,
            I => \N__44386\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__44386\,
            I => \N__44382\
        );

    \I__9436\ : CascadeMux
    port map (
            O => \N__44385\,
            I => \N__44378\
        );

    \I__9435\ : Span4Mux_v
    port map (
            O => \N__44382\,
            I => \N__44375\
        );

    \I__9434\ : InMux
    port map (
            O => \N__44381\,
            I => \N__44372\
        );

    \I__9433\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44369\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__44375\,
            I => n2733
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__44372\,
            I => n2733
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__44369\,
            I => n2733
        );

    \I__9429\ : InMux
    port map (
            O => \N__44362\,
            I => \N__44359\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__44359\,
            I => \N__44356\
        );

    \I__9427\ : Span4Mux_h
    port map (
            O => \N__44356\,
            I => \N__44353\
        );

    \I__9426\ : Odrv4
    port map (
            O => \N__44353\,
            I => n2799
        );

    \I__9425\ : InMux
    port map (
            O => \N__44350\,
            I => \N__44347\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__44347\,
            I => \N__44343\
        );

    \I__9423\ : CascadeMux
    port map (
            O => \N__44346\,
            I => \N__44340\
        );

    \I__9422\ : Span4Mux_h
    port map (
            O => \N__44343\,
            I => \N__44337\
        );

    \I__9421\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44334\
        );

    \I__9420\ : Odrv4
    port map (
            O => \N__44337\,
            I => n2732
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__44334\,
            I => n2732
        );

    \I__9418\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44326\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__44326\,
            I => n14246
        );

    \I__9416\ : CascadeMux
    port map (
            O => \N__44323\,
            I => \n14248_cascade_\
        );

    \I__9415\ : CascadeMux
    port map (
            O => \N__44320\,
            I => \n14254_cascade_\
        );

    \I__9414\ : InMux
    port map (
            O => \N__44317\,
            I => \N__44314\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__44314\,
            I => n14266
        );

    \I__9412\ : CascadeMux
    port map (
            O => \N__44311\,
            I => \n2841_cascade_\
        );

    \I__9411\ : CascadeMux
    port map (
            O => \N__44308\,
            I => \N__44305\
        );

    \I__9410\ : InMux
    port map (
            O => \N__44305\,
            I => \N__44301\
        );

    \I__9409\ : CascadeMux
    port map (
            O => \N__44304\,
            I => \N__44298\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__44301\,
            I => \N__44295\
        );

    \I__9407\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44292\
        );

    \I__9406\ : Span4Mux_h
    port map (
            O => \N__44295\,
            I => \N__44287\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__44292\,
            I => \N__44287\
        );

    \I__9404\ : Span4Mux_v
    port map (
            O => \N__44287\,
            I => \N__44283\
        );

    \I__9403\ : InMux
    port map (
            O => \N__44286\,
            I => \N__44280\
        );

    \I__9402\ : Odrv4
    port map (
            O => \N__44283\,
            I => n2923
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__44280\,
            I => n2923
        );

    \I__9400\ : InMux
    port map (
            O => \N__44275\,
            I => \N__44271\
        );

    \I__9399\ : InMux
    port map (
            O => \N__44274\,
            I => \N__44267\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__44271\,
            I => \N__44264\
        );

    \I__9397\ : InMux
    port map (
            O => \N__44270\,
            I => \N__44261\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__44267\,
            I => \N__44256\
        );

    \I__9395\ : Span4Mux_s1_v
    port map (
            O => \N__44264\,
            I => \N__44256\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__44261\,
            I => pwm_counter_17
        );

    \I__9393\ : Odrv4
    port map (
            O => \N__44256\,
            I => pwm_counter_17
        );

    \I__9392\ : InMux
    port map (
            O => \N__44251\,
            I => \N__44247\
        );

    \I__9391\ : InMux
    port map (
            O => \N__44250\,
            I => \N__44243\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__44247\,
            I => \N__44240\
        );

    \I__9389\ : InMux
    port map (
            O => \N__44246\,
            I => \N__44237\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__44243\,
            I => \N__44234\
        );

    \I__9387\ : Span4Mux_h
    port map (
            O => \N__44240\,
            I => \N__44229\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__44237\,
            I => \N__44229\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__44234\,
            I => n2712
        );

    \I__9384\ : Odrv4
    port map (
            O => \N__44229\,
            I => n2712
        );

    \I__9383\ : CascadeMux
    port map (
            O => \N__44224\,
            I => \N__44221\
        );

    \I__9382\ : InMux
    port map (
            O => \N__44221\,
            I => \N__44218\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__44218\,
            I => \N__44215\
        );

    \I__9380\ : Span4Mux_h
    port map (
            O => \N__44215\,
            I => \N__44212\
        );

    \I__9379\ : Odrv4
    port map (
            O => \N__44212\,
            I => n2779
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__44209\,
            I => \n2811_cascade_\
        );

    \I__9377\ : InMux
    port map (
            O => \N__44206\,
            I => \N__44203\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__44203\,
            I => \N__44200\
        );

    \I__9375\ : Odrv12
    port map (
            O => \N__44200\,
            I => n2794
        );

    \I__9374\ : CascadeMux
    port map (
            O => \N__44197\,
            I => \N__44194\
        );

    \I__9373\ : InMux
    port map (
            O => \N__44194\,
            I => \N__44190\
        );

    \I__9372\ : CascadeMux
    port map (
            O => \N__44193\,
            I => \N__44186\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__44190\,
            I => \N__44183\
        );

    \I__9370\ : InMux
    port map (
            O => \N__44189\,
            I => \N__44180\
        );

    \I__9369\ : InMux
    port map (
            O => \N__44186\,
            I => \N__44177\
        );

    \I__9368\ : Span4Mux_h
    port map (
            O => \N__44183\,
            I => \N__44170\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__44180\,
            I => \N__44170\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__44177\,
            I => \N__44170\
        );

    \I__9365\ : Odrv4
    port map (
            O => \N__44170\,
            I => n2727
        );

    \I__9364\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44162\
        );

    \I__9363\ : InMux
    port map (
            O => \N__44166\,
            I => \N__44159\
        );

    \I__9362\ : InMux
    port map (
            O => \N__44165\,
            I => \N__44156\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__44162\,
            I => \N__44153\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__44159\,
            I => \N__44148\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__44156\,
            I => \N__44148\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__44153\,
            I => n2716
        );

    \I__9357\ : Odrv12
    port map (
            O => \N__44148\,
            I => n2716
        );

    \I__9356\ : CascadeMux
    port map (
            O => \N__44143\,
            I => \N__44140\
        );

    \I__9355\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44137\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__44137\,
            I => \N__44134\
        );

    \I__9353\ : Span4Mux_v
    port map (
            O => \N__44134\,
            I => \N__44131\
        );

    \I__9352\ : Odrv4
    port map (
            O => \N__44131\,
            I => n2783
        );

    \I__9351\ : InMux
    port map (
            O => \N__44128\,
            I => \N__44125\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__44125\,
            I => \N__44122\
        );

    \I__9349\ : Span4Mux_v
    port map (
            O => \N__44122\,
            I => \N__44119\
        );

    \I__9348\ : Odrv4
    port map (
            O => \N__44119\,
            I => n2782
        );

    \I__9347\ : CascadeMux
    port map (
            O => \N__44116\,
            I => \N__44112\
        );

    \I__9346\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44108\
        );

    \I__9345\ : InMux
    port map (
            O => \N__44112\,
            I => \N__44105\
        );

    \I__9344\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44102\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__44108\,
            I => \N__44097\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__44105\,
            I => \N__44097\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__44102\,
            I => \N__44094\
        );

    \I__9340\ : Span4Mux_h
    port map (
            O => \N__44097\,
            I => \N__44091\
        );

    \I__9339\ : Odrv4
    port map (
            O => \N__44094\,
            I => n2715
        );

    \I__9338\ : Odrv4
    port map (
            O => \N__44091\,
            I => n2715
        );

    \I__9337\ : CascadeMux
    port map (
            O => \N__44086\,
            I => \n2814_cascade_\
        );

    \I__9336\ : InMux
    port map (
            O => \N__44083\,
            I => \N__44080\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__44080\,
            I => n14260
        );

    \I__9334\ : InMux
    port map (
            O => \N__44077\,
            I => \N__44074\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__44074\,
            I => \N__44071\
        );

    \I__9332\ : Odrv4
    port map (
            O => \N__44071\,
            I => \pwm_setpoint_23_N_171_15\
        );

    \I__9331\ : InMux
    port map (
            O => \N__44068\,
            I => \N__44065\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__44065\,
            I => \pwm_setpoint_23_N_171_18\
        );

    \I__9329\ : InMux
    port map (
            O => \N__44062\,
            I => \N__44057\
        );

    \I__9328\ : InMux
    port map (
            O => \N__44061\,
            I => \N__44054\
        );

    \I__9327\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44051\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__44057\,
            I => \N__44046\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__44054\,
            I => \N__44046\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__44051\,
            I => pwm_counter_23
        );

    \I__9323\ : Odrv4
    port map (
            O => \N__44046\,
            I => pwm_counter_23
        );

    \I__9322\ : InMux
    port map (
            O => \N__44041\,
            I => \N__44038\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__44038\,
            I => \PWM.n28\
        );

    \I__9320\ : CascadeMux
    port map (
            O => \N__44035\,
            I => \N__44032\
        );

    \I__9319\ : InMux
    port map (
            O => \N__44032\,
            I => \N__44027\
        );

    \I__9318\ : InMux
    port map (
            O => \N__44031\,
            I => \N__44024\
        );

    \I__9317\ : InMux
    port map (
            O => \N__44030\,
            I => \N__44021\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__44027\,
            I => \N__44018\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__44024\,
            I => \N__44015\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__44021\,
            I => \N__44008\
        );

    \I__9313\ : Span4Mux_h
    port map (
            O => \N__44018\,
            I => \N__44008\
        );

    \I__9312\ : Span4Mux_s2_v
    port map (
            O => \N__44015\,
            I => \N__44008\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__44008\,
            I => pwm_counter_15
        );

    \I__9310\ : InMux
    port map (
            O => \N__44005\,
            I => \N__44001\
        );

    \I__9309\ : InMux
    port map (
            O => \N__44004\,
            I => \N__43997\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__44001\,
            I => \N__43994\
        );

    \I__9307\ : InMux
    port map (
            O => \N__44000\,
            I => \N__43991\
        );

    \I__9306\ : LocalMux
    port map (
            O => \N__43997\,
            I => \N__43984\
        );

    \I__9305\ : Span4Mux_v
    port map (
            O => \N__43994\,
            I => \N__43984\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__43991\,
            I => \N__43984\
        );

    \I__9303\ : Odrv4
    port map (
            O => \N__43984\,
            I => pwm_counter_18
        );

    \I__9302\ : InMux
    port map (
            O => \N__43981\,
            I => \N__43978\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__43978\,
            I => n37
        );

    \I__9300\ : InMux
    port map (
            O => \N__43975\,
            I => \N__43969\
        );

    \I__9299\ : InMux
    port map (
            O => \N__43974\,
            I => \N__43969\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__43969\,
            I => pwm_setpoint_18
        );

    \I__9297\ : CascadeMux
    port map (
            O => \N__43966\,
            I => \n37_cascade_\
        );

    \I__9296\ : InMux
    port map (
            O => \N__43963\,
            I => \N__43960\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__43960\,
            I => n14887
        );

    \I__9294\ : InMux
    port map (
            O => \N__43957\,
            I => \N__43954\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__43954\,
            I => \pwm_setpoint_23_N_171_22\
        );

    \I__9292\ : InMux
    port map (
            O => \N__43951\,
            I => \N__43945\
        );

    \I__9291\ : InMux
    port map (
            O => \N__43950\,
            I => \N__43945\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__43945\,
            I => \N__43942\
        );

    \I__9289\ : Odrv12
    port map (
            O => \N__43942\,
            I => pwm_setpoint_22
        );

    \I__9288\ : InMux
    port map (
            O => \N__43939\,
            I => \N__43936\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__43936\,
            I => \N__43933\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__43933\,
            I => \pwm_setpoint_23_N_171_17\
        );

    \I__9285\ : InMux
    port map (
            O => \N__43930\,
            I => \N__43927\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__43927\,
            I => n14870
        );

    \I__9283\ : InMux
    port map (
            O => \N__43924\,
            I => \N__43921\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__43921\,
            I => n14832
        );

    \I__9281\ : InMux
    port map (
            O => \N__43918\,
            I => n12064
        );

    \I__9280\ : InMux
    port map (
            O => \N__43915\,
            I => \bfn_13_30_0_\
        );

    \I__9279\ : InMux
    port map (
            O => \N__43912\,
            I => n12066
        );

    \I__9278\ : InMux
    port map (
            O => \N__43909\,
            I => n12067
        );

    \I__9277\ : InMux
    port map (
            O => \N__43906\,
            I => \N__43903\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__43903\,
            I => \pwm_setpoint_23_N_171_19\
        );

    \I__9275\ : InMux
    port map (
            O => \N__43900\,
            I => n12068
        );

    \I__9274\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43894\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__43894\,
            I => \pwm_setpoint_23_N_171_20\
        );

    \I__9272\ : InMux
    port map (
            O => \N__43891\,
            I => n12069
        );

    \I__9271\ : InMux
    port map (
            O => \N__43888\,
            I => \N__43885\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__43885\,
            I => \N__43882\
        );

    \I__9269\ : Span4Mux_v
    port map (
            O => \N__43882\,
            I => \N__43879\
        );

    \I__9268\ : Odrv4
    port map (
            O => \N__43879\,
            I => n4_adj_570
        );

    \I__9267\ : InMux
    port map (
            O => \N__43876\,
            I => \N__43873\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__43873\,
            I => \N__43870\
        );

    \I__9265\ : Span4Mux_v
    port map (
            O => \N__43870\,
            I => \N__43867\
        );

    \I__9264\ : Odrv4
    port map (
            O => \N__43867\,
            I => \pwm_setpoint_23_N_171_21\
        );

    \I__9263\ : InMux
    port map (
            O => \N__43864\,
            I => n12070
        );

    \I__9262\ : InMux
    port map (
            O => \N__43861\,
            I => n12071
        );

    \I__9261\ : InMux
    port map (
            O => \N__43858\,
            I => n12072
        );

    \I__9260\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43852\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__43852\,
            I => \N__43849\
        );

    \I__9258\ : Odrv4
    port map (
            O => \N__43849\,
            I => pwm_setpoint_23
        );

    \I__9257\ : InMux
    port map (
            O => \N__43846\,
            I => \N__43843\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__43843\,
            I => n18_adj_584
        );

    \I__9255\ : InMux
    port map (
            O => \N__43840\,
            I => n12056
        );

    \I__9254\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43834\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__43834\,
            I => \pwm_setpoint_23_N_171_8\
        );

    \I__9252\ : InMux
    port map (
            O => \N__43831\,
            I => \bfn_13_29_0_\
        );

    \I__9251\ : InMux
    port map (
            O => \N__43828\,
            I => n12058
        );

    \I__9250\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43822\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43819\
        );

    \I__9248\ : Odrv4
    port map (
            O => \N__43819\,
            I => n15_adj_581
        );

    \I__9247\ : InMux
    port map (
            O => \N__43816\,
            I => \N__43813\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__43813\,
            I => \pwm_setpoint_23_N_171_10\
        );

    \I__9245\ : InMux
    port map (
            O => \N__43810\,
            I => n12059
        );

    \I__9244\ : InMux
    port map (
            O => \N__43807\,
            I => \N__43804\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__43804\,
            I => \N__43801\
        );

    \I__9242\ : Odrv4
    port map (
            O => \N__43801\,
            I => n14_adj_580
        );

    \I__9241\ : InMux
    port map (
            O => \N__43798\,
            I => \N__43795\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__43795\,
            I => \pwm_setpoint_23_N_171_11\
        );

    \I__9239\ : InMux
    port map (
            O => \N__43792\,
            I => n12060
        );

    \I__9238\ : CascadeMux
    port map (
            O => \N__43789\,
            I => \N__43786\
        );

    \I__9237\ : InMux
    port map (
            O => \N__43786\,
            I => \N__43783\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__43783\,
            I => \pwm_setpoint_23_N_171_12\
        );

    \I__9235\ : InMux
    port map (
            O => \N__43780\,
            I => n12061
        );

    \I__9234\ : InMux
    port map (
            O => \N__43777\,
            I => n12062
        );

    \I__9233\ : InMux
    port map (
            O => \N__43774\,
            I => \N__43771\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__43771\,
            I => \N__43768\
        );

    \I__9231\ : Odrv4
    port map (
            O => \N__43768\,
            I => n11_adj_577
        );

    \I__9230\ : InMux
    port map (
            O => \N__43765\,
            I => n12063
        );

    \I__9229\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43759\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__43759\,
            I => n25_adj_591
        );

    \I__9227\ : InMux
    port map (
            O => \N__43756\,
            I => \bfn_13_28_0_\
        );

    \I__9226\ : InMux
    port map (
            O => \N__43753\,
            I => n12050
        );

    \I__9225\ : InMux
    port map (
            O => \N__43750\,
            I => \N__43747\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__43747\,
            I => n23_adj_589
        );

    \I__9223\ : InMux
    port map (
            O => \N__43744\,
            I => \N__43741\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__43741\,
            I => \pwm_setpoint_23_N_171_2\
        );

    \I__9221\ : InMux
    port map (
            O => \N__43738\,
            I => n12051
        );

    \I__9220\ : InMux
    port map (
            O => \N__43735\,
            I => \N__43732\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__43732\,
            I => \pwm_setpoint_23_N_171_3\
        );

    \I__9218\ : InMux
    port map (
            O => \N__43729\,
            I => n12052
        );

    \I__9217\ : InMux
    port map (
            O => \N__43726\,
            I => \N__43723\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__43723\,
            I => \N__43720\
        );

    \I__9215\ : Span4Mux_v
    port map (
            O => \N__43720\,
            I => \N__43717\
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__43717\,
            I => n21_adj_587
        );

    \I__9213\ : InMux
    port map (
            O => \N__43714\,
            I => \N__43711\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__43711\,
            I => \pwm_setpoint_23_N_171_4\
        );

    \I__9211\ : InMux
    port map (
            O => \N__43708\,
            I => n12053
        );

    \I__9210\ : InMux
    port map (
            O => \N__43705\,
            I => \N__43702\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__43702\,
            I => n20_adj_586
        );

    \I__9208\ : InMux
    port map (
            O => \N__43699\,
            I => \N__43696\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__43696\,
            I => \N__43693\
        );

    \I__9206\ : Odrv4
    port map (
            O => \N__43693\,
            I => \pwm_setpoint_23_N_171_5\
        );

    \I__9205\ : InMux
    port map (
            O => \N__43690\,
            I => n12054
        );

    \I__9204\ : InMux
    port map (
            O => \N__43687\,
            I => \N__43684\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__43684\,
            I => n19_adj_585
        );

    \I__9202\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43678\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__43678\,
            I => \pwm_setpoint_23_N_171_6\
        );

    \I__9200\ : InMux
    port map (
            O => \N__43675\,
            I => n12055
        );

    \I__9199\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43669\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__43669\,
            I => \N__43665\
        );

    \I__9197\ : CascadeMux
    port map (
            O => \N__43668\,
            I => \N__43662\
        );

    \I__9196\ : Span4Mux_v
    port map (
            O => \N__43665\,
            I => \N__43658\
        );

    \I__9195\ : InMux
    port map (
            O => \N__43662\,
            I => \N__43655\
        );

    \I__9194\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43652\
        );

    \I__9193\ : Sp12to4
    port map (
            O => \N__43658\,
            I => \N__43647\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__43655\,
            I => \N__43647\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__43652\,
            I => n3206
        );

    \I__9190\ : Odrv12
    port map (
            O => \N__43647\,
            I => n3206
        );

    \I__9189\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43639\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__43639\,
            I => \N__43636\
        );

    \I__9187\ : Span4Mux_h
    port map (
            O => \N__43636\,
            I => \N__43633\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__43633\,
            I => n3273
        );

    \I__9185\ : InMux
    port map (
            O => \N__43630\,
            I => n12549
        );

    \I__9184\ : InMux
    port map (
            O => \N__43627\,
            I => \N__43624\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__43624\,
            I => \N__43621\
        );

    \I__9182\ : Span4Mux_h
    port map (
            O => \N__43621\,
            I => \N__43616\
        );

    \I__9181\ : InMux
    port map (
            O => \N__43620\,
            I => \N__43611\
        );

    \I__9180\ : InMux
    port map (
            O => \N__43619\,
            I => \N__43611\
        );

    \I__9179\ : Odrv4
    port map (
            O => \N__43616\,
            I => n3205
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__43611\,
            I => n3205
        );

    \I__9177\ : InMux
    port map (
            O => \N__43606\,
            I => \N__43603\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__43603\,
            I => \N__43600\
        );

    \I__9175\ : Span4Mux_v
    port map (
            O => \N__43600\,
            I => \N__43597\
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__43597\,
            I => n3272
        );

    \I__9173\ : InMux
    port map (
            O => \N__43594\,
            I => n12550
        );

    \I__9172\ : InMux
    port map (
            O => \N__43591\,
            I => \N__43588\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__43588\,
            I => \N__43584\
        );

    \I__9170\ : InMux
    port map (
            O => \N__43587\,
            I => \N__43581\
        );

    \I__9169\ : Span12Mux_s7_v
    port map (
            O => \N__43584\,
            I => \N__43578\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__43581\,
            I => n15163
        );

    \I__9167\ : Odrv12
    port map (
            O => \N__43578\,
            I => n15163
        );

    \I__9166\ : InMux
    port map (
            O => \N__43573\,
            I => n12551
        );

    \I__9165\ : InMux
    port map (
            O => \N__43570\,
            I => \N__43567\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__43567\,
            I => \N__43564\
        );

    \I__9163\ : Span4Mux_h
    port map (
            O => \N__43564\,
            I => \N__43561\
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__43561\,
            I => n14461
        );

    \I__9161\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43555\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__43555\,
            I => \N__43552\
        );

    \I__9159\ : Span4Mux_v
    port map (
            O => \N__43552\,
            I => \N__43549\
        );

    \I__9158\ : Odrv4
    port map (
            O => \N__43549\,
            I => encoder0_position_scaled_3
        );

    \I__9157\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43541\
        );

    \I__9156\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43538\
        );

    \I__9155\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43535\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__43541\,
            I => dti_counter_2
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__43538\,
            I => dti_counter_2
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__43535\,
            I => dti_counter_2
        );

    \I__9151\ : CascadeMux
    port map (
            O => \N__43528\,
            I => \N__43524\
        );

    \I__9150\ : InMux
    port map (
            O => \N__43527\,
            I => \N__43520\
        );

    \I__9149\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43517\
        );

    \I__9148\ : InMux
    port map (
            O => \N__43523\,
            I => \N__43514\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__43520\,
            I => dti_counter_1
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__43517\,
            I => dti_counter_1
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__43514\,
            I => dti_counter_1
        );

    \I__9144\ : InMux
    port map (
            O => \N__43507\,
            I => \N__43504\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__43504\,
            I => n10_adj_680
        );

    \I__9142\ : InMux
    port map (
            O => \N__43501\,
            I => \N__43498\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__43498\,
            I => n3281
        );

    \I__9140\ : InMux
    port map (
            O => \N__43495\,
            I => n12541
        );

    \I__9139\ : InMux
    port map (
            O => \N__43492\,
            I => \N__43489\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__43489\,
            I => n3280
        );

    \I__9137\ : InMux
    port map (
            O => \N__43486\,
            I => n12542
        );

    \I__9136\ : InMux
    port map (
            O => \N__43483\,
            I => \N__43479\
        );

    \I__9135\ : InMux
    port map (
            O => \N__43482\,
            I => \N__43475\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__43479\,
            I => \N__43472\
        );

    \I__9133\ : InMux
    port map (
            O => \N__43478\,
            I => \N__43469\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__43475\,
            I => \N__43466\
        );

    \I__9131\ : Span4Mux_v
    port map (
            O => \N__43472\,
            I => \N__43463\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__43469\,
            I => \N__43460\
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__43466\,
            I => n3212
        );

    \I__9128\ : Odrv4
    port map (
            O => \N__43463\,
            I => n3212
        );

    \I__9127\ : Odrv4
    port map (
            O => \N__43460\,
            I => n3212
        );

    \I__9126\ : InMux
    port map (
            O => \N__43453\,
            I => \N__43450\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__43450\,
            I => \N__43447\
        );

    \I__9124\ : Odrv4
    port map (
            O => \N__43447\,
            I => n3279
        );

    \I__9123\ : InMux
    port map (
            O => \N__43444\,
            I => n12543
        );

    \I__9122\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43437\
        );

    \I__9121\ : InMux
    port map (
            O => \N__43440\,
            I => \N__43434\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__43437\,
            I => \N__43430\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__43434\,
            I => \N__43427\
        );

    \I__9118\ : InMux
    port map (
            O => \N__43433\,
            I => \N__43424\
        );

    \I__9117\ : Odrv4
    port map (
            O => \N__43430\,
            I => n3211
        );

    \I__9116\ : Odrv4
    port map (
            O => \N__43427\,
            I => n3211
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__43424\,
            I => n3211
        );

    \I__9114\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43414\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__43414\,
            I => \N__43411\
        );

    \I__9112\ : Span4Mux_v
    port map (
            O => \N__43411\,
            I => \N__43408\
        );

    \I__9111\ : Odrv4
    port map (
            O => \N__43408\,
            I => n3278
        );

    \I__9110\ : InMux
    port map (
            O => \N__43405\,
            I => \bfn_13_26_0_\
        );

    \I__9109\ : InMux
    port map (
            O => \N__43402\,
            I => \N__43398\
        );

    \I__9108\ : CascadeMux
    port map (
            O => \N__43401\,
            I => \N__43395\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__43398\,
            I => \N__43391\
        );

    \I__9106\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43388\
        );

    \I__9105\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43385\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__43391\,
            I => \N__43380\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__43388\,
            I => \N__43380\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__43385\,
            I => n3210
        );

    \I__9101\ : Odrv4
    port map (
            O => \N__43380\,
            I => n3210
        );

    \I__9100\ : InMux
    port map (
            O => \N__43375\,
            I => \N__43372\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__43372\,
            I => \N__43369\
        );

    \I__9098\ : Span4Mux_v
    port map (
            O => \N__43369\,
            I => \N__43366\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__43366\,
            I => n3277
        );

    \I__9096\ : InMux
    port map (
            O => \N__43363\,
            I => n12545
        );

    \I__9095\ : InMux
    port map (
            O => \N__43360\,
            I => \N__43357\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__43357\,
            I => \N__43354\
        );

    \I__9093\ : Span4Mux_h
    port map (
            O => \N__43354\,
            I => \N__43351\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__43351\,
            I => n3276
        );

    \I__9091\ : InMux
    port map (
            O => \N__43348\,
            I => n12546
        );

    \I__9090\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43342\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__43342\,
            I => \N__43338\
        );

    \I__9088\ : InMux
    port map (
            O => \N__43341\,
            I => \N__43334\
        );

    \I__9087\ : Span4Mux_h
    port map (
            O => \N__43338\,
            I => \N__43331\
        );

    \I__9086\ : InMux
    port map (
            O => \N__43337\,
            I => \N__43328\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__43334\,
            I => n3208
        );

    \I__9084\ : Odrv4
    port map (
            O => \N__43331\,
            I => n3208
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__43328\,
            I => n3208
        );

    \I__9082\ : InMux
    port map (
            O => \N__43321\,
            I => \N__43318\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__43318\,
            I => \N__43315\
        );

    \I__9080\ : Span4Mux_h
    port map (
            O => \N__43315\,
            I => \N__43312\
        );

    \I__9079\ : Odrv4
    port map (
            O => \N__43312\,
            I => n3275
        );

    \I__9078\ : InMux
    port map (
            O => \N__43309\,
            I => n12547
        );

    \I__9077\ : InMux
    port map (
            O => \N__43306\,
            I => \N__43303\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__43303\,
            I => \N__43299\
        );

    \I__9075\ : InMux
    port map (
            O => \N__43302\,
            I => \N__43295\
        );

    \I__9074\ : Span4Mux_h
    port map (
            O => \N__43299\,
            I => \N__43292\
        );

    \I__9073\ : InMux
    port map (
            O => \N__43298\,
            I => \N__43289\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__43295\,
            I => n3207
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__43292\,
            I => n3207
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__43289\,
            I => n3207
        );

    \I__9069\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43279\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__43279\,
            I => \N__43276\
        );

    \I__9067\ : Span4Mux_h
    port map (
            O => \N__43276\,
            I => \N__43273\
        );

    \I__9066\ : Odrv4
    port map (
            O => \N__43273\,
            I => n3274
        );

    \I__9065\ : InMux
    port map (
            O => \N__43270\,
            I => n12548
        );

    \I__9064\ : InMux
    port map (
            O => \N__43267\,
            I => n12533
        );

    \I__9063\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43261\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__43261\,
            I => n3288
        );

    \I__9061\ : InMux
    port map (
            O => \N__43258\,
            I => n12534
        );

    \I__9060\ : InMux
    port map (
            O => \N__43255\,
            I => n12535
        );

    \I__9059\ : InMux
    port map (
            O => \N__43252\,
            I => \bfn_13_25_0_\
        );

    \I__9058\ : InMux
    port map (
            O => \N__43249\,
            I => \N__43246\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__43246\,
            I => n3285
        );

    \I__9056\ : InMux
    port map (
            O => \N__43243\,
            I => n12537
        );

    \I__9055\ : CascadeMux
    port map (
            O => \N__43240\,
            I => \N__43237\
        );

    \I__9054\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43233\
        );

    \I__9053\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43230\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__43233\,
            I => \N__43224\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__43230\,
            I => \N__43224\
        );

    \I__9050\ : InMux
    port map (
            O => \N__43229\,
            I => \N__43221\
        );

    \I__9049\ : Odrv4
    port map (
            O => \N__43224\,
            I => n3217
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__43221\,
            I => n3217
        );

    \I__9047\ : InMux
    port map (
            O => \N__43216\,
            I => \N__43213\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__43213\,
            I => n3284
        );

    \I__9045\ : InMux
    port map (
            O => \N__43210\,
            I => n12538
        );

    \I__9044\ : InMux
    port map (
            O => \N__43207\,
            I => \N__43204\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__43204\,
            I => \N__43200\
        );

    \I__9042\ : InMux
    port map (
            O => \N__43203\,
            I => \N__43196\
        );

    \I__9041\ : Span4Mux_v
    port map (
            O => \N__43200\,
            I => \N__43193\
        );

    \I__9040\ : InMux
    port map (
            O => \N__43199\,
            I => \N__43190\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__43196\,
            I => n3216
        );

    \I__9038\ : Odrv4
    port map (
            O => \N__43193\,
            I => n3216
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__43190\,
            I => n3216
        );

    \I__9036\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43180\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43177\
        );

    \I__9034\ : Odrv4
    port map (
            O => \N__43177\,
            I => n3283
        );

    \I__9033\ : InMux
    port map (
            O => \N__43174\,
            I => n12539
        );

    \I__9032\ : InMux
    port map (
            O => \N__43171\,
            I => \N__43168\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__43168\,
            I => \N__43163\
        );

    \I__9030\ : InMux
    port map (
            O => \N__43167\,
            I => \N__43160\
        );

    \I__9029\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43157\
        );

    \I__9028\ : Span4Mux_v
    port map (
            O => \N__43163\,
            I => \N__43152\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__43160\,
            I => \N__43152\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__43157\,
            I => \N__43149\
        );

    \I__9025\ : Span4Mux_v
    port map (
            O => \N__43152\,
            I => \N__43146\
        );

    \I__9024\ : Odrv12
    port map (
            O => \N__43149\,
            I => n3215
        );

    \I__9023\ : Odrv4
    port map (
            O => \N__43146\,
            I => n3215
        );

    \I__9022\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43138\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__43138\,
            I => n3282
        );

    \I__9020\ : InMux
    port map (
            O => \N__43135\,
            I => n12540
        );

    \I__9019\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43127\
        );

    \I__9018\ : InMux
    port map (
            O => \N__43131\,
            I => \N__43124\
        );

    \I__9017\ : InMux
    port map (
            O => \N__43130\,
            I => \N__43121\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__43127\,
            I => \N__43118\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__43124\,
            I => n3214
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__43121\,
            I => n3214
        );

    \I__9013\ : Odrv4
    port map (
            O => \N__43118\,
            I => n3214
        );

    \I__9012\ : InMux
    port map (
            O => \N__43111\,
            I => \N__43108\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__43108\,
            I => n3298
        );

    \I__9010\ : CascadeMux
    port map (
            O => \N__43105\,
            I => \N__43101\
        );

    \I__9009\ : InMux
    port map (
            O => \N__43104\,
            I => \N__43098\
        );

    \I__9008\ : InMux
    port map (
            O => \N__43101\,
            I => \N__43095\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__43098\,
            I => \N__43091\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__43095\,
            I => \N__43088\
        );

    \I__9005\ : InMux
    port map (
            O => \N__43094\,
            I => \N__43085\
        );

    \I__9004\ : Odrv4
    port map (
            O => \N__43091\,
            I => n3230
        );

    \I__9003\ : Odrv12
    port map (
            O => \N__43088\,
            I => n3230
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__43085\,
            I => n3230
        );

    \I__9001\ : InMux
    port map (
            O => \N__43078\,
            I => \N__43075\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__43075\,
            I => \N__43072\
        );

    \I__8999\ : Span4Mux_h
    port map (
            O => \N__43072\,
            I => \N__43069\
        );

    \I__8998\ : Odrv4
    port map (
            O => \N__43069\,
            I => n14697
        );

    \I__8997\ : InMux
    port map (
            O => \N__43066\,
            I => n12525
        );

    \I__8996\ : InMux
    port map (
            O => \N__43063\,
            I => n12526
        );

    \I__8995\ : InMux
    port map (
            O => \N__43060\,
            I => n12527
        );

    \I__8994\ : InMux
    port map (
            O => \N__43057\,
            I => \bfn_13_24_0_\
        );

    \I__8993\ : InMux
    port map (
            O => \N__43054\,
            I => \N__43051\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__43051\,
            I => n3293
        );

    \I__8991\ : InMux
    port map (
            O => \N__43048\,
            I => n12529
        );

    \I__8990\ : InMux
    port map (
            O => \N__43045\,
            I => n12530
        );

    \I__8989\ : CascadeMux
    port map (
            O => \N__43042\,
            I => \N__43039\
        );

    \I__8988\ : InMux
    port map (
            O => \N__43039\,
            I => \N__43036\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__43036\,
            I => n3291
        );

    \I__8986\ : InMux
    port map (
            O => \N__43033\,
            I => n12531
        );

    \I__8985\ : CascadeMux
    port map (
            O => \N__43030\,
            I => \N__43027\
        );

    \I__8984\ : InMux
    port map (
            O => \N__43027\,
            I => \N__43024\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__43024\,
            I => n3290
        );

    \I__8982\ : InMux
    port map (
            O => \N__43021\,
            I => n12532
        );

    \I__8981\ : CascadeMux
    port map (
            O => \N__43018\,
            I => \n3014_cascade_\
        );

    \I__8980\ : InMux
    port map (
            O => \N__43015\,
            I => \N__43012\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__43012\,
            I => n14408
        );

    \I__8978\ : InMux
    port map (
            O => \N__43009\,
            I => \N__43006\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__43006\,
            I => \N__42990\
        );

    \I__8976\ : InMux
    port map (
            O => \N__43005\,
            I => \N__42981\
        );

    \I__8975\ : InMux
    port map (
            O => \N__43004\,
            I => \N__42981\
        );

    \I__8974\ : InMux
    port map (
            O => \N__43003\,
            I => \N__42981\
        );

    \I__8973\ : InMux
    port map (
            O => \N__43002\,
            I => \N__42981\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__43001\,
            I => \N__42976\
        );

    \I__8971\ : CascadeMux
    port map (
            O => \N__43000\,
            I => \N__42972\
        );

    \I__8970\ : CascadeMux
    port map (
            O => \N__42999\,
            I => \N__42968\
        );

    \I__8969\ : CascadeMux
    port map (
            O => \N__42998\,
            I => \N__42965\
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__42997\,
            I => \N__42957\
        );

    \I__8967\ : CascadeMux
    port map (
            O => \N__42996\,
            I => \N__42954\
        );

    \I__8966\ : CascadeMux
    port map (
            O => \N__42995\,
            I => \N__42950\
        );

    \I__8965\ : CascadeMux
    port map (
            O => \N__42994\,
            I => \N__42947\
        );

    \I__8964\ : CascadeMux
    port map (
            O => \N__42993\,
            I => \N__42942\
        );

    \I__8963\ : Span4Mux_v
    port map (
            O => \N__42990\,
            I => \N__42937\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__42981\,
            I => \N__42934\
        );

    \I__8961\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42931\
        );

    \I__8960\ : InMux
    port map (
            O => \N__42979\,
            I => \N__42920\
        );

    \I__8959\ : InMux
    port map (
            O => \N__42976\,
            I => \N__42920\
        );

    \I__8958\ : InMux
    port map (
            O => \N__42975\,
            I => \N__42920\
        );

    \I__8957\ : InMux
    port map (
            O => \N__42972\,
            I => \N__42920\
        );

    \I__8956\ : InMux
    port map (
            O => \N__42971\,
            I => \N__42920\
        );

    \I__8955\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42913\
        );

    \I__8954\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42913\
        );

    \I__8953\ : InMux
    port map (
            O => \N__42964\,
            I => \N__42913\
        );

    \I__8952\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42906\
        );

    \I__8951\ : InMux
    port map (
            O => \N__42962\,
            I => \N__42906\
        );

    \I__8950\ : InMux
    port map (
            O => \N__42961\,
            I => \N__42906\
        );

    \I__8949\ : InMux
    port map (
            O => \N__42960\,
            I => \N__42897\
        );

    \I__8948\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42897\
        );

    \I__8947\ : InMux
    port map (
            O => \N__42954\,
            I => \N__42897\
        );

    \I__8946\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42897\
        );

    \I__8945\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42888\
        );

    \I__8944\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42888\
        );

    \I__8943\ : InMux
    port map (
            O => \N__42946\,
            I => \N__42888\
        );

    \I__8942\ : InMux
    port map (
            O => \N__42945\,
            I => \N__42888\
        );

    \I__8941\ : InMux
    port map (
            O => \N__42942\,
            I => \N__42881\
        );

    \I__8940\ : InMux
    port map (
            O => \N__42941\,
            I => \N__42881\
        );

    \I__8939\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42881\
        );

    \I__8938\ : Odrv4
    port map (
            O => \N__42937\,
            I => n2940
        );

    \I__8937\ : Odrv4
    port map (
            O => \N__42934\,
            I => n2940
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__42931\,
            I => n2940
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__42920\,
            I => n2940
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__42913\,
            I => n2940
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__42906\,
            I => n2940
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__42897\,
            I => n2940
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__42888\,
            I => n2940
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__42881\,
            I => n2940
        );

    \I__8929\ : InMux
    port map (
            O => \N__42862\,
            I => \N__42859\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__42859\,
            I => \N__42856\
        );

    \I__8927\ : Odrv4
    port map (
            O => \N__42856\,
            I => n2989
        );

    \I__8926\ : CascadeMux
    port map (
            O => \N__42853\,
            I => \n3021_cascade_\
        );

    \I__8925\ : InMux
    port map (
            O => \N__42850\,
            I => \N__42846\
        );

    \I__8924\ : InMux
    port map (
            O => \N__42849\,
            I => \N__42843\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__42846\,
            I => \N__42840\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__42843\,
            I => \N__42837\
        );

    \I__8921\ : Span4Mux_v
    port map (
            O => \N__42840\,
            I => \N__42834\
        );

    \I__8920\ : Span4Mux_v
    port map (
            O => \N__42837\,
            I => \N__42829\
        );

    \I__8919\ : Span4Mux_h
    port map (
            O => \N__42834\,
            I => \N__42829\
        );

    \I__8918\ : Span4Mux_h
    port map (
            O => \N__42829\,
            I => \N__42826\
        );

    \I__8917\ : Odrv4
    port map (
            O => \N__42826\,
            I => n319
        );

    \I__8916\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42819\
        );

    \I__8915\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42815\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__42819\,
            I => \N__42812\
        );

    \I__8913\ : InMux
    port map (
            O => \N__42818\,
            I => \N__42809\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__42815\,
            I => \N__42806\
        );

    \I__8911\ : Span4Mux_v
    port map (
            O => \N__42812\,
            I => \N__42803\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__42809\,
            I => \N__42800\
        );

    \I__8909\ : Span4Mux_h
    port map (
            O => \N__42806\,
            I => \N__42797\
        );

    \I__8908\ : Span4Mux_h
    port map (
            O => \N__42803\,
            I => \N__42792\
        );

    \I__8907\ : Span4Mux_v
    port map (
            O => \N__42800\,
            I => \N__42792\
        );

    \I__8906\ : Odrv4
    port map (
            O => \N__42797\,
            I => n318
        );

    \I__8905\ : Odrv4
    port map (
            O => \N__42792\,
            I => n318
        );

    \I__8904\ : CascadeMux
    port map (
            O => \N__42787\,
            I => \N__42784\
        );

    \I__8903\ : InMux
    port map (
            O => \N__42784\,
            I => \N__42781\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__42781\,
            I => \N__42778\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__42778\,
            I => \N__42775\
        );

    \I__8900\ : Odrv4
    port map (
            O => \N__42775\,
            I => n3301
        );

    \I__8899\ : InMux
    port map (
            O => \N__42772\,
            I => n12521
        );

    \I__8898\ : InMux
    port map (
            O => \N__42769\,
            I => \N__42766\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__42766\,
            I => \N__42762\
        );

    \I__8896\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42758\
        );

    \I__8895\ : Span4Mux_h
    port map (
            O => \N__42762\,
            I => \N__42755\
        );

    \I__8894\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42752\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__42758\,
            I => n3233
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__42755\,
            I => n3233
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__42752\,
            I => n3233
        );

    \I__8890\ : InMux
    port map (
            O => \N__42745\,
            I => \N__42742\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__42742\,
            I => \N__42739\
        );

    \I__8888\ : Span4Mux_v
    port map (
            O => \N__42739\,
            I => \N__42736\
        );

    \I__8887\ : Span4Mux_h
    port map (
            O => \N__42736\,
            I => \N__42733\
        );

    \I__8886\ : Odrv4
    port map (
            O => \N__42733\,
            I => n3300
        );

    \I__8885\ : InMux
    port map (
            O => \N__42730\,
            I => n12522
        );

    \I__8884\ : InMux
    port map (
            O => \N__42727\,
            I => \N__42724\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__42724\,
            I => \N__42720\
        );

    \I__8882\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42717\
        );

    \I__8881\ : Span4Mux_v
    port map (
            O => \N__42720\,
            I => \N__42714\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__42717\,
            I => \N__42711\
        );

    \I__8879\ : Odrv4
    port map (
            O => \N__42714\,
            I => n3232
        );

    \I__8878\ : Odrv12
    port map (
            O => \N__42711\,
            I => n3232
        );

    \I__8877\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42703\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__42703\,
            I => \N__42700\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__42700\,
            I => \N__42697\
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__42697\,
            I => n3299
        );

    \I__8873\ : InMux
    port map (
            O => \N__42694\,
            I => n12523
        );

    \I__8872\ : InMux
    port map (
            O => \N__42691\,
            I => \N__42688\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__42688\,
            I => \N__42684\
        );

    \I__8870\ : InMux
    port map (
            O => \N__42687\,
            I => \N__42680\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__42684\,
            I => \N__42677\
        );

    \I__8868\ : InMux
    port map (
            O => \N__42683\,
            I => \N__42674\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__42680\,
            I => n3231
        );

    \I__8866\ : Odrv4
    port map (
            O => \N__42677\,
            I => n3231
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__42674\,
            I => n3231
        );

    \I__8864\ : InMux
    port map (
            O => \N__42667\,
            I => n12524
        );

    \I__8863\ : InMux
    port map (
            O => \N__42664\,
            I => \N__42661\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__42661\,
            I => \N__42658\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__42658\,
            I => \N__42655\
        );

    \I__8860\ : Odrv4
    port map (
            O => \N__42655\,
            I => n2992
        );

    \I__8859\ : InMux
    port map (
            O => \N__42652\,
            I => \N__42649\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__42649\,
            I => \N__42646\
        );

    \I__8857\ : Span4Mux_v
    port map (
            O => \N__42646\,
            I => \N__42643\
        );

    \I__8856\ : Odrv4
    port map (
            O => \N__42643\,
            I => n2991
        );

    \I__8855\ : CascadeMux
    port map (
            O => \N__42640\,
            I => \n3023_cascade_\
        );

    \I__8854\ : InMux
    port map (
            O => \N__42637\,
            I => \N__42634\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__42634\,
            I => n14320
        );

    \I__8852\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42628\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__42628\,
            I => \N__42625\
        );

    \I__8850\ : Odrv12
    port map (
            O => \N__42625\,
            I => n2995
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__42622\,
            I => \N__42619\
        );

    \I__8848\ : InMux
    port map (
            O => \N__42619\,
            I => \N__42616\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__42616\,
            I => \N__42613\
        );

    \I__8846\ : Span4Mux_h
    port map (
            O => \N__42613\,
            I => \N__42610\
        );

    \I__8845\ : Odrv4
    port map (
            O => \N__42610\,
            I => n2994
        );

    \I__8844\ : InMux
    port map (
            O => \N__42607\,
            I => \N__42603\
        );

    \I__8843\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42600\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__42603\,
            I => \N__42595\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__42600\,
            I => \N__42595\
        );

    \I__8840\ : Span4Mux_h
    port map (
            O => \N__42595\,
            I => \N__42591\
        );

    \I__8839\ : InMux
    port map (
            O => \N__42594\,
            I => \N__42588\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__42591\,
            I => n2913
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__42588\,
            I => n2913
        );

    \I__8836\ : InMux
    port map (
            O => \N__42583\,
            I => \N__42580\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__42580\,
            I => \N__42577\
        );

    \I__8834\ : Odrv12
    port map (
            O => \N__42577\,
            I => n2990
        );

    \I__8833\ : CascadeMux
    port map (
            O => \N__42574\,
            I => \N__42571\
        );

    \I__8832\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42568\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__42568\,
            I => \N__42565\
        );

    \I__8830\ : Span4Mux_h
    port map (
            O => \N__42565\,
            I => \N__42562\
        );

    \I__8829\ : Odrv4
    port map (
            O => \N__42562\,
            I => n2982
        );

    \I__8828\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42555\
        );

    \I__8827\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42552\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__42555\,
            I => \N__42549\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__42552\,
            I => \N__42545\
        );

    \I__8824\ : Span4Mux_v
    port map (
            O => \N__42549\,
            I => \N__42542\
        );

    \I__8823\ : InMux
    port map (
            O => \N__42548\,
            I => \N__42539\
        );

    \I__8822\ : Odrv4
    port map (
            O => \N__42545\,
            I => n2915
        );

    \I__8821\ : Odrv4
    port map (
            O => \N__42542\,
            I => n2915
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__42539\,
            I => n2915
        );

    \I__8819\ : InMux
    port map (
            O => \N__42532\,
            I => \N__42528\
        );

    \I__8818\ : InMux
    port map (
            O => \N__42531\,
            I => \N__42525\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__42528\,
            I => \N__42519\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__42525\,
            I => \N__42519\
        );

    \I__8815\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42516\
        );

    \I__8814\ : Span4Mux_v
    port map (
            O => \N__42519\,
            I => \N__42511\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__42516\,
            I => \N__42511\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__42511\,
            I => n2916
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__42508\,
            I => \n13934_cascade_\
        );

    \I__8810\ : InMux
    port map (
            O => \N__42505\,
            I => \N__42502\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__42502\,
            I => \N__42499\
        );

    \I__8808\ : Odrv4
    port map (
            O => \N__42499\,
            I => n13942
        );

    \I__8807\ : InMux
    port map (
            O => \N__42496\,
            I => \N__42493\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__42493\,
            I => \N__42490\
        );

    \I__8805\ : Span4Mux_h
    port map (
            O => \N__42490\,
            I => \N__42487\
        );

    \I__8804\ : Odrv4
    port map (
            O => \N__42487\,
            I => n2679
        );

    \I__8803\ : CascadeMux
    port map (
            O => \N__42484\,
            I => \N__42481\
        );

    \I__8802\ : InMux
    port map (
            O => \N__42481\,
            I => \N__42478\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__42478\,
            I => \N__42475\
        );

    \I__8800\ : Span4Mux_v
    port map (
            O => \N__42475\,
            I => \N__42470\
        );

    \I__8799\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42467\
        );

    \I__8798\ : InMux
    port map (
            O => \N__42473\,
            I => \N__42464\
        );

    \I__8797\ : Span4Mux_h
    port map (
            O => \N__42470\,
            I => \N__42461\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__42467\,
            I => \N__42458\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__42464\,
            I => \N__42455\
        );

    \I__8794\ : Odrv4
    port map (
            O => \N__42461\,
            I => n2612
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__42458\,
            I => n2612
        );

    \I__8792\ : Odrv4
    port map (
            O => \N__42455\,
            I => n2612
        );

    \I__8791\ : InMux
    port map (
            O => \N__42448\,
            I => \N__42445\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__42445\,
            I => \N__42439\
        );

    \I__8789\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42436\
        );

    \I__8788\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42433\
        );

    \I__8787\ : CascadeMux
    port map (
            O => \N__42442\,
            I => \N__42424\
        );

    \I__8786\ : Span4Mux_v
    port map (
            O => \N__42439\,
            I => \N__42419\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__42436\,
            I => \N__42416\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__42433\,
            I => \N__42413\
        );

    \I__8783\ : CascadeMux
    port map (
            O => \N__42432\,
            I => \N__42409\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__42431\,
            I => \N__42406\
        );

    \I__8781\ : CascadeMux
    port map (
            O => \N__42430\,
            I => \N__42399\
        );

    \I__8780\ : CascadeMux
    port map (
            O => \N__42429\,
            I => \N__42392\
        );

    \I__8779\ : CascadeMux
    port map (
            O => \N__42428\,
            I => \N__42387\
        );

    \I__8778\ : CascadeMux
    port map (
            O => \N__42427\,
            I => \N__42384\
        );

    \I__8777\ : InMux
    port map (
            O => \N__42424\,
            I => \N__42375\
        );

    \I__8776\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42375\
        );

    \I__8775\ : InMux
    port map (
            O => \N__42422\,
            I => \N__42375\
        );

    \I__8774\ : Span4Mux_v
    port map (
            O => \N__42419\,
            I => \N__42368\
        );

    \I__8773\ : Span4Mux_v
    port map (
            O => \N__42416\,
            I => \N__42368\
        );

    \I__8772\ : Span4Mux_v
    port map (
            O => \N__42413\,
            I => \N__42368\
        );

    \I__8771\ : InMux
    port map (
            O => \N__42412\,
            I => \N__42357\
        );

    \I__8770\ : InMux
    port map (
            O => \N__42409\,
            I => \N__42357\
        );

    \I__8769\ : InMux
    port map (
            O => \N__42406\,
            I => \N__42357\
        );

    \I__8768\ : InMux
    port map (
            O => \N__42405\,
            I => \N__42357\
        );

    \I__8767\ : InMux
    port map (
            O => \N__42404\,
            I => \N__42357\
        );

    \I__8766\ : InMux
    port map (
            O => \N__42403\,
            I => \N__42346\
        );

    \I__8765\ : InMux
    port map (
            O => \N__42402\,
            I => \N__42346\
        );

    \I__8764\ : InMux
    port map (
            O => \N__42399\,
            I => \N__42346\
        );

    \I__8763\ : InMux
    port map (
            O => \N__42398\,
            I => \N__42346\
        );

    \I__8762\ : InMux
    port map (
            O => \N__42397\,
            I => \N__42346\
        );

    \I__8761\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42341\
        );

    \I__8760\ : InMux
    port map (
            O => \N__42395\,
            I => \N__42341\
        );

    \I__8759\ : InMux
    port map (
            O => \N__42392\,
            I => \N__42336\
        );

    \I__8758\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42336\
        );

    \I__8757\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42325\
        );

    \I__8756\ : InMux
    port map (
            O => \N__42387\,
            I => \N__42325\
        );

    \I__8755\ : InMux
    port map (
            O => \N__42384\,
            I => \N__42325\
        );

    \I__8754\ : InMux
    port map (
            O => \N__42383\,
            I => \N__42325\
        );

    \I__8753\ : InMux
    port map (
            O => \N__42382\,
            I => \N__42325\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__42375\,
            I => n2643
        );

    \I__8751\ : Odrv4
    port map (
            O => \N__42368\,
            I => n2643
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__42357\,
            I => n2643
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__42346\,
            I => n2643
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__42341\,
            I => n2643
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__42336\,
            I => n2643
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__42325\,
            I => n2643
        );

    \I__8745\ : CascadeMux
    port map (
            O => \N__42310\,
            I => \N__42306\
        );

    \I__8744\ : CascadeMux
    port map (
            O => \N__42309\,
            I => \N__42302\
        );

    \I__8743\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42299\
        );

    \I__8742\ : InMux
    port map (
            O => \N__42305\,
            I => \N__42296\
        );

    \I__8741\ : InMux
    port map (
            O => \N__42302\,
            I => \N__42293\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__42299\,
            I => \N__42288\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__42296\,
            I => \N__42288\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__42293\,
            I => n2711
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__42288\,
            I => n2711
        );

    \I__8736\ : InMux
    port map (
            O => \N__42283\,
            I => \N__42280\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__42280\,
            I => \N__42277\
        );

    \I__8734\ : Span4Mux_v
    port map (
            O => \N__42277\,
            I => \N__42274\
        );

    \I__8733\ : Span4Mux_h
    port map (
            O => \N__42274\,
            I => \N__42270\
        );

    \I__8732\ : InMux
    port map (
            O => \N__42273\,
            I => \N__42267\
        );

    \I__8731\ : Odrv4
    port map (
            O => \N__42270\,
            I => n15467
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__42267\,
            I => n15467
        );

    \I__8729\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42258\
        );

    \I__8728\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42255\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__42258\,
            I => \N__42252\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__42255\,
            I => \N__42249\
        );

    \I__8725\ : Span4Mux_v
    port map (
            O => \N__42252\,
            I => \N__42245\
        );

    \I__8724\ : Span4Mux_v
    port map (
            O => \N__42249\,
            I => \N__42242\
        );

    \I__8723\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42239\
        );

    \I__8722\ : Odrv4
    port map (
            O => \N__42245\,
            I => n2909
        );

    \I__8721\ : Odrv4
    port map (
            O => \N__42242\,
            I => n2909
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__42239\,
            I => n2909
        );

    \I__8719\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42228\
        );

    \I__8718\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42224\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__42228\,
            I => \N__42221\
        );

    \I__8716\ : InMux
    port map (
            O => \N__42227\,
            I => \N__42218\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__42224\,
            I => \N__42215\
        );

    \I__8714\ : Span4Mux_v
    port map (
            O => \N__42221\,
            I => \N__42212\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__42218\,
            I => \N__42207\
        );

    \I__8712\ : Span4Mux_v
    port map (
            O => \N__42215\,
            I => \N__42207\
        );

    \I__8711\ : Odrv4
    port map (
            O => \N__42212\,
            I => n2713
        );

    \I__8710\ : Odrv4
    port map (
            O => \N__42207\,
            I => n2713
        );

    \I__8709\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42199\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__42199\,
            I => n2780
        );

    \I__8707\ : CascadeMux
    port map (
            O => \N__42196\,
            I => \n14322_cascade_\
        );

    \I__8706\ : CascadeMux
    port map (
            O => \N__42193\,
            I => \N__42190\
        );

    \I__8705\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42187\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__42187\,
            I => n14328
        );

    \I__8703\ : CascadeMux
    port map (
            O => \N__42184\,
            I => \N__42180\
        );

    \I__8702\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42177\
        );

    \I__8701\ : InMux
    port map (
            O => \N__42180\,
            I => \N__42174\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__42177\,
            I => \N__42168\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__42174\,
            I => \N__42168\
        );

    \I__8698\ : InMux
    port map (
            O => \N__42173\,
            I => \N__42165\
        );

    \I__8697\ : Odrv12
    port map (
            O => \N__42168\,
            I => n2724
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__42165\,
            I => n2724
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__42160\,
            I => \N__42157\
        );

    \I__8694\ : InMux
    port map (
            O => \N__42157\,
            I => \N__42154\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__42154\,
            I => \N__42151\
        );

    \I__8692\ : Odrv4
    port map (
            O => \N__42151\,
            I => n2791
        );

    \I__8691\ : InMux
    port map (
            O => \N__42148\,
            I => \N__42145\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__42145\,
            I => n2786
        );

    \I__8689\ : InMux
    port map (
            O => \N__42142\,
            I => \N__42139\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__42139\,
            I => \N__42135\
        );

    \I__8687\ : InMux
    port map (
            O => \N__42138\,
            I => \N__42132\
        );

    \I__8686\ : Span4Mux_h
    port map (
            O => \N__42135\,
            I => \N__42126\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__42132\,
            I => \N__42126\
        );

    \I__8684\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42123\
        );

    \I__8683\ : Odrv4
    port map (
            O => \N__42126\,
            I => n2719
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__42123\,
            I => n2719
        );

    \I__8681\ : InMux
    port map (
            O => \N__42118\,
            I => \N__42114\
        );

    \I__8680\ : InMux
    port map (
            O => \N__42117\,
            I => \N__42111\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__42114\,
            I => \N__42106\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__42111\,
            I => \N__42106\
        );

    \I__8677\ : Span4Mux_v
    port map (
            O => \N__42106\,
            I => \N__42103\
        );

    \I__8676\ : Odrv4
    port map (
            O => \N__42103\,
            I => n2921
        );

    \I__8675\ : CascadeMux
    port map (
            O => \N__42100\,
            I => \n2921_cascade_\
        );

    \I__8674\ : InMux
    port map (
            O => \N__42097\,
            I => \N__42094\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__42094\,
            I => n2778
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__42091\,
            I => \N__42087\
        );

    \I__8671\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42084\
        );

    \I__8670\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42081\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__42084\,
            I => \N__42078\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__42081\,
            I => \N__42075\
        );

    \I__8667\ : Span4Mux_h
    port map (
            O => \N__42078\,
            I => \N__42072\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__42075\,
            I => \N__42069\
        );

    \I__8665\ : Odrv4
    port map (
            O => \N__42072\,
            I => n2917
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__42069\,
            I => n2917
        );

    \I__8663\ : InMux
    port map (
            O => \N__42064\,
            I => \N__42060\
        );

    \I__8662\ : CascadeMux
    port map (
            O => \N__42063\,
            I => \N__42057\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__42060\,
            I => \N__42054\
        );

    \I__8660\ : InMux
    port map (
            O => \N__42057\,
            I => \N__42050\
        );

    \I__8659\ : Span4Mux_v
    port map (
            O => \N__42054\,
            I => \N__42047\
        );

    \I__8658\ : InMux
    port map (
            O => \N__42053\,
            I => \N__42044\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__42050\,
            I => n2918
        );

    \I__8656\ : Odrv4
    port map (
            O => \N__42047\,
            I => n2918
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__42044\,
            I => n2918
        );

    \I__8654\ : InMux
    port map (
            O => \N__42037\,
            I => \N__42034\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__42034\,
            I => n13926
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__42031\,
            I => \n2917_cascade_\
        );

    \I__8651\ : CascadeMux
    port map (
            O => \N__42028\,
            I => \N__42024\
        );

    \I__8650\ : InMux
    port map (
            O => \N__42027\,
            I => \N__42021\
        );

    \I__8649\ : InMux
    port map (
            O => \N__42024\,
            I => \N__42018\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__42021\,
            I => \N__42015\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__42018\,
            I => \N__42012\
        );

    \I__8646\ : Span4Mux_v
    port map (
            O => \N__42015\,
            I => \N__42009\
        );

    \I__8645\ : Span4Mux_h
    port map (
            O => \N__42012\,
            I => \N__42006\
        );

    \I__8644\ : Span4Mux_h
    port map (
            O => \N__42009\,
            I => \N__42003\
        );

    \I__8643\ : Odrv4
    port map (
            O => \N__42006\,
            I => n2709
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__42003\,
            I => n2709
        );

    \I__8641\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41995\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__41995\,
            I => n2798
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__41992\,
            I => \n2742_cascade_\
        );

    \I__8638\ : InMux
    port map (
            O => \N__41989\,
            I => \N__41986\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__41986\,
            I => \N__41982\
        );

    \I__8636\ : CascadeMux
    port map (
            O => \N__41985\,
            I => \N__41978\
        );

    \I__8635\ : Span4Mux_v
    port map (
            O => \N__41982\,
            I => \N__41975\
        );

    \I__8634\ : InMux
    port map (
            O => \N__41981\,
            I => \N__41972\
        );

    \I__8633\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41969\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__41975\,
            I => n2731
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__41972\,
            I => n2731
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__41969\,
            I => n2731
        );

    \I__8629\ : CascadeMux
    port map (
            O => \N__41962\,
            I => \N__41958\
        );

    \I__8628\ : InMux
    port map (
            O => \N__41961\,
            I => \N__41955\
        );

    \I__8627\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41952\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__41955\,
            I => \N__41946\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__41952\,
            I => \N__41946\
        );

    \I__8624\ : InMux
    port map (
            O => \N__41951\,
            I => \N__41943\
        );

    \I__8623\ : Odrv4
    port map (
            O => \N__41946\,
            I => n2728
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__41943\,
            I => n2728
        );

    \I__8621\ : CascadeMux
    port map (
            O => \N__41938\,
            I => \N__41935\
        );

    \I__8620\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41932\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__41932\,
            I => n2795
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__41929\,
            I => \n14238_cascade_\
        );

    \I__8617\ : CascadeMux
    port map (
            O => \N__41926\,
            I => \n14240_cascade_\
        );

    \I__8616\ : CascadeMux
    port map (
            O => \N__41923\,
            I => \N__41920\
        );

    \I__8615\ : InMux
    port map (
            O => \N__41920\,
            I => \N__41916\
        );

    \I__8614\ : InMux
    port map (
            O => \N__41919\,
            I => \N__41913\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41908\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__41913\,
            I => \N__41908\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__41908\,
            I => n2720
        );

    \I__8610\ : InMux
    port map (
            O => \N__41905\,
            I => \N__41902\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__41902\,
            I => \N__41899\
        );

    \I__8608\ : Odrv4
    port map (
            O => \N__41899\,
            I => n2787
        );

    \I__8607\ : InMux
    port map (
            O => \N__41896\,
            I => \N__41893\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__41893\,
            I => n2789
        );

    \I__8605\ : CascadeMux
    port map (
            O => \N__41890\,
            I => \N__41887\
        );

    \I__8604\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41883\
        );

    \I__8603\ : CascadeMux
    port map (
            O => \N__41886\,
            I => \N__41880\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41876\
        );

    \I__8601\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41873\
        );

    \I__8600\ : InMux
    port map (
            O => \N__41879\,
            I => \N__41870\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__41876\,
            I => n2722
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__41873\,
            I => n2722
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__41870\,
            I => n2722
        );

    \I__8596\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41860\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__41860\,
            I => n2797
        );

    \I__8594\ : InMux
    port map (
            O => \N__41857\,
            I => \N__41853\
        );

    \I__8593\ : CascadeMux
    port map (
            O => \N__41856\,
            I => \N__41849\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__41853\,
            I => \N__41846\
        );

    \I__8591\ : InMux
    port map (
            O => \N__41852\,
            I => \N__41843\
        );

    \I__8590\ : InMux
    port map (
            O => \N__41849\,
            I => \N__41840\
        );

    \I__8589\ : Odrv4
    port map (
            O => \N__41846\,
            I => n2730
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__41843\,
            I => n2730
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__41840\,
            I => n2730
        );

    \I__8586\ : CascadeMux
    port map (
            O => \N__41833\,
            I => \N__41829\
        );

    \I__8585\ : InMux
    port map (
            O => \N__41832\,
            I => \N__41825\
        );

    \I__8584\ : InMux
    port map (
            O => \N__41829\,
            I => \N__41820\
        );

    \I__8583\ : InMux
    port map (
            O => \N__41828\,
            I => \N__41820\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__41825\,
            I => \N__41817\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__41820\,
            I => \N__41812\
        );

    \I__8580\ : Span4Mux_h
    port map (
            O => \N__41817\,
            I => \N__41812\
        );

    \I__8579\ : Odrv4
    port map (
            O => \N__41812\,
            I => n23_adj_618
        );

    \I__8578\ : CascadeMux
    port map (
            O => \N__41809\,
            I => \n14800_cascade_\
        );

    \I__8577\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41803\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__41803\,
            I => n19_adj_616
        );

    \I__8575\ : InMux
    port map (
            O => \N__41800\,
            I => \N__41794\
        );

    \I__8574\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41794\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__41794\,
            I => \N__41791\
        );

    \I__8572\ : Span4Mux_h
    port map (
            O => \N__41791\,
            I => \N__41788\
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__41788\,
            I => n17_adj_615
        );

    \I__8570\ : CascadeMux
    port map (
            O => \N__41785\,
            I => \N__41782\
        );

    \I__8569\ : InMux
    port map (
            O => \N__41782\,
            I => \N__41779\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__41779\,
            I => \N__41775\
        );

    \I__8567\ : InMux
    port map (
            O => \N__41778\,
            I => \N__41772\
        );

    \I__8566\ : Span4Mux_s2_v
    port map (
            O => \N__41775\,
            I => \N__41767\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__41772\,
            I => \N__41767\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__41767\,
            I => n9_adj_608
        );

    \I__8563\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41758\
        );

    \I__8562\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41758\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__41758\,
            I => \N__41755\
        );

    \I__8560\ : Odrv4
    port map (
            O => \N__41755\,
            I => n21_adj_617
        );

    \I__8559\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41749\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__41749\,
            I => \N__41746\
        );

    \I__8557\ : Odrv4
    port map (
            O => \N__41746\,
            I => n14734
        );

    \I__8556\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41740\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__41740\,
            I => \N__41737\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__41737\,
            I => \N__41734\
        );

    \I__8553\ : Odrv4
    port map (
            O => \N__41734\,
            I => n14874
        );

    \I__8552\ : InMux
    port map (
            O => \N__41731\,
            I => \N__41728\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__41728\,
            I => \N__41724\
        );

    \I__8550\ : InMux
    port map (
            O => \N__41727\,
            I => \N__41721\
        );

    \I__8549\ : Span4Mux_h
    port map (
            O => \N__41724\,
            I => \N__41716\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__41721\,
            I => \N__41716\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__41716\,
            I => pwm_setpoint_12
        );

    \I__8546\ : InMux
    port map (
            O => \N__41713\,
            I => \N__41708\
        );

    \I__8545\ : InMux
    port map (
            O => \N__41712\,
            I => \N__41705\
        );

    \I__8544\ : InMux
    port map (
            O => \N__41711\,
            I => \N__41702\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__41708\,
            I => \N__41699\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__41705\,
            I => pwm_counter_12
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__41702\,
            I => pwm_counter_12
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__41699\,
            I => pwm_counter_12
        );

    \I__8539\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41686\
        );

    \I__8538\ : InMux
    port map (
            O => \N__41691\,
            I => \N__41686\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__41686\,
            I => \N__41682\
        );

    \I__8536\ : InMux
    port map (
            O => \N__41685\,
            I => \N__41679\
        );

    \I__8535\ : Odrv4
    port map (
            O => \N__41682\,
            I => n25_adj_620
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__41679\,
            I => n25_adj_620
        );

    \I__8533\ : InMux
    port map (
            O => \N__41674\,
            I => \N__41670\
        );

    \I__8532\ : CascadeMux
    port map (
            O => \N__41673\,
            I => \N__41667\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__41670\,
            I => \N__41663\
        );

    \I__8530\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41660\
        );

    \I__8529\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41657\
        );

    \I__8528\ : Odrv4
    port map (
            O => \N__41663\,
            I => n2723
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__41660\,
            I => n2723
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__41657\,
            I => n2723
        );

    \I__8525\ : CascadeMux
    port map (
            O => \N__41650\,
            I => \N__41647\
        );

    \I__8524\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41644\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__41644\,
            I => n2790
        );

    \I__8522\ : CascadeMux
    port map (
            O => \N__41641\,
            I => \N__41638\
        );

    \I__8521\ : InMux
    port map (
            O => \N__41638\,
            I => \N__41634\
        );

    \I__8520\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41631\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__41634\,
            I => \N__41628\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__41631\,
            I => \N__41625\
        );

    \I__8517\ : Span4Mux_h
    port map (
            O => \N__41628\,
            I => \N__41622\
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__41625\,
            I => n2725
        );

    \I__8515\ : Odrv4
    port map (
            O => \N__41622\,
            I => n2725
        );

    \I__8514\ : InMux
    port map (
            O => \N__41617\,
            I => \N__41614\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__41614\,
            I => n2792
        );

    \I__8512\ : InMux
    port map (
            O => \N__41611\,
            I => \N__41608\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__41608\,
            I => \N__41605\
        );

    \I__8510\ : Odrv4
    port map (
            O => \N__41605\,
            I => n13403
        );

    \I__8509\ : InMux
    port map (
            O => \N__41602\,
            I => \N__41599\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__41599\,
            I => \N__41596\
        );

    \I__8507\ : Odrv4
    port map (
            O => \N__41596\,
            I => n14048
        );

    \I__8506\ : InMux
    port map (
            O => \N__41593\,
            I => \N__41590\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__41590\,
            I => \N__41586\
        );

    \I__8504\ : InMux
    port map (
            O => \N__41589\,
            I => \N__41583\
        );

    \I__8503\ : Span4Mux_h
    port map (
            O => \N__41586\,
            I => \N__41580\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__41583\,
            I => n2714
        );

    \I__8501\ : Odrv4
    port map (
            O => \N__41580\,
            I => n2714
        );

    \I__8500\ : CascadeMux
    port map (
            O => \N__41575\,
            I => \n14054_cascade_\
        );

    \I__8499\ : CascadeMux
    port map (
            O => \N__41572\,
            I => \N__41569\
        );

    \I__8498\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41564\
        );

    \I__8497\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41561\
        );

    \I__8496\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41558\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__41564\,
            I => \N__41555\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__41561\,
            I => \N__41552\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__41558\,
            I => \N__41549\
        );

    \I__8492\ : Span4Mux_v
    port map (
            O => \N__41555\,
            I => \N__41544\
        );

    \I__8491\ : Span4Mux_v
    port map (
            O => \N__41552\,
            I => \N__41544\
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__41549\,
            I => n2710
        );

    \I__8489\ : Odrv4
    port map (
            O => \N__41544\,
            I => n2710
        );

    \I__8488\ : CascadeMux
    port map (
            O => \N__41539\,
            I => \n14060_cascade_\
        );

    \I__8487\ : CascadeMux
    port map (
            O => \N__41536\,
            I => \PWM.n13596_cascade_\
        );

    \I__8486\ : InMux
    port map (
            O => \N__41533\,
            I => \N__41527\
        );

    \I__8485\ : InMux
    port map (
            O => \N__41532\,
            I => \N__41524\
        );

    \I__8484\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41519\
        );

    \I__8483\ : InMux
    port map (
            O => \N__41530\,
            I => \N__41519\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__41527\,
            I => pwm_counter_8
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__41524\,
            I => pwm_counter_8
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__41519\,
            I => pwm_counter_8
        );

    \I__8479\ : InMux
    port map (
            O => \N__41512\,
            I => \N__41509\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__41509\,
            I => \N__41506\
        );

    \I__8477\ : Span4Mux_h
    port map (
            O => \N__41506\,
            I => \N__41503\
        );

    \I__8476\ : Odrv4
    port map (
            O => \N__41503\,
            I => \PWM.n26\
        );

    \I__8475\ : InMux
    port map (
            O => \N__41500\,
            I => \N__41497\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__41497\,
            I => \N__41493\
        );

    \I__8473\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41490\
        );

    \I__8472\ : Span4Mux_h
    port map (
            O => \N__41493\,
            I => \N__41487\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__41490\,
            I => \N__41484\
        );

    \I__8470\ : Odrv4
    port map (
            O => \N__41487\,
            I => n4823
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__41484\,
            I => n4823
        );

    \I__8468\ : CascadeMux
    port map (
            O => \N__41479\,
            I => \PWM.n17_cascade_\
        );

    \I__8467\ : InMux
    port map (
            O => \N__41476\,
            I => \N__41471\
        );

    \I__8466\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41468\
        );

    \I__8465\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41465\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__41471\,
            I => \N__41462\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__41468\,
            I => pwm_counter_31
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__41465\,
            I => pwm_counter_31
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__41462\,
            I => pwm_counter_31
        );

    \I__8460\ : CascadeMux
    port map (
            O => \N__41455\,
            I => \PWM.n29_cascade_\
        );

    \I__8459\ : InMux
    port map (
            O => \N__41452\,
            I => \N__41449\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__41449\,
            I => \N__41446\
        );

    \I__8457\ : Span4Mux_s2_v
    port map (
            O => \N__41446\,
            I => \N__41443\
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__41443\,
            I => \PWM.n27\
        );

    \I__8455\ : SRMux
    port map (
            O => \N__41440\,
            I => \N__41437\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__41437\,
            I => \N__41433\
        );

    \I__8453\ : SRMux
    port map (
            O => \N__41436\,
            I => \N__41430\
        );

    \I__8452\ : Span4Mux_v
    port map (
            O => \N__41433\,
            I => \N__41424\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__41430\,
            I => \N__41424\
        );

    \I__8450\ : SRMux
    port map (
            O => \N__41429\,
            I => \N__41420\
        );

    \I__8449\ : Span4Mux_s1_v
    port map (
            O => \N__41424\,
            I => \N__41417\
        );

    \I__8448\ : SRMux
    port map (
            O => \N__41423\,
            I => \N__41414\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__41420\,
            I => \N__41407\
        );

    \I__8446\ : Span4Mux_h
    port map (
            O => \N__41417\,
            I => \N__41407\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__41414\,
            I => \N__41407\
        );

    \I__8444\ : Span4Mux_v
    port map (
            O => \N__41407\,
            I => \N__41404\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__41404\,
            I => \PWM.pwm_counter_31__N_401\
        );

    \I__8442\ : InMux
    port map (
            O => \N__41401\,
            I => \N__41396\
        );

    \I__8441\ : InMux
    port map (
            O => \N__41400\,
            I => \N__41391\
        );

    \I__8440\ : InMux
    port map (
            O => \N__41399\,
            I => \N__41391\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__41396\,
            I => pwm_counter_19
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__41391\,
            I => pwm_counter_19
        );

    \I__8437\ : InMux
    port map (
            O => \N__41386\,
            I => \N__41383\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__41383\,
            I => \N__41380\
        );

    \I__8435\ : Span4Mux_h
    port map (
            O => \N__41380\,
            I => \N__41377\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__41377\,
            I => n39
        );

    \I__8433\ : InMux
    port map (
            O => \N__41374\,
            I => \N__41368\
        );

    \I__8432\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41368\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__41368\,
            I => pwm_setpoint_19
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__41365\,
            I => \n39_cascade_\
        );

    \I__8429\ : InMux
    port map (
            O => \N__41362\,
            I => \N__41359\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__41359\,
            I => \N__41356\
        );

    \I__8427\ : Span4Mux_h
    port map (
            O => \N__41356\,
            I => \N__41353\
        );

    \I__8426\ : Odrv4
    port map (
            O => \N__41353\,
            I => n14883
        );

    \I__8425\ : CascadeMux
    port map (
            O => \N__41350\,
            I => \N__41347\
        );

    \I__8424\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41344\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__41344\,
            I => \N__41338\
        );

    \I__8422\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41335\
        );

    \I__8421\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41332\
        );

    \I__8420\ : InMux
    port map (
            O => \N__41341\,
            I => \N__41329\
        );

    \I__8419\ : Span4Mux_h
    port map (
            O => \N__41338\,
            I => \N__41324\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__41335\,
            I => \N__41324\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__41332\,
            I => pwm_counter_9
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__41329\,
            I => pwm_counter_9
        );

    \I__8415\ : Odrv4
    port map (
            O => \N__41324\,
            I => pwm_counter_9
        );

    \I__8414\ : InMux
    port map (
            O => \N__41317\,
            I => \N__41314\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__41314\,
            I => \N__41311\
        );

    \I__8412\ : Odrv4
    port map (
            O => \N__41311\,
            I => n14804
        );

    \I__8411\ : CascadeMux
    port map (
            O => \N__41308\,
            I => \n19_adj_616_cascade_\
        );

    \I__8410\ : InMux
    port map (
            O => \N__41305\,
            I => \N__41301\
        );

    \I__8409\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41298\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__41301\,
            I => n15_adj_613
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__41298\,
            I => n15_adj_613
        );

    \I__8406\ : InMux
    port map (
            O => \N__41293\,
            I => \N__41287\
        );

    \I__8405\ : InMux
    port map (
            O => \N__41292\,
            I => \N__41287\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__41287\,
            I => pwm_setpoint_10
        );

    \I__8403\ : CascadeMux
    port map (
            O => \N__41284\,
            I => \n11_adj_610_cascade_\
        );

    \I__8402\ : InMux
    port map (
            O => \N__41281\,
            I => \N__41275\
        );

    \I__8401\ : InMux
    port map (
            O => \N__41280\,
            I => \N__41275\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__41275\,
            I => pwm_setpoint_5
        );

    \I__8399\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41268\
        );

    \I__8398\ : InMux
    port map (
            O => \N__41271\,
            I => \N__41265\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__41268\,
            I => \N__41262\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__41265\,
            I => \N__41259\
        );

    \I__8395\ : Span4Mux_h
    port map (
            O => \N__41262\,
            I => \N__41256\
        );

    \I__8394\ : Odrv4
    port map (
            O => \N__41259\,
            I => pwm_setpoint_6
        );

    \I__8393\ : Odrv4
    port map (
            O => \N__41256\,
            I => pwm_setpoint_6
        );

    \I__8392\ : SRMux
    port map (
            O => \N__41251\,
            I => \N__41248\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__41248\,
            I => \N__41245\
        );

    \I__8390\ : Span4Mux_h
    port map (
            O => \N__41245\,
            I => \N__41242\
        );

    \I__8389\ : Span4Mux_s2_v
    port map (
            O => \N__41242\,
            I => \N__41239\
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__41239\,
            I => n4825
        );

    \I__8387\ : InMux
    port map (
            O => \N__41236\,
            I => \N__41230\
        );

    \I__8386\ : InMux
    port map (
            O => \N__41235\,
            I => \N__41230\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__41230\,
            I => \N__41227\
        );

    \I__8384\ : Span4Mux_s3_v
    port map (
            O => \N__41227\,
            I => \N__41224\
        );

    \I__8383\ : Odrv4
    port map (
            O => \N__41224\,
            I => n13_adj_612
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__41221\,
            I => \N__41218\
        );

    \I__8381\ : InMux
    port map (
            O => \N__41218\,
            I => \N__41215\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__41215\,
            I => n11_adj_610
        );

    \I__8379\ : InMux
    port map (
            O => \N__41212\,
            I => \N__41209\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__41209\,
            I => \N__41206\
        );

    \I__8377\ : Odrv4
    port map (
            O => \N__41206\,
            I => n14745
        );

    \I__8376\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41197\
        );

    \I__8375\ : InMux
    port map (
            O => \N__41202\,
            I => \N__41197\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__41197\,
            I => \N__41194\
        );

    \I__8373\ : Odrv4
    port map (
            O => \N__41194\,
            I => pwm_setpoint_20
        );

    \I__8372\ : InMux
    port map (
            O => \N__41191\,
            I => \N__41187\
        );

    \I__8371\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41183\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__41187\,
            I => \N__41180\
        );

    \I__8369\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41177\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__41183\,
            I => pwm_counter_5
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__41180\,
            I => pwm_counter_5
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__41177\,
            I => pwm_counter_5
        );

    \I__8365\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41166\
        );

    \I__8364\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41161\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__41166\,
            I => \N__41158\
        );

    \I__8362\ : InMux
    port map (
            O => \N__41165\,
            I => \N__41155\
        );

    \I__8361\ : InMux
    port map (
            O => \N__41164\,
            I => \N__41152\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__41161\,
            I => pwm_counter_6
        );

    \I__8359\ : Odrv4
    port map (
            O => \N__41158\,
            I => pwm_counter_6
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__41155\,
            I => pwm_counter_6
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__41152\,
            I => pwm_counter_6
        );

    \I__8356\ : CascadeMux
    port map (
            O => \N__41143\,
            I => \N__41136\
        );

    \I__8355\ : CascadeMux
    port map (
            O => \N__41142\,
            I => \N__41133\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__41141\,
            I => \N__41128\
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__41140\,
            I => \N__41125\
        );

    \I__8352\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41121\
        );

    \I__8351\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41116\
        );

    \I__8350\ : InMux
    port map (
            O => \N__41133\,
            I => \N__41116\
        );

    \I__8349\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41107\
        );

    \I__8348\ : InMux
    port map (
            O => \N__41131\,
            I => \N__41107\
        );

    \I__8347\ : InMux
    port map (
            O => \N__41128\,
            I => \N__41107\
        );

    \I__8346\ : InMux
    port map (
            O => \N__41125\,
            I => \N__41107\
        );

    \I__8345\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41104\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__41121\,
            I => n4_adj_698
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__41116\,
            I => n4_adj_698
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__41107\,
            I => n4_adj_698
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__41104\,
            I => n4_adj_698
        );

    \I__8340\ : CascadeMux
    port map (
            O => \N__41095\,
            I => \N__41091\
        );

    \I__8339\ : CascadeMux
    port map (
            O => \N__41094\,
            I => \N__41088\
        );

    \I__8338\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41085\
        );

    \I__8337\ : InMux
    port map (
            O => \N__41088\,
            I => \N__41081\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__41085\,
            I => \N__41078\
        );

    \I__8335\ : InMux
    port map (
            O => \N__41084\,
            I => \N__41075\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__41081\,
            I => dti_counter_5
        );

    \I__8333\ : Odrv4
    port map (
            O => \N__41078\,
            I => dti_counter_5
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__41075\,
            I => dti_counter_5
        );

    \I__8331\ : InMux
    port map (
            O => \N__41068\,
            I => \N__41061\
        );

    \I__8330\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41061\
        );

    \I__8329\ : InMux
    port map (
            O => \N__41066\,
            I => \N__41052\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__41061\,
            I => \N__41049\
        );

    \I__8327\ : InMux
    port map (
            O => \N__41060\,
            I => \N__41046\
        );

    \I__8326\ : InMux
    port map (
            O => \N__41059\,
            I => \N__41035\
        );

    \I__8325\ : InMux
    port map (
            O => \N__41058\,
            I => \N__41035\
        );

    \I__8324\ : InMux
    port map (
            O => \N__41057\,
            I => \N__41035\
        );

    \I__8323\ : InMux
    port map (
            O => \N__41056\,
            I => \N__41035\
        );

    \I__8322\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41035\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__41052\,
            I => commutation_state_prev_0
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__41049\,
            I => commutation_state_prev_0
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__41046\,
            I => commutation_state_prev_0
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__41035\,
            I => commutation_state_prev_0
        );

    \I__8317\ : InMux
    port map (
            O => \N__41026\,
            I => \N__41023\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__41023\,
            I => n14689
        );

    \I__8315\ : InMux
    port map (
            O => \N__41020\,
            I => \N__41014\
        );

    \I__8314\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41014\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__41014\,
            I => pwm_setpoint_2
        );

    \I__8312\ : InMux
    port map (
            O => \N__41011\,
            I => \N__41008\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__41008\,
            I => \N__41004\
        );

    \I__8310\ : InMux
    port map (
            O => \N__41007\,
            I => \N__41001\
        );

    \I__8309\ : Span4Mux_s3_v
    port map (
            O => \N__41004\,
            I => \N__40996\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__41001\,
            I => \N__40996\
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__40996\,
            I => pwm_setpoint_11
        );

    \I__8306\ : InMux
    port map (
            O => \N__40993\,
            I => \N__40989\
        );

    \I__8305\ : InMux
    port map (
            O => \N__40992\,
            I => \N__40986\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__40989\,
            I => \N__40981\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__40986\,
            I => \N__40981\
        );

    \I__8302\ : Span4Mux_s3_v
    port map (
            O => \N__40981\,
            I => \N__40978\
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__40978\,
            I => pwm_setpoint_8
        );

    \I__8300\ : InMux
    port map (
            O => \N__40975\,
            I => \N__40970\
        );

    \I__8299\ : InMux
    port map (
            O => \N__40974\,
            I => \N__40967\
        );

    \I__8298\ : InMux
    port map (
            O => \N__40973\,
            I => \N__40964\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__40970\,
            I => pwm_counter_10
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__40967\,
            I => pwm_counter_10
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__40964\,
            I => pwm_counter_10
        );

    \I__8294\ : CascadeMux
    port map (
            O => \N__40957\,
            I => \n21_adj_617_cascade_\
        );

    \I__8293\ : InMux
    port map (
            O => \N__40954\,
            I => \N__40951\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__40951\,
            I => n6_adj_606
        );

    \I__8291\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40945\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__40945\,
            I => \N__40942\
        );

    \I__8289\ : Span4Mux_h
    port map (
            O => \N__40942\,
            I => \N__40939\
        );

    \I__8288\ : Odrv4
    port map (
            O => \N__40939\,
            I => n14842
        );

    \I__8287\ : InMux
    port map (
            O => \N__40936\,
            I => \N__40933\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__40933\,
            I => \N__40930\
        );

    \I__8285\ : Odrv4
    port map (
            O => \N__40930\,
            I => n14690
        );

    \I__8284\ : CascadeMux
    port map (
            O => \N__40927\,
            I => \N__40922\
        );

    \I__8283\ : InMux
    port map (
            O => \N__40926\,
            I => \N__40919\
        );

    \I__8282\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40916\
        );

    \I__8281\ : InMux
    port map (
            O => \N__40922\,
            I => \N__40913\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__40919\,
            I => dti_counter_4
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__40916\,
            I => dti_counter_4
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__40913\,
            I => dti_counter_4
        );

    \I__8277\ : InMux
    port map (
            O => \N__40906\,
            I => n12745
        );

    \I__8276\ : InMux
    port map (
            O => \N__40903\,
            I => n12746
        );

    \I__8275\ : InMux
    port map (
            O => \N__40900\,
            I => \N__40897\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__40897\,
            I => n14688
        );

    \I__8273\ : InMux
    port map (
            O => \N__40894\,
            I => \N__40889\
        );

    \I__8272\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40884\
        );

    \I__8271\ : InMux
    port map (
            O => \N__40892\,
            I => \N__40884\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__40889\,
            I => dti_counter_6
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__40884\,
            I => dti_counter_6
        );

    \I__8268\ : InMux
    port map (
            O => \N__40879\,
            I => n12747
        );

    \I__8267\ : InMux
    port map (
            O => \N__40876\,
            I => \N__40873\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__40873\,
            I => n14687
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__40870\,
            I => \N__40864\
        );

    \I__8264\ : CascadeMux
    port map (
            O => \N__40869\,
            I => \N__40860\
        );

    \I__8263\ : CascadeMux
    port map (
            O => \N__40868\,
            I => \N__40856\
        );

    \I__8262\ : InMux
    port map (
            O => \N__40867\,
            I => \N__40840\
        );

    \I__8261\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40840\
        );

    \I__8260\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40840\
        );

    \I__8259\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40840\
        );

    \I__8258\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40840\
        );

    \I__8257\ : InMux
    port map (
            O => \N__40856\,
            I => \N__40840\
        );

    \I__8256\ : InMux
    port map (
            O => \N__40855\,
            I => \N__40840\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__40840\,
            I => \N__40837\
        );

    \I__8254\ : Odrv4
    port map (
            O => \N__40837\,
            I => n11202
        );

    \I__8253\ : InMux
    port map (
            O => \N__40834\,
            I => n12748
        );

    \I__8252\ : CascadeMux
    port map (
            O => \N__40831\,
            I => \N__40827\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__40830\,
            I => \N__40824\
        );

    \I__8250\ : InMux
    port map (
            O => \N__40827\,
            I => \N__40821\
        );

    \I__8249\ : InMux
    port map (
            O => \N__40824\,
            I => \N__40817\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__40821\,
            I => \N__40814\
        );

    \I__8247\ : InMux
    port map (
            O => \N__40820\,
            I => \N__40811\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__40817\,
            I => dti_counter_7
        );

    \I__8245\ : Odrv4
    port map (
            O => \N__40814\,
            I => dti_counter_7
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__40811\,
            I => dti_counter_7
        );

    \I__8243\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40801\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__40801\,
            I => \N__40798\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__40798\,
            I => \N__40794\
        );

    \I__8240\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40791\
        );

    \I__8239\ : Odrv4
    port map (
            O => \N__40794\,
            I => pwm_setpoint_4
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__40791\,
            I => pwm_setpoint_4
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__40786\,
            I => \N__40783\
        );

    \I__8236\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40779\
        );

    \I__8235\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40776\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__40779\,
            I => \N__40773\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__40776\,
            I => pwm_counter_2
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__40773\,
            I => pwm_counter_2
        );

    \I__8231\ : InMux
    port map (
            O => \N__40768\,
            I => \N__40763\
        );

    \I__8230\ : InMux
    port map (
            O => \N__40767\,
            I => \N__40758\
        );

    \I__8229\ : InMux
    port map (
            O => \N__40766\,
            I => \N__40758\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__40763\,
            I => pwm_counter_3
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__40758\,
            I => pwm_counter_3
        );

    \I__8226\ : CascadeMux
    port map (
            O => \N__40753\,
            I => \N__40750\
        );

    \I__8225\ : InMux
    port map (
            O => \N__40750\,
            I => \N__40744\
        );

    \I__8224\ : InMux
    port map (
            O => \N__40749\,
            I => \N__40744\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__40744\,
            I => pwm_setpoint_3
        );

    \I__8222\ : CascadeMux
    port map (
            O => \N__40741\,
            I => \n14_adj_679_cascade_\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__40738\,
            I => \n4781_cascade_\
        );

    \I__8220\ : InMux
    port map (
            O => \N__40735\,
            I => \N__40732\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__40732\,
            I => n14700
        );

    \I__8218\ : InMux
    port map (
            O => \N__40729\,
            I => \N__40726\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__40726\,
            I => n1259
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__40723\,
            I => \N__40719\
        );

    \I__8215\ : InMux
    port map (
            O => \N__40722\,
            I => \N__40715\
        );

    \I__8214\ : InMux
    port map (
            O => \N__40719\,
            I => \N__40712\
        );

    \I__8213\ : InMux
    port map (
            O => \N__40718\,
            I => \N__40709\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__40715\,
            I => dti_counter_0
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__40712\,
            I => dti_counter_0
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__40709\,
            I => dti_counter_0
        );

    \I__8209\ : InMux
    port map (
            O => \N__40702\,
            I => \bfn_12_27_0_\
        );

    \I__8208\ : InMux
    port map (
            O => \N__40699\,
            I => \N__40696\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__40696\,
            I => n14693
        );

    \I__8206\ : InMux
    port map (
            O => \N__40693\,
            I => n12742
        );

    \I__8205\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40687\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__40687\,
            I => n14692
        );

    \I__8203\ : InMux
    port map (
            O => \N__40684\,
            I => n12743
        );

    \I__8202\ : InMux
    port map (
            O => \N__40681\,
            I => \N__40678\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__40678\,
            I => n14691
        );

    \I__8200\ : CascadeMux
    port map (
            O => \N__40675\,
            I => \N__40671\
        );

    \I__8199\ : CascadeMux
    port map (
            O => \N__40674\,
            I => \N__40668\
        );

    \I__8198\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40665\
        );

    \I__8197\ : InMux
    port map (
            O => \N__40668\,
            I => \N__40661\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__40665\,
            I => \N__40658\
        );

    \I__8195\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40655\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__40661\,
            I => dti_counter_3
        );

    \I__8193\ : Odrv12
    port map (
            O => \N__40658\,
            I => dti_counter_3
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__40655\,
            I => dti_counter_3
        );

    \I__8191\ : InMux
    port map (
            O => \N__40648\,
            I => n12744
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__40645\,
            I => \n13848_cascade_\
        );

    \I__8189\ : InMux
    port map (
            O => \N__40642\,
            I => \N__40639\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__40639\,
            I => \N__40636\
        );

    \I__8187\ : Odrv4
    port map (
            O => \N__40636\,
            I => n5_adj_713
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__40633\,
            I => \n13850_cascade_\
        );

    \I__8185\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40627\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__40627\,
            I => \N__40624\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__40624\,
            I => n11656
        );

    \I__8182\ : CascadeMux
    port map (
            O => \N__40621\,
            I => \n13852_cascade_\
        );

    \I__8181\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40615\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__40615\,
            I => n13854
        );

    \I__8179\ : InMux
    port map (
            O => \N__40612\,
            I => \N__40609\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__40609\,
            I => n37_adj_710
        );

    \I__8177\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40603\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__40603\,
            I => n7_adj_703
        );

    \I__8175\ : CascadeMux
    port map (
            O => \N__40600\,
            I => \n23_adj_707_cascade_\
        );

    \I__8174\ : CascadeMux
    port map (
            O => \N__40597\,
            I => \n25_adj_708_cascade_\
        );

    \I__8173\ : CascadeMux
    port map (
            O => \N__40594\,
            I => \n13832_cascade_\
        );

    \I__8172\ : InMux
    port map (
            O => \N__40591\,
            I => \N__40588\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__40588\,
            I => n13828
        );

    \I__8170\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40582\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__40582\,
            I => n13826
        );

    \I__8168\ : CascadeMux
    port map (
            O => \N__40579\,
            I => \n13840_cascade_\
        );

    \I__8167\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__40573\,
            I => n13846
        );

    \I__8165\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40567\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__40567\,
            I => \N__40564\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__40564\,
            I => n13466
        );

    \I__8162\ : InMux
    port map (
            O => \N__40561\,
            I => \N__40558\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__40558\,
            I => n14334
        );

    \I__8160\ : CascadeMux
    port map (
            O => \N__40555\,
            I => \n3121_cascade_\
        );

    \I__8159\ : CascadeMux
    port map (
            O => \N__40552\,
            I => \n3112_cascade_\
        );

    \I__8158\ : CascadeMux
    port map (
            O => \N__40549\,
            I => \N__40546\
        );

    \I__8157\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40542\
        );

    \I__8156\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40539\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__40542\,
            I => \N__40534\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__40539\,
            I => \N__40534\
        );

    \I__8153\ : Span4Mux_h
    port map (
            O => \N__40534\,
            I => \N__40530\
        );

    \I__8152\ : InMux
    port map (
            O => \N__40533\,
            I => \N__40527\
        );

    \I__8151\ : Odrv4
    port map (
            O => \N__40530\,
            I => n2911
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__40527\,
            I => n2911
        );

    \I__8149\ : CascadeMux
    port map (
            O => \N__40522\,
            I => \N__40519\
        );

    \I__8148\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40515\
        );

    \I__8147\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40512\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__40515\,
            I => n2912
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__40512\,
            I => n2912
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__40507\,
            I => \n13948_cascade_\
        );

    \I__8143\ : CascadeMux
    port map (
            O => \N__40504\,
            I => \n13954_cascade_\
        );

    \I__8142\ : InMux
    port map (
            O => \N__40501\,
            I => \N__40498\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__40498\,
            I => \N__40495\
        );

    \I__8140\ : Odrv4
    port map (
            O => \N__40495\,
            I => n2999
        );

    \I__8139\ : CascadeMux
    port map (
            O => \N__40492\,
            I => \n2940_cascade_\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__40489\,
            I => \N__40486\
        );

    \I__8137\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40483\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__40483\,
            I => \N__40480\
        );

    \I__8135\ : Odrv4
    port map (
            O => \N__40480\,
            I => n2996
        );

    \I__8134\ : CascadeMux
    port map (
            O => \N__40477\,
            I => \n14340_cascade_\
        );

    \I__8133\ : InMux
    port map (
            O => \N__40474\,
            I => \N__40471\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__40471\,
            I => \N__40467\
        );

    \I__8131\ : InMux
    port map (
            O => \N__40470\,
            I => \N__40463\
        );

    \I__8130\ : Span4Mux_v
    port map (
            O => \N__40467\,
            I => \N__40460\
        );

    \I__8129\ : InMux
    port map (
            O => \N__40466\,
            I => \N__40457\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__40463\,
            I => n2908
        );

    \I__8127\ : Odrv4
    port map (
            O => \N__40460\,
            I => n2908
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__40457\,
            I => n2908
        );

    \I__8125\ : InMux
    port map (
            O => \N__40450\,
            I => \N__40447\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__40447\,
            I => n14344
        );

    \I__8123\ : CascadeMux
    port map (
            O => \N__40444\,
            I => \n3039_cascade_\
        );

    \I__8122\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40438\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40435\
        );

    \I__8120\ : Span4Mux_h
    port map (
            O => \N__40435\,
            I => \N__40432\
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__40432\,
            I => n2777
        );

    \I__8118\ : InMux
    port map (
            O => \N__40429\,
            I => \bfn_12_20_0_\
        );

    \I__8117\ : InMux
    port map (
            O => \N__40426\,
            I => n12410
        );

    \I__8116\ : InMux
    port map (
            O => \N__40423\,
            I => \N__40420\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__40420\,
            I => \N__40417\
        );

    \I__8114\ : Span4Mux_h
    port map (
            O => \N__40417\,
            I => \N__40414\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__40414\,
            I => n2985
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__40411\,
            I => \n3017_cascade_\
        );

    \I__8111\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40405\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__40405\,
            I => \N__40402\
        );

    \I__8109\ : Span4Mux_v
    port map (
            O => \N__40402\,
            I => \N__40399\
        );

    \I__8108\ : Odrv4
    port map (
            O => \N__40399\,
            I => n2977
        );

    \I__8107\ : CascadeMux
    port map (
            O => \N__40396\,
            I => \N__40393\
        );

    \I__8106\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40390\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__40390\,
            I => \N__40387\
        );

    \I__8104\ : Span4Mux_v
    port map (
            O => \N__40387\,
            I => \N__40384\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__40384\,
            I => n2993
        );

    \I__8102\ : InMux
    port map (
            O => \N__40381\,
            I => n12400
        );

    \I__8101\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40374\
        );

    \I__8100\ : InMux
    port map (
            O => \N__40377\,
            I => \N__40371\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__40374\,
            I => \N__40366\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__40371\,
            I => \N__40366\
        );

    \I__8097\ : Span4Mux_h
    port map (
            O => \N__40366\,
            I => \N__40362\
        );

    \I__8096\ : InMux
    port map (
            O => \N__40365\,
            I => \N__40359\
        );

    \I__8095\ : Odrv4
    port map (
            O => \N__40362\,
            I => n2718
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__40359\,
            I => n2718
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__40354\,
            I => \N__40351\
        );

    \I__8092\ : InMux
    port map (
            O => \N__40351\,
            I => \N__40348\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__40348\,
            I => n2785
        );

    \I__8090\ : InMux
    port map (
            O => \N__40345\,
            I => \bfn_12_19_0_\
        );

    \I__8089\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40337\
        );

    \I__8088\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40334\
        );

    \I__8087\ : InMux
    port map (
            O => \N__40340\,
            I => \N__40331\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40328\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__40334\,
            I => \N__40325\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__40331\,
            I => n2717
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__40328\,
            I => n2717
        );

    \I__8082\ : Odrv4
    port map (
            O => \N__40325\,
            I => n2717
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__40318\,
            I => \N__40315\
        );

    \I__8080\ : InMux
    port map (
            O => \N__40315\,
            I => \N__40312\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__40312\,
            I => n2784
        );

    \I__8078\ : InMux
    port map (
            O => \N__40309\,
            I => n12402
        );

    \I__8077\ : InMux
    port map (
            O => \N__40306\,
            I => n12403
        );

    \I__8076\ : InMux
    port map (
            O => \N__40303\,
            I => n12404
        );

    \I__8075\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40297\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__40297\,
            I => n2781
        );

    \I__8073\ : InMux
    port map (
            O => \N__40294\,
            I => n12405
        );

    \I__8072\ : InMux
    port map (
            O => \N__40291\,
            I => n12406
        );

    \I__8071\ : InMux
    port map (
            O => \N__40288\,
            I => n12407
        );

    \I__8070\ : InMux
    port map (
            O => \N__40285\,
            I => n12408
        );

    \I__8069\ : InMux
    port map (
            O => \N__40282\,
            I => n12391
        );

    \I__8068\ : InMux
    port map (
            O => \N__40279\,
            I => n12392
        );

    \I__8067\ : InMux
    port map (
            O => \N__40276\,
            I => \bfn_12_18_0_\
        );

    \I__8066\ : InMux
    port map (
            O => \N__40273\,
            I => n12394
        );

    \I__8065\ : InMux
    port map (
            O => \N__40270\,
            I => n12395
        );

    \I__8064\ : InMux
    port map (
            O => \N__40267\,
            I => n12396
        );

    \I__8063\ : InMux
    port map (
            O => \N__40264\,
            I => n12397
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__40261\,
            I => \N__40258\
        );

    \I__8061\ : InMux
    port map (
            O => \N__40258\,
            I => \N__40255\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__40255\,
            I => \N__40251\
        );

    \I__8059\ : InMux
    port map (
            O => \N__40254\,
            I => \N__40248\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__40251\,
            I => n2721
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__40248\,
            I => n2721
        );

    \I__8056\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40240\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__40240\,
            I => \N__40237\
        );

    \I__8054\ : Odrv4
    port map (
            O => \N__40237\,
            I => n2788
        );

    \I__8053\ : InMux
    port map (
            O => \N__40234\,
            I => n12398
        );

    \I__8052\ : InMux
    port map (
            O => \N__40231\,
            I => n12399
        );

    \I__8051\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40224\
        );

    \I__8050\ : InMux
    port map (
            O => \N__40227\,
            I => \N__40221\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__40224\,
            I => pwm_counter_29
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__40221\,
            I => pwm_counter_29
        );

    \I__8047\ : InMux
    port map (
            O => \N__40216\,
            I => \PWM.n12714\
        );

    \I__8046\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40209\
        );

    \I__8045\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40206\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__40209\,
            I => pwm_counter_30
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__40206\,
            I => pwm_counter_30
        );

    \I__8042\ : InMux
    port map (
            O => \N__40201\,
            I => \PWM.n12715\
        );

    \I__8041\ : InMux
    port map (
            O => \N__40198\,
            I => \PWM.n12716\
        );

    \I__8040\ : InMux
    port map (
            O => \N__40195\,
            I => \bfn_12_17_0_\
        );

    \I__8039\ : InMux
    port map (
            O => \N__40192\,
            I => n12386
        );

    \I__8038\ : InMux
    port map (
            O => \N__40189\,
            I => n12387
        );

    \I__8037\ : InMux
    port map (
            O => \N__40186\,
            I => n12388
        );

    \I__8036\ : InMux
    port map (
            O => \N__40183\,
            I => n12389
        );

    \I__8035\ : InMux
    port map (
            O => \N__40180\,
            I => n12390
        );

    \I__8034\ : InMux
    port map (
            O => \N__40177\,
            I => \N__40170\
        );

    \I__8033\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40170\
        );

    \I__8032\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40165\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__40170\,
            I => \N__40162\
        );

    \I__8030\ : InMux
    port map (
            O => \N__40169\,
            I => \N__40159\
        );

    \I__8029\ : InMux
    port map (
            O => \N__40168\,
            I => \N__40156\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__40165\,
            I => \N__40153\
        );

    \I__8027\ : Span4Mux_h
    port map (
            O => \N__40162\,
            I => \N__40150\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__40159\,
            I => pwm_counter_21
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__40156\,
            I => pwm_counter_21
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__40153\,
            I => pwm_counter_21
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__40150\,
            I => pwm_counter_21
        );

    \I__8022\ : InMux
    port map (
            O => \N__40141\,
            I => \PWM.n12706\
        );

    \I__8021\ : InMux
    port map (
            O => \N__40138\,
            I => \N__40135\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__40135\,
            I => \N__40131\
        );

    \I__8019\ : InMux
    port map (
            O => \N__40134\,
            I => \N__40127\
        );

    \I__8018\ : Span4Mux_h
    port map (
            O => \N__40131\,
            I => \N__40124\
        );

    \I__8017\ : InMux
    port map (
            O => \N__40130\,
            I => \N__40121\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__40127\,
            I => pwm_counter_22
        );

    \I__8015\ : Odrv4
    port map (
            O => \N__40124\,
            I => pwm_counter_22
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__40121\,
            I => pwm_counter_22
        );

    \I__8013\ : InMux
    port map (
            O => \N__40114\,
            I => \PWM.n12707\
        );

    \I__8012\ : InMux
    port map (
            O => \N__40111\,
            I => \PWM.n12708\
        );

    \I__8011\ : InMux
    port map (
            O => \N__40108\,
            I => \N__40104\
        );

    \I__8010\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40101\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__40104\,
            I => pwm_counter_24
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__40101\,
            I => pwm_counter_24
        );

    \I__8007\ : InMux
    port map (
            O => \N__40096\,
            I => \bfn_11_32_0_\
        );

    \I__8006\ : InMux
    port map (
            O => \N__40093\,
            I => \N__40089\
        );

    \I__8005\ : InMux
    port map (
            O => \N__40092\,
            I => \N__40086\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__40089\,
            I => pwm_counter_25
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__40086\,
            I => pwm_counter_25
        );

    \I__8002\ : InMux
    port map (
            O => \N__40081\,
            I => \PWM.n12710\
        );

    \I__8001\ : InMux
    port map (
            O => \N__40078\,
            I => \N__40074\
        );

    \I__8000\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40071\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__40074\,
            I => pwm_counter_26
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__40071\,
            I => pwm_counter_26
        );

    \I__7997\ : InMux
    port map (
            O => \N__40066\,
            I => \PWM.n12711\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__40063\,
            I => \N__40059\
        );

    \I__7995\ : InMux
    port map (
            O => \N__40062\,
            I => \N__40056\
        );

    \I__7994\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40053\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__40056\,
            I => pwm_counter_27
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__40053\,
            I => pwm_counter_27
        );

    \I__7991\ : InMux
    port map (
            O => \N__40048\,
            I => \PWM.n12712\
        );

    \I__7990\ : InMux
    port map (
            O => \N__40045\,
            I => \N__40041\
        );

    \I__7989\ : InMux
    port map (
            O => \N__40044\,
            I => \N__40038\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__40041\,
            I => pwm_counter_28
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__40038\,
            I => pwm_counter_28
        );

    \I__7986\ : InMux
    port map (
            O => \N__40033\,
            I => \PWM.n12713\
        );

    \I__7985\ : InMux
    port map (
            O => \N__40030\,
            I => \PWM.n12697\
        );

    \I__7984\ : InMux
    port map (
            O => \N__40027\,
            I => \PWM.n12698\
        );

    \I__7983\ : InMux
    port map (
            O => \N__40024\,
            I => \PWM.n12699\
        );

    \I__7982\ : InMux
    port map (
            O => \N__40021\,
            I => \PWM.n12700\
        );

    \I__7981\ : InMux
    port map (
            O => \N__40018\,
            I => \bfn_11_31_0_\
        );

    \I__7980\ : InMux
    port map (
            O => \N__40015\,
            I => \PWM.n12702\
        );

    \I__7979\ : InMux
    port map (
            O => \N__40012\,
            I => \PWM.n12703\
        );

    \I__7978\ : InMux
    port map (
            O => \N__40009\,
            I => \PWM.n12704\
        );

    \I__7977\ : InMux
    port map (
            O => \N__40006\,
            I => \N__40001\
        );

    \I__7976\ : InMux
    port map (
            O => \N__40005\,
            I => \N__39996\
        );

    \I__7975\ : InMux
    port map (
            O => \N__40004\,
            I => \N__39996\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__40001\,
            I => pwm_counter_20
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__39996\,
            I => pwm_counter_20
        );

    \I__7972\ : InMux
    port map (
            O => \N__39991\,
            I => \PWM.n12705\
        );

    \I__7971\ : InMux
    port map (
            O => \N__39988\,
            I => \PWM.n12688\
        );

    \I__7970\ : InMux
    port map (
            O => \N__39985\,
            I => \N__39981\
        );

    \I__7969\ : InMux
    port map (
            O => \N__39984\,
            I => \N__39978\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__39981\,
            I => pwm_counter_4
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__39978\,
            I => pwm_counter_4
        );

    \I__7966\ : InMux
    port map (
            O => \N__39973\,
            I => \PWM.n12689\
        );

    \I__7965\ : InMux
    port map (
            O => \N__39970\,
            I => \PWM.n12690\
        );

    \I__7964\ : InMux
    port map (
            O => \N__39967\,
            I => \PWM.n12691\
        );

    \I__7963\ : InMux
    port map (
            O => \N__39964\,
            I => \PWM.n12692\
        );

    \I__7962\ : InMux
    port map (
            O => \N__39961\,
            I => \bfn_11_30_0_\
        );

    \I__7961\ : InMux
    port map (
            O => \N__39958\,
            I => \PWM.n12694\
        );

    \I__7960\ : InMux
    port map (
            O => \N__39955\,
            I => \PWM.n12695\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__39952\,
            I => \N__39948\
        );

    \I__7958\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39944\
        );

    \I__7957\ : InMux
    port map (
            O => \N__39948\,
            I => \N__39941\
        );

    \I__7956\ : InMux
    port map (
            O => \N__39947\,
            I => \N__39938\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__39944\,
            I => pwm_counter_11
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__39941\,
            I => pwm_counter_11
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__39938\,
            I => pwm_counter_11
        );

    \I__7952\ : InMux
    port map (
            O => \N__39931\,
            I => \PWM.n12696\
        );

    \I__7951\ : InMux
    port map (
            O => \N__39928\,
            I => \N__39925\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__39925\,
            I => \N__39922\
        );

    \I__7949\ : Span4Mux_h
    port map (
            O => \N__39922\,
            I => \N__39919\
        );

    \I__7948\ : Odrv4
    port map (
            O => \N__39919\,
            I => encoder0_position_scaled_14
        );

    \I__7947\ : InMux
    port map (
            O => \N__39916\,
            I => \N__39913\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__39913\,
            I => \N__39910\
        );

    \I__7945\ : Span4Mux_h
    port map (
            O => \N__39910\,
            I => \N__39907\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__39907\,
            I => encoder0_position_scaled_16
        );

    \I__7943\ : InMux
    port map (
            O => \N__39904\,
            I => \N__39901\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__39901\,
            I => \N__39898\
        );

    \I__7941\ : Span4Mux_h
    port map (
            O => \N__39898\,
            I => \N__39895\
        );

    \I__7940\ : Odrv4
    port map (
            O => \N__39895\,
            I => encoder0_position_scaled_18
        );

    \I__7939\ : InMux
    port map (
            O => \N__39892\,
            I => \N__39889\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__39889\,
            I => commutation_state_prev_2
        );

    \I__7937\ : InMux
    port map (
            O => \N__39886\,
            I => \bfn_11_29_0_\
        );

    \I__7936\ : InMux
    port map (
            O => \N__39883\,
            I => \PWM.n12686\
        );

    \I__7935\ : InMux
    port map (
            O => \N__39880\,
            I => \PWM.n12687\
        );

    \I__7934\ : InMux
    port map (
            O => \N__39877\,
            I => \N__39874\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__39874\,
            I => \N__39871\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__39871\,
            I => \N__39868\
        );

    \I__7931\ : Odrv4
    port map (
            O => \N__39868\,
            I => encoder0_position_scaled_7
        );

    \I__7930\ : InMux
    port map (
            O => \N__39865\,
            I => \N__39862\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__39862\,
            I => \N__39859\
        );

    \I__7928\ : Span4Mux_v
    port map (
            O => \N__39859\,
            I => \N__39856\
        );

    \I__7927\ : Odrv4
    port map (
            O => \N__39856\,
            I => encoder0_position_scaled_1
        );

    \I__7926\ : CascadeMux
    port map (
            O => \N__39853\,
            I => \n4_adj_698_cascade_\
        );

    \I__7925\ : InMux
    port map (
            O => \N__39850\,
            I => \N__39845\
        );

    \I__7924\ : InMux
    port map (
            O => \N__39849\,
            I => \N__39842\
        );

    \I__7923\ : InMux
    port map (
            O => \N__39848\,
            I => \N__39839\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__39845\,
            I => \N__39836\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__39842\,
            I => \N__39833\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__39839\,
            I => \N__39830\
        );

    \I__7919\ : Span4Mux_s3_v
    port map (
            O => \N__39836\,
            I => \N__39827\
        );

    \I__7918\ : Span4Mux_s2_v
    port map (
            O => \N__39833\,
            I => \N__39822\
        );

    \I__7917\ : Span4Mux_h
    port map (
            O => \N__39830\,
            I => \N__39822\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__39827\,
            I => pwm_setpoint_21
        );

    \I__7915\ : Odrv4
    port map (
            O => \N__39822\,
            I => pwm_setpoint_21
        );

    \I__7914\ : CascadeMux
    port map (
            O => \N__39817\,
            I => \n13856_cascade_\
        );

    \I__7913\ : CascadeMux
    port map (
            O => \N__39814\,
            I => \n13858_cascade_\
        );

    \I__7912\ : CascadeMux
    port map (
            O => \N__39811\,
            I => \n13860_cascade_\
        );

    \I__7911\ : CascadeMux
    port map (
            O => \N__39808\,
            I => \n13862_cascade_\
        );

    \I__7910\ : CascadeMux
    port map (
            O => \N__39805\,
            I => \n13864_cascade_\
        );

    \I__7909\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39799\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__39799\,
            I => n13866
        );

    \I__7907\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39793\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__39793\,
            I => \N__39790\
        );

    \I__7905\ : Span4Mux_h
    port map (
            O => \N__39790\,
            I => \N__39787\
        );

    \I__7904\ : Odrv4
    port map (
            O => \N__39787\,
            I => encoder0_position_scaled_5
        );

    \I__7903\ : InMux
    port map (
            O => \N__39784\,
            I => \N__39781\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__39781\,
            I => \N__39778\
        );

    \I__7901\ : Odrv4
    port map (
            O => \N__39778\,
            I => encoder0_position_scaled_8
        );

    \I__7900\ : InMux
    port map (
            O => \N__39775\,
            I => \N__39772\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__39772\,
            I => \N__39769\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__39769\,
            I => encoder0_position_scaled_11
        );

    \I__7897\ : CascadeMux
    port map (
            O => \N__39766\,
            I => \n3010_cascade_\
        );

    \I__7896\ : InMux
    port map (
            O => \N__39763\,
            I => \N__39760\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__39760\,
            I => \N__39757\
        );

    \I__7894\ : Span4Mux_h
    port map (
            O => \N__39757\,
            I => \N__39753\
        );

    \I__7893\ : InMux
    port map (
            O => \N__39756\,
            I => \N__39750\
        );

    \I__7892\ : Odrv4
    port map (
            O => \N__39753\,
            I => n15090
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__39750\,
            I => n15090
        );

    \I__7890\ : CascadeMux
    port map (
            O => \N__39745\,
            I => \n14392_cascade_\
        );

    \I__7889\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39739\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__39739\,
            I => \N__39736\
        );

    \I__7887\ : Odrv4
    port map (
            O => \N__39736\,
            I => n13470
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__39733\,
            I => \n14380_cascade_\
        );

    \I__7885\ : InMux
    port map (
            O => \N__39730\,
            I => \N__39727\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__39727\,
            I => n14386
        );

    \I__7883\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39721\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__39721\,
            I => n14398
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__39718\,
            I => \n3237_cascade_\
        );

    \I__7880\ : InMux
    port map (
            O => \N__39715\,
            I => \N__39712\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__39712\,
            I => n61
        );

    \I__7878\ : InMux
    port map (
            O => \N__39709\,
            I => \N__39706\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__39706\,
            I => n2981
        );

    \I__7876\ : InMux
    port map (
            O => \N__39703\,
            I => \N__39700\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__39700\,
            I => n2984
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__39697\,
            I => \n2912_cascade_\
        );

    \I__7873\ : InMux
    port map (
            O => \N__39694\,
            I => \N__39691\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__39691\,
            I => n2979
        );

    \I__7871\ : CascadeMux
    port map (
            O => \N__39688\,
            I => \N__39685\
        );

    \I__7870\ : InMux
    port map (
            O => \N__39685\,
            I => \N__39682\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__39682\,
            I => \N__39679\
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__39679\,
            I => n2975
        );

    \I__7867\ : CascadeMux
    port map (
            O => \N__39676\,
            I => \N__39673\
        );

    \I__7866\ : InMux
    port map (
            O => \N__39673\,
            I => \N__39670\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__39670\,
            I => n2980
        );

    \I__7864\ : CascadeMux
    port map (
            O => \N__39667\,
            I => \N__39664\
        );

    \I__7863\ : InMux
    port map (
            O => \N__39664\,
            I => \N__39661\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__39661\,
            I => n2976
        );

    \I__7861\ : InMux
    port map (
            O => \N__39658\,
            I => \N__39655\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__39655\,
            I => n2978
        );

    \I__7859\ : InMux
    port map (
            O => \N__39652\,
            I => \N__39649\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__39649\,
            I => n2998
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__39646\,
            I => \n3115_cascade_\
        );

    \I__7856\ : InMux
    port map (
            O => \N__39643\,
            I => \N__39640\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__39640\,
            I => n13894
        );

    \I__7854\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39634\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__39634\,
            I => \N__39631\
        );

    \I__7852\ : Span4Mux_v
    port map (
            O => \N__39631\,
            I => \N__39628\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__39628\,
            I => n13898
        );

    \I__7850\ : InMux
    port map (
            O => \N__39625\,
            I => \N__39622\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__39622\,
            I => n2988
        );

    \I__7848\ : InMux
    port map (
            O => \N__39619\,
            I => \N__39616\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__39616\,
            I => n2987
        );

    \I__7846\ : CascadeMux
    port map (
            O => \N__39613\,
            I => \n3019_cascade_\
        );

    \I__7845\ : CascadeMux
    port map (
            O => \N__39610\,
            I => \N__39607\
        );

    \I__7844\ : InMux
    port map (
            O => \N__39607\,
            I => \N__39604\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__39604\,
            I => n2983
        );

    \I__7842\ : CascadeMux
    port map (
            O => \N__39601\,
            I => \n2817_cascade_\
        );

    \I__7841\ : InMux
    port map (
            O => \N__39598\,
            I => \N__39595\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__39595\,
            I => n3000
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__39592\,
            I => \n3032_cascade_\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__39589\,
            I => \n11660_cascade_\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__39586\,
            I => \N__39583\
        );

    \I__7836\ : InMux
    port map (
            O => \N__39583\,
            I => \N__39580\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__39580\,
            I => \N__39577\
        );

    \I__7834\ : Odrv4
    port map (
            O => \N__39577\,
            I => n2986
        );

    \I__7833\ : InMux
    port map (
            O => \N__39574\,
            I => \N__39571\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__39571\,
            I => n2997
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__39568\,
            I => \n3029_cascade_\
        );

    \I__7830\ : InMux
    port map (
            O => \N__39565\,
            I => \N__39559\
        );

    \I__7829\ : InMux
    port map (
            O => \N__39564\,
            I => \N__39551\
        );

    \I__7828\ : InMux
    port map (
            O => \N__39563\,
            I => \N__39551\
        );

    \I__7827\ : InMux
    port map (
            O => \N__39562\,
            I => \N__39551\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__39559\,
            I => \N__39543\
        );

    \I__7825\ : InMux
    port map (
            O => \N__39558\,
            I => \N__39539\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__39551\,
            I => \N__39536\
        );

    \I__7823\ : InMux
    port map (
            O => \N__39550\,
            I => \N__39519\
        );

    \I__7822\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39519\
        );

    \I__7821\ : InMux
    port map (
            O => \N__39548\,
            I => \N__39519\
        );

    \I__7820\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39519\
        );

    \I__7819\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39513\
        );

    \I__7818\ : Span4Mux_h
    port map (
            O => \N__39543\,
            I => \N__39510\
        );

    \I__7817\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39507\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__39539\,
            I => \N__39504\
        );

    \I__7815\ : Span4Mux_v
    port map (
            O => \N__39536\,
            I => \N__39501\
        );

    \I__7814\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39498\
        );

    \I__7813\ : InMux
    port map (
            O => \N__39534\,
            I => \N__39493\
        );

    \I__7812\ : InMux
    port map (
            O => \N__39533\,
            I => \N__39490\
        );

    \I__7811\ : InMux
    port map (
            O => \N__39532\,
            I => \N__39487\
        );

    \I__7810\ : CascadeMux
    port map (
            O => \N__39531\,
            I => \N__39482\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__39530\,
            I => \N__39477\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__39529\,
            I => \N__39472\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__39528\,
            I => \N__39468\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__39519\,
            I => \N__39462\
        );

    \I__7805\ : InMux
    port map (
            O => \N__39518\,
            I => \N__39455\
        );

    \I__7804\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39455\
        );

    \I__7803\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39455\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__39513\,
            I => \N__39452\
        );

    \I__7801\ : Span4Mux_v
    port map (
            O => \N__39510\,
            I => \N__39449\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__39507\,
            I => \N__39446\
        );

    \I__7799\ : Span4Mux_v
    port map (
            O => \N__39504\,
            I => \N__39437\
        );

    \I__7798\ : Span4Mux_v
    port map (
            O => \N__39501\,
            I => \N__39437\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__39498\,
            I => \N__39434\
        );

    \I__7796\ : InMux
    port map (
            O => \N__39497\,
            I => \N__39429\
        );

    \I__7795\ : InMux
    port map (
            O => \N__39496\,
            I => \N__39429\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__39493\,
            I => \N__39422\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__39490\,
            I => \N__39422\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__39487\,
            I => \N__39422\
        );

    \I__7791\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39419\
        );

    \I__7790\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39408\
        );

    \I__7789\ : InMux
    port map (
            O => \N__39482\,
            I => \N__39408\
        );

    \I__7788\ : InMux
    port map (
            O => \N__39481\,
            I => \N__39408\
        );

    \I__7787\ : InMux
    port map (
            O => \N__39480\,
            I => \N__39408\
        );

    \I__7786\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39408\
        );

    \I__7785\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39397\
        );

    \I__7784\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39397\
        );

    \I__7783\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39397\
        );

    \I__7782\ : InMux
    port map (
            O => \N__39471\,
            I => \N__39397\
        );

    \I__7781\ : InMux
    port map (
            O => \N__39468\,
            I => \N__39397\
        );

    \I__7780\ : InMux
    port map (
            O => \N__39467\,
            I => \N__39391\
        );

    \I__7779\ : InMux
    port map (
            O => \N__39466\,
            I => \N__39386\
        );

    \I__7778\ : InMux
    port map (
            O => \N__39465\,
            I => \N__39386\
        );

    \I__7777\ : Span4Mux_v
    port map (
            O => \N__39462\,
            I => \N__39379\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__39455\,
            I => \N__39379\
        );

    \I__7775\ : Span4Mux_h
    port map (
            O => \N__39452\,
            I => \N__39379\
        );

    \I__7774\ : Span4Mux_h
    port map (
            O => \N__39449\,
            I => \N__39374\
        );

    \I__7773\ : Span4Mux_h
    port map (
            O => \N__39446\,
            I => \N__39374\
        );

    \I__7772\ : InMux
    port map (
            O => \N__39445\,
            I => \N__39367\
        );

    \I__7771\ : InMux
    port map (
            O => \N__39444\,
            I => \N__39367\
        );

    \I__7770\ : InMux
    port map (
            O => \N__39443\,
            I => \N__39367\
        );

    \I__7769\ : InMux
    port map (
            O => \N__39442\,
            I => \N__39364\
        );

    \I__7768\ : Span4Mux_h
    port map (
            O => \N__39437\,
            I => \N__39349\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__39434\,
            I => \N__39349\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__39429\,
            I => \N__39349\
        );

    \I__7765\ : Span4Mux_s3_v
    port map (
            O => \N__39422\,
            I => \N__39349\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39349\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__39408\,
            I => \N__39349\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__39397\,
            I => \N__39349\
        );

    \I__7761\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39342\
        );

    \I__7760\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39342\
        );

    \I__7759\ : InMux
    port map (
            O => \N__39394\,
            I => \N__39342\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__39391\,
            I => encoder0_position_31
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__39386\,
            I => encoder0_position_31
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__39379\,
            I => encoder0_position_31
        );

    \I__7755\ : Odrv4
    port map (
            O => \N__39374\,
            I => encoder0_position_31
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__39367\,
            I => encoder0_position_31
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__39364\,
            I => encoder0_position_31
        );

    \I__7752\ : Odrv4
    port map (
            O => \N__39349\,
            I => encoder0_position_31
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__39342\,
            I => encoder0_position_31
        );

    \I__7750\ : InMux
    port map (
            O => \N__39325\,
            I => \N__39322\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__39322\,
            I => \N__39319\
        );

    \I__7748\ : Span12Mux_v
    port map (
            O => \N__39319\,
            I => \N__39316\
        );

    \I__7747\ : Odrv12
    port map (
            O => \N__39316\,
            I => n29
        );

    \I__7746\ : InMux
    port map (
            O => \N__39313\,
            I => \N__39310\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__39310\,
            I => \N__39306\
        );

    \I__7744\ : CascadeMux
    port map (
            O => \N__39309\,
            I => \N__39303\
        );

    \I__7743\ : Span4Mux_v
    port map (
            O => \N__39306\,
            I => \N__39299\
        );

    \I__7742\ : InMux
    port map (
            O => \N__39303\,
            I => \N__39296\
        );

    \I__7741\ : InMux
    port map (
            O => \N__39302\,
            I => \N__39293\
        );

    \I__7740\ : Span4Mux_h
    port map (
            O => \N__39299\,
            I => \N__39290\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__39296\,
            I => \N__39287\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__39293\,
            I => encoder0_position_4
        );

    \I__7737\ : Odrv4
    port map (
            O => \N__39290\,
            I => encoder0_position_4
        );

    \I__7736\ : Odrv4
    port map (
            O => \N__39287\,
            I => encoder0_position_4
        );

    \I__7735\ : InMux
    port map (
            O => \N__39280\,
            I => \N__39277\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__39277\,
            I => n3001
        );

    \I__7733\ : CascadeMux
    port map (
            O => \N__39274\,
            I => \n315_cascade_\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__39271\,
            I => \n2714_cascade_\
        );

    \I__7731\ : CascadeMux
    port map (
            O => \N__39268\,
            I => \N__39265\
        );

    \I__7730\ : InMux
    port map (
            O => \N__39265\,
            I => \N__39261\
        );

    \I__7729\ : InMux
    port map (
            O => \N__39264\,
            I => \N__39258\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__39261\,
            I => \N__39255\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__39258\,
            I => \N__39251\
        );

    \I__7726\ : Span4Mux_h
    port map (
            O => \N__39255\,
            I => \N__39248\
        );

    \I__7725\ : InMux
    port map (
            O => \N__39254\,
            I => \N__39245\
        );

    \I__7724\ : Odrv12
    port map (
            O => \N__39251\,
            I => n2623
        );

    \I__7723\ : Odrv4
    port map (
            O => \N__39248\,
            I => n2623
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__39245\,
            I => n2623
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__39238\,
            I => \N__39235\
        );

    \I__7720\ : InMux
    port map (
            O => \N__39235\,
            I => \N__39232\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__39232\,
            I => \N__39229\
        );

    \I__7718\ : Span4Mux_v
    port map (
            O => \N__39229\,
            I => \N__39226\
        );

    \I__7717\ : Odrv4
    port map (
            O => \N__39226\,
            I => n2690
        );

    \I__7716\ : InMux
    port map (
            O => \N__39223\,
            I => \N__39220\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__39220\,
            I => \N__39217\
        );

    \I__7714\ : Span4Mux_h
    port map (
            O => \N__39217\,
            I => \N__39214\
        );

    \I__7713\ : Odrv4
    port map (
            O => \N__39214\,
            I => n2698
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__39211\,
            I => \N__39208\
        );

    \I__7711\ : InMux
    port map (
            O => \N__39208\,
            I => \N__39205\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__39205\,
            I => \N__39202\
        );

    \I__7709\ : Span4Mux_h
    port map (
            O => \N__39202\,
            I => \N__39199\
        );

    \I__7708\ : Odrv4
    port map (
            O => \N__39199\,
            I => n2699
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__39196\,
            I => \N__39192\
        );

    \I__7706\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39189\
        );

    \I__7705\ : InMux
    port map (
            O => \N__39192\,
            I => \N__39186\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__39189\,
            I => \N__39183\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__39186\,
            I => \N__39180\
        );

    \I__7702\ : Span4Mux_h
    port map (
            O => \N__39183\,
            I => \N__39174\
        );

    \I__7701\ : Span4Mux_v
    port map (
            O => \N__39180\,
            I => \N__39174\
        );

    \I__7700\ : InMux
    port map (
            O => \N__39179\,
            I => \N__39171\
        );

    \I__7699\ : Odrv4
    port map (
            O => \N__39174\,
            I => n2217
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__39171\,
            I => n2217
        );

    \I__7697\ : CascadeMux
    port map (
            O => \N__39166\,
            I => \N__39163\
        );

    \I__7696\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39160\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39157\
        );

    \I__7694\ : Span4Mux_h
    port map (
            O => \N__39157\,
            I => \N__39154\
        );

    \I__7693\ : Odrv4
    port map (
            O => \N__39154\,
            I => n2284
        );

    \I__7692\ : InMux
    port map (
            O => \N__39151\,
            I => \N__39146\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__39150\,
            I => \N__39140\
        );

    \I__7690\ : InMux
    port map (
            O => \N__39149\,
            I => \N__39135\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__39146\,
            I => \N__39129\
        );

    \I__7688\ : InMux
    port map (
            O => \N__39145\,
            I => \N__39126\
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__39144\,
            I => \N__39123\
        );

    \I__7686\ : CascadeMux
    port map (
            O => \N__39143\,
            I => \N__39120\
        );

    \I__7685\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39112\
        );

    \I__7684\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39112\
        );

    \I__7683\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39112\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__39135\,
            I => \N__39109\
        );

    \I__7681\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39106\
        );

    \I__7680\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39099\
        );

    \I__7679\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39099\
        );

    \I__7678\ : Span4Mux_h
    port map (
            O => \N__39129\,
            I => \N__39092\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__39126\,
            I => \N__39089\
        );

    \I__7676\ : InMux
    port map (
            O => \N__39123\,
            I => \N__39082\
        );

    \I__7675\ : InMux
    port map (
            O => \N__39120\,
            I => \N__39082\
        );

    \I__7674\ : InMux
    port map (
            O => \N__39119\,
            I => \N__39082\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__39112\,
            I => \N__39079\
        );

    \I__7672\ : Span4Mux_h
    port map (
            O => \N__39109\,
            I => \N__39076\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__39106\,
            I => \N__39073\
        );

    \I__7670\ : CascadeMux
    port map (
            O => \N__39105\,
            I => \N__39068\
        );

    \I__7669\ : InMux
    port map (
            O => \N__39104\,
            I => \N__39064\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__39099\,
            I => \N__39061\
        );

    \I__7667\ : InMux
    port map (
            O => \N__39098\,
            I => \N__39056\
        );

    \I__7666\ : InMux
    port map (
            O => \N__39097\,
            I => \N__39056\
        );

    \I__7665\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39051\
        );

    \I__7664\ : InMux
    port map (
            O => \N__39095\,
            I => \N__39051\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__39092\,
            I => \N__39042\
        );

    \I__7662\ : Span4Mux_h
    port map (
            O => \N__39089\,
            I => \N__39042\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__39082\,
            I => \N__39042\
        );

    \I__7660\ : Span4Mux_h
    port map (
            O => \N__39079\,
            I => \N__39042\
        );

    \I__7659\ : Span4Mux_h
    port map (
            O => \N__39076\,
            I => \N__39037\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__39073\,
            I => \N__39037\
        );

    \I__7657\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39028\
        );

    \I__7656\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39028\
        );

    \I__7655\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39028\
        );

    \I__7654\ : InMux
    port map (
            O => \N__39067\,
            I => \N__39028\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__39064\,
            I => n2247
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__39061\,
            I => n2247
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__39056\,
            I => n2247
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__39051\,
            I => n2247
        );

    \I__7649\ : Odrv4
    port map (
            O => \N__39042\,
            I => n2247
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__39037\,
            I => n2247
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__39028\,
            I => n2247
        );

    \I__7646\ : InMux
    port map (
            O => \N__39013\,
            I => \N__39008\
        );

    \I__7645\ : InMux
    port map (
            O => \N__39012\,
            I => \N__39005\
        );

    \I__7644\ : InMux
    port map (
            O => \N__39011\,
            I => \N__39002\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__39008\,
            I => \N__38995\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__39005\,
            I => \N__38995\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__39002\,
            I => \N__38995\
        );

    \I__7640\ : Span12Mux_s6_h
    port map (
            O => \N__38995\,
            I => \N__38992\
        );

    \I__7639\ : Odrv12
    port map (
            O => \N__38992\,
            I => n2316
        );

    \I__7638\ : InMux
    port map (
            O => \N__38989\,
            I => \N__38986\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__38986\,
            I => \N__38982\
        );

    \I__7636\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38979\
        );

    \I__7635\ : Span4Mux_h
    port map (
            O => \N__38982\,
            I => \N__38976\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__38979\,
            I => \N__38973\
        );

    \I__7633\ : Span4Mux_h
    port map (
            O => \N__38976\,
            I => \N__38970\
        );

    \I__7632\ : Span4Mux_v
    port map (
            O => \N__38973\,
            I => \N__38967\
        );

    \I__7631\ : Odrv4
    port map (
            O => \N__38970\,
            I => n2533
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__38967\,
            I => n2533
        );

    \I__7629\ : CascadeMux
    port map (
            O => \N__38962\,
            I => \N__38959\
        );

    \I__7628\ : InMux
    port map (
            O => \N__38959\,
            I => \N__38956\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__38956\,
            I => \N__38953\
        );

    \I__7626\ : Span4Mux_v
    port map (
            O => \N__38953\,
            I => \N__38950\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__38950\,
            I => \N__38947\
        );

    \I__7624\ : Odrv4
    port map (
            O => \N__38947\,
            I => n2600
        );

    \I__7623\ : InMux
    port map (
            O => \N__38944\,
            I => \N__38940\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__38943\,
            I => \N__38937\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__38940\,
            I => \N__38927\
        );

    \I__7620\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38924\
        );

    \I__7619\ : InMux
    port map (
            O => \N__38936\,
            I => \N__38919\
        );

    \I__7618\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38919\
        );

    \I__7617\ : InMux
    port map (
            O => \N__38934\,
            I => \N__38916\
        );

    \I__7616\ : CascadeMux
    port map (
            O => \N__38933\,
            I => \N__38913\
        );

    \I__7615\ : CascadeMux
    port map (
            O => \N__38932\,
            I => \N__38910\
        );

    \I__7614\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38904\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__38930\,
            I => \N__38901\
        );

    \I__7612\ : Span4Mux_v
    port map (
            O => \N__38927\,
            I => \N__38894\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__38924\,
            I => \N__38891\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__38919\,
            I => \N__38888\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__38916\,
            I => \N__38885\
        );

    \I__7608\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38874\
        );

    \I__7607\ : InMux
    port map (
            O => \N__38910\,
            I => \N__38874\
        );

    \I__7606\ : InMux
    port map (
            O => \N__38909\,
            I => \N__38874\
        );

    \I__7605\ : InMux
    port map (
            O => \N__38908\,
            I => \N__38874\
        );

    \I__7604\ : InMux
    port map (
            O => \N__38907\,
            I => \N__38874\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__38904\,
            I => \N__38871\
        );

    \I__7602\ : InMux
    port map (
            O => \N__38901\,
            I => \N__38863\
        );

    \I__7601\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38863\
        );

    \I__7600\ : CascadeMux
    port map (
            O => \N__38899\,
            I => \N__38857\
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__38898\,
            I => \N__38854\
        );

    \I__7598\ : CascadeMux
    port map (
            O => \N__38897\,
            I => \N__38851\
        );

    \I__7597\ : Span4Mux_v
    port map (
            O => \N__38894\,
            I => \N__38838\
        );

    \I__7596\ : Span4Mux_v
    port map (
            O => \N__38891\,
            I => \N__38838\
        );

    \I__7595\ : Span4Mux_v
    port map (
            O => \N__38888\,
            I => \N__38838\
        );

    \I__7594\ : Span4Mux_h
    port map (
            O => \N__38885\,
            I => \N__38838\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__38874\,
            I => \N__38838\
        );

    \I__7592\ : Span4Mux_h
    port map (
            O => \N__38871\,
            I => \N__38835\
        );

    \I__7591\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38828\
        );

    \I__7590\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38828\
        );

    \I__7589\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38828\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__38863\,
            I => \N__38825\
        );

    \I__7587\ : InMux
    port map (
            O => \N__38862\,
            I => \N__38820\
        );

    \I__7586\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38820\
        );

    \I__7585\ : InMux
    port map (
            O => \N__38860\,
            I => \N__38807\
        );

    \I__7584\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38807\
        );

    \I__7583\ : InMux
    port map (
            O => \N__38854\,
            I => \N__38807\
        );

    \I__7582\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38807\
        );

    \I__7581\ : InMux
    port map (
            O => \N__38850\,
            I => \N__38807\
        );

    \I__7580\ : InMux
    port map (
            O => \N__38849\,
            I => \N__38807\
        );

    \I__7579\ : Odrv4
    port map (
            O => \N__38838\,
            I => n2544
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__38835\,
            I => n2544
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__38828\,
            I => n2544
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__38825\,
            I => n2544
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__38820\,
            I => n2544
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__38807\,
            I => n2544
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__38794\,
            I => \N__38791\
        );

    \I__7572\ : InMux
    port map (
            O => \N__38791\,
            I => \N__38787\
        );

    \I__7571\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38784\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__38787\,
            I => \N__38781\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__38784\,
            I => n2632
        );

    \I__7568\ : Odrv4
    port map (
            O => \N__38781\,
            I => n2632
        );

    \I__7567\ : InMux
    port map (
            O => \N__38776\,
            I => \N__38771\
        );

    \I__7566\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38768\
        );

    \I__7565\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38765\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__38771\,
            I => \N__38762\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__38768\,
            I => \N__38759\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__38765\,
            I => \N__38756\
        );

    \I__7561\ : Span4Mux_v
    port map (
            O => \N__38762\,
            I => \N__38753\
        );

    \I__7560\ : Span4Mux_h
    port map (
            O => \N__38759\,
            I => \N__38748\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__38756\,
            I => \N__38748\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__38753\,
            I => \N__38745\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__38748\,
            I => \N__38742\
        );

    \I__7556\ : Odrv4
    port map (
            O => \N__38745\,
            I => n312
        );

    \I__7555\ : Odrv4
    port map (
            O => \N__38742\,
            I => n312
        );

    \I__7554\ : InMux
    port map (
            O => \N__38737\,
            I => \N__38733\
        );

    \I__7553\ : CascadeMux
    port map (
            O => \N__38736\,
            I => \N__38730\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__38733\,
            I => \N__38726\
        );

    \I__7551\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38723\
        );

    \I__7550\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38720\
        );

    \I__7549\ : Span4Mux_h
    port map (
            O => \N__38726\,
            I => \N__38717\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__38723\,
            I => \N__38712\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__38720\,
            I => \N__38712\
        );

    \I__7546\ : Odrv4
    port map (
            O => \N__38717\,
            I => n2633
        );

    \I__7545\ : Odrv12
    port map (
            O => \N__38712\,
            I => n2633
        );

    \I__7544\ : CascadeMux
    port map (
            O => \N__38707\,
            I => \n2632_cascade_\
        );

    \I__7543\ : InMux
    port map (
            O => \N__38704\,
            I => \N__38700\
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__38703\,
            I => \N__38697\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__38700\,
            I => \N__38693\
        );

    \I__7540\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38690\
        );

    \I__7539\ : InMux
    port map (
            O => \N__38696\,
            I => \N__38687\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__38693\,
            I => \N__38684\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__38690\,
            I => \N__38679\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__38687\,
            I => \N__38679\
        );

    \I__7535\ : Odrv4
    port map (
            O => \N__38684\,
            I => n2631
        );

    \I__7534\ : Odrv12
    port map (
            O => \N__38679\,
            I => n2631
        );

    \I__7533\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38671\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__38671\,
            I => \N__38668\
        );

    \I__7531\ : Span4Mux_v
    port map (
            O => \N__38668\,
            I => \N__38665\
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__38665\,
            I => n11760
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__38662\,
            I => \n2732_cascade_\
        );

    \I__7528\ : CascadeMux
    port map (
            O => \N__38659\,
            I => \n11666_cascade_\
        );

    \I__7527\ : InMux
    port map (
            O => \N__38656\,
            I => \N__38653\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__38653\,
            I => \N__38650\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__38650\,
            I => \N__38647\
        );

    \I__7524\ : Odrv4
    port map (
            O => \N__38647\,
            I => n2691
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__38644\,
            I => \N__38640\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__38643\,
            I => \N__38637\
        );

    \I__7521\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38634\
        );

    \I__7520\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38631\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__38634\,
            I => \N__38628\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__38631\,
            I => \N__38625\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__38628\,
            I => \N__38619\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__38625\,
            I => \N__38619\
        );

    \I__7515\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38616\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__38619\,
            I => n2624
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__38616\,
            I => n2624
        );

    \I__7512\ : InMux
    port map (
            O => \N__38611\,
            I => \N__38607\
        );

    \I__7511\ : InMux
    port map (
            O => \N__38610\,
            I => \N__38604\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__38607\,
            I => \N__38600\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__38604\,
            I => \N__38597\
        );

    \I__7508\ : InMux
    port map (
            O => \N__38603\,
            I => \N__38594\
        );

    \I__7507\ : Span4Mux_h
    port map (
            O => \N__38600\,
            I => \N__38591\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__38597\,
            I => \N__38586\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__38594\,
            I => \N__38586\
        );

    \I__7504\ : Odrv4
    port map (
            O => \N__38591\,
            I => n2617
        );

    \I__7503\ : Odrv4
    port map (
            O => \N__38586\,
            I => n2617
        );

    \I__7502\ : InMux
    port map (
            O => \N__38581\,
            I => \N__38578\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__38578\,
            I => \N__38575\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__38575\,
            I => \N__38572\
        );

    \I__7499\ : Odrv4
    port map (
            O => \N__38572\,
            I => n2684
        );

    \I__7498\ : InMux
    port map (
            O => \N__38569\,
            I => \N__38566\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__38566\,
            I => \N__38563\
        );

    \I__7496\ : Span4Mux_v
    port map (
            O => \N__38563\,
            I => \N__38560\
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__38560\,
            I => n2701
        );

    \I__7494\ : CascadeMux
    port map (
            O => \N__38557\,
            I => \N__38554\
        );

    \I__7493\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38551\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__38551\,
            I => \N__38546\
        );

    \I__7491\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38543\
        );

    \I__7490\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38540\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__38546\,
            I => \N__38537\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__38543\,
            I => \N__38532\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__38540\,
            I => \N__38532\
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__38537\,
            I => n2613
        );

    \I__7485\ : Odrv12
    port map (
            O => \N__38532\,
            I => n2613
        );

    \I__7484\ : CascadeMux
    port map (
            O => \N__38527\,
            I => \N__38524\
        );

    \I__7483\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38521\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__38521\,
            I => \N__38518\
        );

    \I__7481\ : Span4Mux_h
    port map (
            O => \N__38518\,
            I => \N__38515\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__38515\,
            I => n2680
        );

    \I__7479\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38508\
        );

    \I__7478\ : InMux
    port map (
            O => \N__38511\,
            I => \N__38505\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__38508\,
            I => \N__38501\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__38505\,
            I => \N__38498\
        );

    \I__7475\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38495\
        );

    \I__7474\ : Span4Mux_h
    port map (
            O => \N__38501\,
            I => \N__38492\
        );

    \I__7473\ : Span4Mux_h
    port map (
            O => \N__38498\,
            I => \N__38487\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__38495\,
            I => \N__38487\
        );

    \I__7471\ : Odrv4
    port map (
            O => \N__38492\,
            I => n2611
        );

    \I__7470\ : Odrv4
    port map (
            O => \N__38487\,
            I => n2611
        );

    \I__7469\ : InMux
    port map (
            O => \N__38482\,
            I => \N__38479\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__38479\,
            I => \N__38476\
        );

    \I__7467\ : Span4Mux_h
    port map (
            O => \N__38476\,
            I => \N__38473\
        );

    \I__7466\ : Odrv4
    port map (
            O => \N__38473\,
            I => n2678
        );

    \I__7465\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38465\
        );

    \I__7464\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38462\
        );

    \I__7463\ : CascadeMux
    port map (
            O => \N__38468\,
            I => \N__38459\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__38465\,
            I => \N__38456\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__38462\,
            I => \N__38453\
        );

    \I__7460\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38450\
        );

    \I__7459\ : Span4Mux_v
    port map (
            O => \N__38456\,
            I => \N__38447\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__38453\,
            I => \N__38442\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__38450\,
            I => \N__38442\
        );

    \I__7456\ : Odrv4
    port map (
            O => \N__38447\,
            I => n2615
        );

    \I__7455\ : Odrv4
    port map (
            O => \N__38442\,
            I => n2615
        );

    \I__7454\ : CascadeMux
    port map (
            O => \N__38437\,
            I => \N__38434\
        );

    \I__7453\ : InMux
    port map (
            O => \N__38434\,
            I => \N__38431\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__38431\,
            I => \N__38428\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__38428\,
            I => \N__38425\
        );

    \I__7450\ : Odrv4
    port map (
            O => \N__38425\,
            I => n2682
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__38422\,
            I => \n45_cascade_\
        );

    \I__7448\ : InMux
    port map (
            O => \N__38419\,
            I => \N__38416\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__38416\,
            I => n16_adj_614
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__38413\,
            I => \n14843_cascade_\
        );

    \I__7445\ : InMux
    port map (
            O => \N__38410\,
            I => \N__38407\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__38407\,
            I => n24_adj_619
        );

    \I__7443\ : CascadeMux
    port map (
            O => \N__38404\,
            I => \n14711_cascade_\
        );

    \I__7442\ : InMux
    port map (
            O => \N__38401\,
            I => \N__38398\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__38398\,
            I => n8_adj_607
        );

    \I__7440\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38390\
        );

    \I__7439\ : InMux
    port map (
            O => \N__38394\,
            I => \N__38385\
        );

    \I__7438\ : InMux
    port map (
            O => \N__38393\,
            I => \N__38385\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__38390\,
            I => n45
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__38385\,
            I => n45
        );

    \I__7435\ : CascadeMux
    port map (
            O => \N__38380\,
            I => \n14826_cascade_\
        );

    \I__7434\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38374\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__38374\,
            I => n14779
        );

    \I__7432\ : InMux
    port map (
            O => \N__38371\,
            I => \N__38368\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__38368\,
            I => \N__38365\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__38365\,
            I => n14864
        );

    \I__7429\ : CascadeMux
    port map (
            O => \N__38362\,
            I => \N__38359\
        );

    \I__7428\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38355\
        );

    \I__7427\ : InMux
    port map (
            O => \N__38358\,
            I => \N__38352\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__38355\,
            I => n43
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__38352\,
            I => n43
        );

    \I__7424\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38344\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__38344\,
            I => n14713
        );

    \I__7422\ : InMux
    port map (
            O => \N__38341\,
            I => \N__38338\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__38338\,
            I => \N__38335\
        );

    \I__7420\ : Span4Mux_h
    port map (
            O => \N__38335\,
            I => \N__38332\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__38332\,
            I => n2700
        );

    \I__7418\ : CascadeMux
    port map (
            O => \N__38329\,
            I => \n41_cascade_\
        );

    \I__7417\ : InMux
    port map (
            O => \N__38326\,
            I => \N__38323\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__38323\,
            I => n41
        );

    \I__7415\ : CascadeMux
    port map (
            O => \N__38320\,
            I => \n14715_cascade_\
        );

    \I__7414\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38314\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__38314\,
            I => n40
        );

    \I__7412\ : CascadeMux
    port map (
            O => \N__38311\,
            I => \n14866_cascade_\
        );

    \I__7411\ : CascadeMux
    port map (
            O => \N__38308\,
            I => \n12_adj_598_cascade_\
        );

    \I__7410\ : InMux
    port map (
            O => \N__38305\,
            I => \N__38301\
        );

    \I__7409\ : InMux
    port map (
            O => \N__38304\,
            I => \N__38298\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__38301\,
            I => \N__38294\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__38298\,
            I => \N__38291\
        );

    \I__7406\ : InMux
    port map (
            O => \N__38297\,
            I => \N__38288\
        );

    \I__7405\ : Span4Mux_v
    port map (
            O => \N__38294\,
            I => \N__38283\
        );

    \I__7404\ : Span4Mux_v
    port map (
            O => \N__38291\,
            I => \N__38283\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__38288\,
            I => encoder0_position_13
        );

    \I__7402\ : Odrv4
    port map (
            O => \N__38283\,
            I => encoder0_position_13
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__38278\,
            I => \N__38275\
        );

    \I__7400\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38272\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__38272\,
            I => \N__38269\
        );

    \I__7398\ : Span4Mux_h
    port map (
            O => \N__38269\,
            I => \N__38266\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__38266\,
            I => n20_adj_644
        );

    \I__7396\ : InMux
    port map (
            O => \N__38263\,
            I => \N__38258\
        );

    \I__7395\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38252\
        );

    \I__7394\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38252\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__38258\,
            I => \N__38249\
        );

    \I__7392\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38246\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__38252\,
            I => \N__38243\
        );

    \I__7390\ : Span4Mux_h
    port map (
            O => \N__38249\,
            I => \N__38240\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__38246\,
            I => encoder0_position_28
        );

    \I__7388\ : Odrv4
    port map (
            O => \N__38243\,
            I => encoder0_position_28
        );

    \I__7387\ : Odrv4
    port map (
            O => \N__38240\,
            I => encoder0_position_28
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__38233\,
            I => \N__38230\
        );

    \I__7385\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38227\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38224\
        );

    \I__7383\ : Odrv4
    port map (
            O => \N__38224\,
            I => n5_adj_629
        );

    \I__7382\ : InMux
    port map (
            O => \N__38221\,
            I => \N__38218\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__38218\,
            I => \N__38215\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__38215\,
            I => encoder0_position_scaled_9
        );

    \I__7379\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38209\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__38209\,
            I => \N__38206\
        );

    \I__7377\ : Odrv4
    port map (
            O => \N__38206\,
            I => encoder0_position_scaled_10
        );

    \I__7376\ : CascadeMux
    port map (
            O => \N__38203\,
            I => \N__38200\
        );

    \I__7375\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38193\
        );

    \I__7374\ : InMux
    port map (
            O => \N__38199\,
            I => \N__38193\
        );

    \I__7373\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38188\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__38193\,
            I => \N__38185\
        );

    \I__7371\ : InMux
    port map (
            O => \N__38192\,
            I => \N__38182\
        );

    \I__7370\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38179\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__38188\,
            I => \N__38172\
        );

    \I__7368\ : Span4Mux_h
    port map (
            O => \N__38185\,
            I => \N__38172\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__38182\,
            I => \N__38172\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__38179\,
            I => \N__38166\
        );

    \I__7365\ : Span4Mux_v
    port map (
            O => \N__38172\,
            I => \N__38166\
        );

    \I__7364\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38163\
        );

    \I__7363\ : Span4Mux_h
    port map (
            O => \N__38166\,
            I => \N__38160\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__38163\,
            I => h2
        );

    \I__7361\ : Odrv4
    port map (
            O => \N__38160\,
            I => h2
        );

    \I__7360\ : InMux
    port map (
            O => \N__38155\,
            I => \N__38151\
        );

    \I__7359\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38145\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__38151\,
            I => \N__38142\
        );

    \I__7357\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38139\
        );

    \I__7356\ : InMux
    port map (
            O => \N__38149\,
            I => \N__38136\
        );

    \I__7355\ : InMux
    port map (
            O => \N__38148\,
            I => \N__38133\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__38145\,
            I => \N__38129\
        );

    \I__7353\ : Span4Mux_s2_v
    port map (
            O => \N__38142\,
            I => \N__38126\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__38139\,
            I => \N__38119\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__38136\,
            I => \N__38119\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__38133\,
            I => \N__38119\
        );

    \I__7349\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38116\
        );

    \I__7348\ : Span12Mux_s6_v
    port map (
            O => \N__38129\,
            I => \N__38113\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__38126\,
            I => \N__38110\
        );

    \I__7346\ : Span4Mux_v
    port map (
            O => \N__38119\,
            I => \N__38107\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__38116\,
            I => h3
        );

    \I__7344\ : Odrv12
    port map (
            O => \N__38113\,
            I => h3
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__38110\,
            I => h3
        );

    \I__7342\ : Odrv4
    port map (
            O => \N__38107\,
            I => h3
        );

    \I__7341\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38092\
        );

    \I__7340\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38089\
        );

    \I__7339\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38083\
        );

    \I__7338\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38083\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__38092\,
            I => \N__38080\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__38089\,
            I => \N__38077\
        );

    \I__7335\ : InMux
    port map (
            O => \N__38088\,
            I => \N__38074\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__38083\,
            I => \N__38071\
        );

    \I__7333\ : Span4Mux_h
    port map (
            O => \N__38080\,
            I => \N__38065\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__38077\,
            I => \N__38065\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__38074\,
            I => \N__38062\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__38071\,
            I => \N__38059\
        );

    \I__7329\ : InMux
    port map (
            O => \N__38070\,
            I => \N__38056\
        );

    \I__7328\ : Span4Mux_h
    port map (
            O => \N__38065\,
            I => \N__38053\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__38062\,
            I => \N__38048\
        );

    \I__7326\ : Span4Mux_h
    port map (
            O => \N__38059\,
            I => \N__38048\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__38056\,
            I => h1
        );

    \I__7324\ : Odrv4
    port map (
            O => \N__38053\,
            I => h1
        );

    \I__7323\ : Odrv4
    port map (
            O => \N__38048\,
            I => h1
        );

    \I__7322\ : CEMux
    port map (
            O => \N__38041\,
            I => \N__38038\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__38038\,
            I => \N__38035\
        );

    \I__7320\ : Span4Mux_v
    port map (
            O => \N__38035\,
            I => \N__38032\
        );

    \I__7319\ : Odrv4
    port map (
            O => \N__38032\,
            I => n6_adj_592
        );

    \I__7318\ : SRMux
    port map (
            O => \N__38029\,
            I => \N__38026\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38023\
        );

    \I__7316\ : Span4Mux_h
    port map (
            O => \N__38023\,
            I => \N__38020\
        );

    \I__7315\ : Odrv4
    port map (
            O => \N__38020\,
            I => \commutation_state_7__N_261\
        );

    \I__7314\ : InMux
    port map (
            O => \N__38017\,
            I => \N__38014\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__38014\,
            I => encoder0_position_scaled_4
        );

    \I__7312\ : CascadeMux
    port map (
            O => \N__38011\,
            I => \dti_N_333_cascade_\
        );

    \I__7311\ : InMux
    port map (
            O => \N__38008\,
            I => \N__38005\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__38005\,
            I => encoder0_position_scaled_22
        );

    \I__7309\ : InMux
    port map (
            O => \N__38002\,
            I => \N__37999\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__37999\,
            I => \N__37996\
        );

    \I__7307\ : Span4Mux_h
    port map (
            O => \N__37996\,
            I => \N__37993\
        );

    \I__7306\ : Odrv4
    port map (
            O => \N__37993\,
            I => n26
        );

    \I__7305\ : InMux
    port map (
            O => \N__37990\,
            I => \N__37987\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__37987\,
            I => \N__37983\
        );

    \I__7303\ : CascadeMux
    port map (
            O => \N__37986\,
            I => \N__37980\
        );

    \I__7302\ : Span4Mux_h
    port map (
            O => \N__37983\,
            I => \N__37977\
        );

    \I__7301\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37973\
        );

    \I__7300\ : Span4Mux_v
    port map (
            O => \N__37977\,
            I => \N__37970\
        );

    \I__7299\ : InMux
    port map (
            O => \N__37976\,
            I => \N__37967\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__37973\,
            I => encoder0_position_7
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__37970\,
            I => encoder0_position_7
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__37967\,
            I => encoder0_position_7
        );

    \I__7295\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37957\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__37957\,
            I => encoder0_position_scaled_19
        );

    \I__7293\ : InMux
    port map (
            O => \N__37954\,
            I => \N__37951\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__37951\,
            I => encoder0_position_scaled_21
        );

    \I__7291\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37945\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__37945\,
            I => encoder0_position_scaled_13
        );

    \I__7289\ : CEMux
    port map (
            O => \N__37942\,
            I => \N__37939\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__37939\,
            I => \N__37936\
        );

    \I__7287\ : Span4Mux_h
    port map (
            O => \N__37936\,
            I => \N__37933\
        );

    \I__7286\ : Odrv4
    port map (
            O => \N__37933\,
            I => n4828
        );

    \I__7285\ : CascadeMux
    port map (
            O => \N__37930\,
            I => \n11593_cascade_\
        );

    \I__7284\ : CascadeMux
    port map (
            O => \N__37927\,
            I => \n59_cascade_\
        );

    \I__7283\ : CascadeMux
    port map (
            O => \N__37924\,
            I => \N__37920\
        );

    \I__7282\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37917\
        );

    \I__7281\ : InMux
    port map (
            O => \N__37920\,
            I => \N__37914\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__37917\,
            I => n11838
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__37914\,
            I => n11838
        );

    \I__7278\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37906\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__37906\,
            I => encoder0_position_scaled_0
        );

    \I__7276\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37900\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__37900\,
            I => encoder0_position_scaled_15
        );

    \I__7274\ : InMux
    port map (
            O => \N__37897\,
            I => \N__37894\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__37894\,
            I => encoder0_position_scaled_12
        );

    \I__7272\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37888\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__37888\,
            I => encoder0_position_scaled_2
        );

    \I__7270\ : InMux
    port map (
            O => \N__37885\,
            I => n12461
        );

    \I__7269\ : InMux
    port map (
            O => \N__37882\,
            I => n12462
        );

    \I__7268\ : InMux
    port map (
            O => \N__37879\,
            I => n12463
        );

    \I__7267\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37873\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__37873\,
            I => n15197
        );

    \I__7265\ : InMux
    port map (
            O => \N__37870\,
            I => \bfn_10_23_0_\
        );

    \I__7264\ : InMux
    port map (
            O => \N__37867\,
            I => n12453
        );

    \I__7263\ : InMux
    port map (
            O => \N__37864\,
            I => n12454
        );

    \I__7262\ : InMux
    port map (
            O => \N__37861\,
            I => n12455
        );

    \I__7261\ : InMux
    port map (
            O => \N__37858\,
            I => n12456
        );

    \I__7260\ : InMux
    port map (
            O => \N__37855\,
            I => n12457
        );

    \I__7259\ : InMux
    port map (
            O => \N__37852\,
            I => n12458
        );

    \I__7258\ : InMux
    port map (
            O => \N__37849\,
            I => n12459
        );

    \I__7257\ : InMux
    port map (
            O => \N__37846\,
            I => \bfn_10_24_0_\
        );

    \I__7256\ : InMux
    port map (
            O => \N__37843\,
            I => n12443
        );

    \I__7255\ : InMux
    port map (
            O => \N__37840\,
            I => \bfn_10_22_0_\
        );

    \I__7254\ : InMux
    port map (
            O => \N__37837\,
            I => n12445
        );

    \I__7253\ : InMux
    port map (
            O => \N__37834\,
            I => n12446
        );

    \I__7252\ : InMux
    port map (
            O => \N__37831\,
            I => n12447
        );

    \I__7251\ : InMux
    port map (
            O => \N__37828\,
            I => n12448
        );

    \I__7250\ : InMux
    port map (
            O => \N__37825\,
            I => n12449
        );

    \I__7249\ : InMux
    port map (
            O => \N__37822\,
            I => n12450
        );

    \I__7248\ : InMux
    port map (
            O => \N__37819\,
            I => n12451
        );

    \I__7247\ : CascadeMux
    port map (
            O => \N__37816\,
            I => \n3117_cascade_\
        );

    \I__7246\ : InMux
    port map (
            O => \N__37813\,
            I => \N__37810\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__37810\,
            I => n13888
        );

    \I__7244\ : InMux
    port map (
            O => \N__37807\,
            I => \N__37804\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__37804\,
            I => n13886
        );

    \I__7242\ : InMux
    port map (
            O => \N__37801\,
            I => \bfn_10_21_0_\
        );

    \I__7241\ : InMux
    port map (
            O => \N__37798\,
            I => n12437
        );

    \I__7240\ : InMux
    port map (
            O => \N__37795\,
            I => n12438
        );

    \I__7239\ : InMux
    port map (
            O => \N__37792\,
            I => n12439
        );

    \I__7238\ : InMux
    port map (
            O => \N__37789\,
            I => n12440
        );

    \I__7237\ : InMux
    port map (
            O => \N__37786\,
            I => n12441
        );

    \I__7236\ : InMux
    port map (
            O => \N__37783\,
            I => n12442
        );

    \I__7235\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37777\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__37777\,
            I => \N__37773\
        );

    \I__7233\ : InMux
    port map (
            O => \N__37776\,
            I => \N__37769\
        );

    \I__7232\ : Span4Mux_h
    port map (
            O => \N__37773\,
            I => \N__37766\
        );

    \I__7231\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37763\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__37769\,
            I => \N__37758\
        );

    \I__7229\ : Span4Mux_v
    port map (
            O => \N__37766\,
            I => \N__37758\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__37763\,
            I => encoder0_position_6
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__37758\,
            I => encoder0_position_6
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__37753\,
            I => \N__37750\
        );

    \I__7225\ : InMux
    port map (
            O => \N__37750\,
            I => \N__37747\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__37747\,
            I => \N__37744\
        );

    \I__7223\ : Span4Mux_v
    port map (
            O => \N__37744\,
            I => \N__37741\
        );

    \I__7222\ : Span4Mux_h
    port map (
            O => \N__37741\,
            I => \N__37738\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__37738\,
            I => n27_adj_651
        );

    \I__7220\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37732\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__37732\,
            I => \N__37729\
        );

    \I__7218\ : Span4Mux_v
    port map (
            O => \N__37729\,
            I => \N__37726\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__37726\,
            I => \N__37723\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__37723\,
            I => n24
        );

    \I__7215\ : InMux
    port map (
            O => \N__37720\,
            I => \N__37717\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__37717\,
            I => \N__37714\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__37714\,
            I => \N__37709\
        );

    \I__7212\ : InMux
    port map (
            O => \N__37713\,
            I => \N__37706\
        );

    \I__7211\ : InMux
    port map (
            O => \N__37712\,
            I => \N__37703\
        );

    \I__7210\ : Span4Mux_h
    port map (
            O => \N__37709\,
            I => \N__37700\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__37706\,
            I => \N__37697\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__37703\,
            I => encoder0_position_9
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__37700\,
            I => encoder0_position_9
        );

    \I__7206\ : Odrv12
    port map (
            O => \N__37697\,
            I => encoder0_position_9
        );

    \I__7205\ : InMux
    port map (
            O => \N__37690\,
            I => \N__37687\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__37687\,
            I => \N__37683\
        );

    \I__7203\ : InMux
    port map (
            O => \N__37686\,
            I => \N__37680\
        );

    \I__7202\ : Span4Mux_v
    port map (
            O => \N__37683\,
            I => \N__37674\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__37680\,
            I => \N__37674\
        );

    \I__7200\ : InMux
    port map (
            O => \N__37679\,
            I => \N__37671\
        );

    \I__7199\ : Span4Mux_h
    port map (
            O => \N__37674\,
            I => \N__37668\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__37671\,
            I => \N__37665\
        );

    \I__7197\ : Span4Mux_h
    port map (
            O => \N__37668\,
            I => \N__37662\
        );

    \I__7196\ : Span12Mux_s9_h
    port map (
            O => \N__37665\,
            I => \N__37659\
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__37662\,
            I => n310
        );

    \I__7194\ : Odrv12
    port map (
            O => \N__37659\,
            I => n310
        );

    \I__7193\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37651\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__37651\,
            I => \N__37648\
        );

    \I__7191\ : Span4Mux_v
    port map (
            O => \N__37648\,
            I => \N__37645\
        );

    \I__7190\ : Span4Mux_v
    port map (
            O => \N__37645\,
            I => \N__37642\
        );

    \I__7189\ : Span4Mux_h
    port map (
            O => \N__37642\,
            I => \N__37639\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__37639\,
            I => n19
        );

    \I__7187\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37633\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__37633\,
            I => \N__37629\
        );

    \I__7185\ : CascadeMux
    port map (
            O => \N__37632\,
            I => \N__37625\
        );

    \I__7184\ : Span4Mux_h
    port map (
            O => \N__37629\,
            I => \N__37622\
        );

    \I__7183\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37619\
        );

    \I__7182\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37616\
        );

    \I__7181\ : Span4Mux_v
    port map (
            O => \N__37622\,
            I => \N__37613\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__37619\,
            I => \N__37610\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__37616\,
            I => encoder0_position_14
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__37613\,
            I => encoder0_position_14
        );

    \I__7177\ : Odrv4
    port map (
            O => \N__37610\,
            I => encoder0_position_14
        );

    \I__7176\ : InMux
    port map (
            O => \N__37603\,
            I => \N__37600\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__37600\,
            I => \N__37595\
        );

    \I__7174\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37592\
        );

    \I__7173\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37589\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__37595\,
            I => \N__37586\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__37592\,
            I => \N__37581\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__37589\,
            I => \N__37581\
        );

    \I__7169\ : Span4Mux_h
    port map (
            O => \N__37586\,
            I => \N__37576\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__37581\,
            I => \N__37576\
        );

    \I__7167\ : Span4Mux_h
    port map (
            O => \N__37576\,
            I => \N__37573\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__37573\,
            I => n305
        );

    \I__7165\ : InMux
    port map (
            O => \N__37570\,
            I => \N__37567\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__37567\,
            I => \N__37564\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__37564\,
            I => \N__37561\
        );

    \I__7162\ : Span4Mux_v
    port map (
            O => \N__37561\,
            I => \N__37558\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__37558\,
            I => n23
        );

    \I__7160\ : InMux
    port map (
            O => \N__37555\,
            I => \N__37551\
        );

    \I__7159\ : InMux
    port map (
            O => \N__37554\,
            I => \N__37548\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__37551\,
            I => \N__37544\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__37548\,
            I => \N__37541\
        );

    \I__7156\ : CascadeMux
    port map (
            O => \N__37547\,
            I => \N__37538\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__37544\,
            I => \N__37535\
        );

    \I__7154\ : Span4Mux_v
    port map (
            O => \N__37541\,
            I => \N__37532\
        );

    \I__7153\ : InMux
    port map (
            O => \N__37538\,
            I => \N__37529\
        );

    \I__7152\ : Span4Mux_v
    port map (
            O => \N__37535\,
            I => \N__37526\
        );

    \I__7151\ : Span4Mux_v
    port map (
            O => \N__37532\,
            I => \N__37523\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__37529\,
            I => encoder0_position_10
        );

    \I__7149\ : Odrv4
    port map (
            O => \N__37526\,
            I => encoder0_position_10
        );

    \I__7148\ : Odrv4
    port map (
            O => \N__37523\,
            I => encoder0_position_10
        );

    \I__7147\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37513\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__37513\,
            I => \N__37509\
        );

    \I__7145\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37506\
        );

    \I__7144\ : Span4Mux_v
    port map (
            O => \N__37509\,
            I => \N__37500\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__37506\,
            I => \N__37500\
        );

    \I__7142\ : InMux
    port map (
            O => \N__37505\,
            I => \N__37497\
        );

    \I__7141\ : Span4Mux_h
    port map (
            O => \N__37500\,
            I => \N__37494\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__37497\,
            I => \N__37491\
        );

    \I__7139\ : Span4Mux_h
    port map (
            O => \N__37494\,
            I => \N__37488\
        );

    \I__7138\ : Odrv12
    port map (
            O => \N__37491\,
            I => n309
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__37488\,
            I => n309
        );

    \I__7136\ : CascadeMux
    port map (
            O => \N__37483\,
            I => \N__37479\
        );

    \I__7135\ : InMux
    port map (
            O => \N__37482\,
            I => \N__37476\
        );

    \I__7134\ : InMux
    port map (
            O => \N__37479\,
            I => \N__37473\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__37476\,
            I => \N__37467\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37467\
        );

    \I__7131\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37464\
        );

    \I__7130\ : Span4Mux_v
    port map (
            O => \N__37467\,
            I => \N__37459\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__37464\,
            I => \N__37459\
        );

    \I__7128\ : Odrv4
    port map (
            O => \N__37459\,
            I => n2616
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__37456\,
            I => \N__37453\
        );

    \I__7126\ : InMux
    port map (
            O => \N__37453\,
            I => \N__37450\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__37450\,
            I => \N__37447\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__37447\,
            I => n2683
        );

    \I__7123\ : CascadeMux
    port map (
            O => \N__37444\,
            I => \n13884_cascade_\
        );

    \I__7122\ : CascadeMux
    port map (
            O => \N__37441\,
            I => \N__37437\
        );

    \I__7121\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37434\
        );

    \I__7120\ : InMux
    port map (
            O => \N__37437\,
            I => \N__37431\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37426\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__37431\,
            I => \N__37426\
        );

    \I__7117\ : Span4Mux_v
    port map (
            O => \N__37426\,
            I => \N__37422\
        );

    \I__7116\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37419\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__37422\,
            I => n2627
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__37419\,
            I => n2627
        );

    \I__7113\ : CascadeMux
    port map (
            O => \N__37414\,
            I => \N__37411\
        );

    \I__7112\ : InMux
    port map (
            O => \N__37411\,
            I => \N__37408\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__37408\,
            I => n2694
        );

    \I__7110\ : InMux
    port map (
            O => \N__37405\,
            I => \N__37401\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__37404\,
            I => \N__37398\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__37401\,
            I => \N__37395\
        );

    \I__7107\ : InMux
    port map (
            O => \N__37398\,
            I => \N__37392\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__37395\,
            I => \N__37388\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__37392\,
            I => \N__37385\
        );

    \I__7104\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37382\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__37388\,
            I => n2521
        );

    \I__7102\ : Odrv4
    port map (
            O => \N__37385\,
            I => n2521
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__37382\,
            I => n2521
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__37375\,
            I => \N__37372\
        );

    \I__7099\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37369\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__37369\,
            I => \N__37366\
        );

    \I__7097\ : Span4Mux_v
    port map (
            O => \N__37366\,
            I => \N__37363\
        );

    \I__7096\ : Odrv4
    port map (
            O => \N__37363\,
            I => n2588
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__37360\,
            I => \N__37357\
        );

    \I__7094\ : InMux
    port map (
            O => \N__37357\,
            I => \N__37354\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__37354\,
            I => \N__37350\
        );

    \I__7092\ : InMux
    port map (
            O => \N__37353\,
            I => \N__37347\
        );

    \I__7091\ : Odrv4
    port map (
            O => \N__37350\,
            I => n2620
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__37347\,
            I => n2620
        );

    \I__7089\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37339\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__37339\,
            I => \N__37336\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__37336\,
            I => n2687
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__37333\,
            I => \n2620_cascade_\
        );

    \I__7085\ : InMux
    port map (
            O => \N__37330\,
            I => \N__37327\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__37327\,
            I => \N__37323\
        );

    \I__7083\ : InMux
    port map (
            O => \N__37326\,
            I => \N__37320\
        );

    \I__7082\ : Span4Mux_h
    port map (
            O => \N__37323\,
            I => \N__37317\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__37320\,
            I => \N__37314\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__37317\,
            I => \N__37309\
        );

    \I__7079\ : Span4Mux_h
    port map (
            O => \N__37314\,
            I => \N__37309\
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__37309\,
            I => n2610
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__37306\,
            I => \N__37303\
        );

    \I__7076\ : InMux
    port map (
            O => \N__37303\,
            I => \N__37300\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__37300\,
            I => n14300
        );

    \I__7074\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37293\
        );

    \I__7073\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37289\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__37293\,
            I => \N__37286\
        );

    \I__7071\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37283\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__37289\,
            I => n2621
        );

    \I__7069\ : Odrv4
    port map (
            O => \N__37286\,
            I => n2621
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__37283\,
            I => n2621
        );

    \I__7067\ : CascadeMux
    port map (
            O => \N__37276\,
            I => \n2643_cascade_\
        );

    \I__7066\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37270\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__37270\,
            I => \N__37267\
        );

    \I__7064\ : Span4Mux_v
    port map (
            O => \N__37267\,
            I => \N__37264\
        );

    \I__7063\ : Span4Mux_h
    port map (
            O => \N__37264\,
            I => \N__37261\
        );

    \I__7062\ : Odrv4
    port map (
            O => \N__37261\,
            I => n2688
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__37258\,
            I => \n2720_cascade_\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__37255\,
            I => \n14038_cascade_\
        );

    \I__7059\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37249\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__37249\,
            I => n14042
        );

    \I__7057\ : InMux
    port map (
            O => \N__37246\,
            I => \N__37241\
        );

    \I__7056\ : InMux
    port map (
            O => \N__37245\,
            I => \N__37238\
        );

    \I__7055\ : InMux
    port map (
            O => \N__37244\,
            I => \N__37235\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__37241\,
            I => \N__37232\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__37238\,
            I => \N__37229\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37226\
        );

    \I__7051\ : Span4Mux_h
    port map (
            O => \N__37232\,
            I => \N__37223\
        );

    \I__7050\ : Span4Mux_h
    port map (
            O => \N__37229\,
            I => \N__37218\
        );

    \I__7049\ : Span4Mux_h
    port map (
            O => \N__37226\,
            I => \N__37218\
        );

    \I__7048\ : Odrv4
    port map (
            O => \N__37223\,
            I => n2614
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__37218\,
            I => n2614
        );

    \I__7046\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37210\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__37210\,
            I => \N__37207\
        );

    \I__7044\ : Span4Mux_h
    port map (
            O => \N__37207\,
            I => \N__37204\
        );

    \I__7043\ : Odrv4
    port map (
            O => \N__37204\,
            I => n2681
        );

    \I__7042\ : InMux
    port map (
            O => \N__37201\,
            I => \N__37198\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__37198\,
            I => \N__37195\
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__37195\,
            I => n2685
        );

    \I__7039\ : CascadeMux
    port map (
            O => \N__37192\,
            I => \N__37187\
        );

    \I__7038\ : InMux
    port map (
            O => \N__37191\,
            I => \N__37184\
        );

    \I__7037\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37181\
        );

    \I__7036\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37178\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__37184\,
            I => \N__37175\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__37181\,
            I => \N__37172\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__37178\,
            I => \N__37169\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__37175\,
            I => \N__37164\
        );

    \I__7031\ : Span4Mux_h
    port map (
            O => \N__37172\,
            I => \N__37164\
        );

    \I__7030\ : Odrv4
    port map (
            O => \N__37169\,
            I => n2618
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__37164\,
            I => n2618
        );

    \I__7028\ : InMux
    port map (
            O => \N__37159\,
            I => \N__37156\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__37156\,
            I => n14294
        );

    \I__7026\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37150\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__37150\,
            I => \N__37147\
        );

    \I__7024\ : Odrv4
    port map (
            O => \N__37147\,
            I => n2693
        );

    \I__7023\ : InMux
    port map (
            O => \N__37144\,
            I => \N__37140\
        );

    \I__7022\ : InMux
    port map (
            O => \N__37143\,
            I => \N__37137\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__37140\,
            I => \N__37134\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__37137\,
            I => n2626
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__37134\,
            I => n2626
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__37129\,
            I => \n2725_cascade_\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__37126\,
            I => \n14040_cascade_\
        );

    \I__7016\ : CascadeMux
    port map (
            O => \N__37123\,
            I => \N__37119\
        );

    \I__7015\ : InMux
    port map (
            O => \N__37122\,
            I => \N__37115\
        );

    \I__7014\ : InMux
    port map (
            O => \N__37119\,
            I => \N__37112\
        );

    \I__7013\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37109\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__37115\,
            I => n2629
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__37112\,
            I => n2629
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__37109\,
            I => n2629
        );

    \I__7009\ : CascadeMux
    port map (
            O => \N__37102\,
            I => \N__37099\
        );

    \I__7008\ : InMux
    port map (
            O => \N__37099\,
            I => \N__37096\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__37096\,
            I => \N__37093\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__37093\,
            I => n2696
        );

    \I__7005\ : CascadeMux
    port map (
            O => \N__37090\,
            I => \N__37087\
        );

    \I__7004\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37083\
        );

    \I__7003\ : InMux
    port map (
            O => \N__37086\,
            I => \N__37080\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__37083\,
            I => \N__37077\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__37080\,
            I => n2630
        );

    \I__7000\ : Odrv4
    port map (
            O => \N__37077\,
            I => n2630
        );

    \I__6999\ : InMux
    port map (
            O => \N__37072\,
            I => \N__37069\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__37069\,
            I => \N__37066\
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__37066\,
            I => n2697
        );

    \I__6996\ : InMux
    port map (
            O => \N__37063\,
            I => \N__37060\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__37060\,
            I => \N__37057\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__37057\,
            I => n2695
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__37054\,
            I => \N__37050\
        );

    \I__6992\ : CascadeMux
    port map (
            O => \N__37053\,
            I => \N__37047\
        );

    \I__6991\ : InMux
    port map (
            O => \N__37050\,
            I => \N__37044\
        );

    \I__6990\ : InMux
    port map (
            O => \N__37047\,
            I => \N__37041\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__37044\,
            I => \N__37038\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__37041\,
            I => \N__37035\
        );

    \I__6987\ : Span4Mux_h
    port map (
            O => \N__37038\,
            I => \N__37032\
        );

    \I__6986\ : Odrv12
    port map (
            O => \N__37035\,
            I => n2628
        );

    \I__6985\ : Odrv4
    port map (
            O => \N__37032\,
            I => n2628
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__37027\,
            I => \N__37023\
        );

    \I__6983\ : InMux
    port map (
            O => \N__37026\,
            I => \N__37020\
        );

    \I__6982\ : InMux
    port map (
            O => \N__37023\,
            I => \N__37016\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__37020\,
            I => \N__37013\
        );

    \I__6980\ : InMux
    port map (
            O => \N__37019\,
            I => \N__37010\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__37016\,
            I => n2619
        );

    \I__6978\ : Odrv4
    port map (
            O => \N__37013\,
            I => n2619
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__37010\,
            I => n2619
        );

    \I__6976\ : InMux
    port map (
            O => \N__37003\,
            I => \N__37000\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__37000\,
            I => \N__36997\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__36997\,
            I => \N__36994\
        );

    \I__6973\ : Odrv4
    port map (
            O => \N__36994\,
            I => n2686
        );

    \I__6972\ : InMux
    port map (
            O => \N__36991\,
            I => \N__36988\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__36988\,
            I => encoder0_position_scaled_23
        );

    \I__6970\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36982\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__36982\,
            I => \N__36979\
        );

    \I__6968\ : Span4Mux_h
    port map (
            O => \N__36979\,
            I => \N__36976\
        );

    \I__6967\ : Span4Mux_h
    port map (
            O => \N__36976\,
            I => \N__36973\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__36973\,
            I => \ENCODER0_A_N\
        );

    \I__6965\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36967\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__36967\,
            I => \N__36963\
        );

    \I__6963\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36960\
        );

    \I__6962\ : Span4Mux_v
    port map (
            O => \N__36963\,
            I => \N__36952\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__36960\,
            I => \N__36952\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__36959\,
            I => \N__36945\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__36958\,
            I => \N__36942\
        );

    \I__6958\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36938\
        );

    \I__6957\ : Span4Mux_h
    port map (
            O => \N__36952\,
            I => \N__36935\
        );

    \I__6956\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36932\
        );

    \I__6955\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36925\
        );

    \I__6954\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36925\
        );

    \I__6953\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36925\
        );

    \I__6952\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36918\
        );

    \I__6951\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36918\
        );

    \I__6950\ : InMux
    port map (
            O => \N__36941\,
            I => \N__36918\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__36938\,
            I => \N__36915\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__36935\,
            I => n1059
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__36932\,
            I => n1059
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__36925\,
            I => n1059
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__36918\,
            I => n1059
        );

    \I__6944\ : Odrv4
    port map (
            O => \N__36915\,
            I => n1059
        );

    \I__6943\ : InMux
    port map (
            O => \N__36904\,
            I => \N__36901\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__36901\,
            I => \N__36898\
        );

    \I__6941\ : Span4Mux_h
    port map (
            O => \N__36898\,
            I => \N__36895\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__36895\,
            I => n15210
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__36892\,
            I => \n14536_cascade_\
        );

    \I__6938\ : InMux
    port map (
            O => \N__36889\,
            I => \N__36886\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__36886\,
            I => \N__36883\
        );

    \I__6936\ : Span12Mux_v
    port map (
            O => \N__36883\,
            I => \N__36879\
        );

    \I__6935\ : InMux
    port map (
            O => \N__36882\,
            I => \N__36876\
        );

    \I__6934\ : Odrv12
    port map (
            O => \N__36879\,
            I => blink_counter_25
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__36876\,
            I => blink_counter_25
        );

    \I__6932\ : IoInMux
    port map (
            O => \N__36871\,
            I => \N__36868\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36865\
        );

    \I__6930\ : Span4Mux_s2_v
    port map (
            O => \N__36865\,
            I => \N__36862\
        );

    \I__6929\ : Span4Mux_h
    port map (
            O => \N__36862\,
            I => \N__36859\
        );

    \I__6928\ : Odrv4
    port map (
            O => \N__36859\,
            I => \LED_c\
        );

    \I__6927\ : InMux
    port map (
            O => \N__36856\,
            I => \N__36850\
        );

    \I__6926\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36850\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__36850\,
            I => \N__36847\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__36847\,
            I => \N__36844\
        );

    \I__6923\ : Span4Mux_h
    port map (
            O => \N__36844\,
            I => \N__36840\
        );

    \I__6922\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36837\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__36840\,
            I => blink_counter_24
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__36837\,
            I => blink_counter_24
        );

    \I__6919\ : InMux
    port map (
            O => \N__36832\,
            I => \N__36826\
        );

    \I__6918\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36826\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__36826\,
            I => \N__36822\
        );

    \I__6916\ : InMux
    port map (
            O => \N__36825\,
            I => \N__36819\
        );

    \I__6915\ : Odrv12
    port map (
            O => \N__36822\,
            I => blink_counter_21
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__36819\,
            I => blink_counter_21
        );

    \I__6913\ : CascadeMux
    port map (
            O => \N__36814\,
            I => \N__36810\
        );

    \I__6912\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36805\
        );

    \I__6911\ : InMux
    port map (
            O => \N__36810\,
            I => \N__36805\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__36805\,
            I => \N__36801\
        );

    \I__6909\ : InMux
    port map (
            O => \N__36804\,
            I => \N__36798\
        );

    \I__6908\ : Odrv12
    port map (
            O => \N__36801\,
            I => blink_counter_22
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__36798\,
            I => blink_counter_22
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__36793\,
            I => \N__36790\
        );

    \I__6905\ : InMux
    port map (
            O => \N__36790\,
            I => \N__36784\
        );

    \I__6904\ : InMux
    port map (
            O => \N__36789\,
            I => \N__36784\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__36784\,
            I => \N__36780\
        );

    \I__6902\ : InMux
    port map (
            O => \N__36783\,
            I => \N__36777\
        );

    \I__6901\ : Odrv12
    port map (
            O => \N__36780\,
            I => blink_counter_23
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__36777\,
            I => blink_counter_23
        );

    \I__6899\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36769\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__36769\,
            I => n14535
        );

    \I__6897\ : InMux
    port map (
            O => \N__36766\,
            I => \N__36763\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__36763\,
            I => \N__36760\
        );

    \I__6895\ : Span4Mux_v
    port map (
            O => \N__36760\,
            I => \N__36757\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__36757\,
            I => \N__36753\
        );

    \I__6893\ : InMux
    port map (
            O => \N__36756\,
            I => \N__36750\
        );

    \I__6892\ : Odrv4
    port map (
            O => \N__36753\,
            I => n15259
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__36750\,
            I => n15259
        );

    \I__6890\ : InMux
    port map (
            O => \N__36745\,
            I => \N__36740\
        );

    \I__6889\ : InMux
    port map (
            O => \N__36744\,
            I => \N__36734\
        );

    \I__6888\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36734\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__36740\,
            I => \N__36729\
        );

    \I__6886\ : CascadeMux
    port map (
            O => \N__36739\,
            I => \N__36726\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__36734\,
            I => \N__36722\
        );

    \I__6884\ : CascadeMux
    port map (
            O => \N__36733\,
            I => \N__36716\
        );

    \I__6883\ : CascadeMux
    port map (
            O => \N__36732\,
            I => \N__36712\
        );

    \I__6882\ : Span12Mux_v
    port map (
            O => \N__36729\,
            I => \N__36708\
        );

    \I__6881\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36703\
        );

    \I__6880\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36703\
        );

    \I__6879\ : Span4Mux_s3_h
    port map (
            O => \N__36722\,
            I => \N__36700\
        );

    \I__6878\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36695\
        );

    \I__6877\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36695\
        );

    \I__6876\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36684\
        );

    \I__6875\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36684\
        );

    \I__6874\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36684\
        );

    \I__6873\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36684\
        );

    \I__6872\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36684\
        );

    \I__6871\ : Odrv12
    port map (
            O => \N__36708\,
            I => n1356
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__36703\,
            I => n1356
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__36700\,
            I => n1356
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__36695\,
            I => n1356
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__36684\,
            I => n1356
        );

    \I__6866\ : InMux
    port map (
            O => \N__36673\,
            I => n12571
        );

    \I__6865\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36667\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__36667\,
            I => \N__36664\
        );

    \I__6863\ : Span4Mux_v
    port map (
            O => \N__36664\,
            I => \N__36660\
        );

    \I__6862\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36657\
        );

    \I__6861\ : Span4Mux_h
    port map (
            O => \N__36660\,
            I => \N__36654\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__36657\,
            I => \N__36651\
        );

    \I__6859\ : Odrv4
    port map (
            O => \N__36654\,
            I => n15243
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__36651\,
            I => n15243
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__36646\,
            I => \N__36643\
        );

    \I__6856\ : InMux
    port map (
            O => \N__36643\,
            I => \N__36640\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__36640\,
            I => \N__36637\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__36637\,
            I => \N__36632\
        );

    \I__6853\ : CascadeMux
    port map (
            O => \N__36636\,
            I => \N__36622\
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__36635\,
            I => \N__36619\
        );

    \I__6851\ : Span4Mux_h
    port map (
            O => \N__36632\,
            I => \N__36615\
        );

    \I__6850\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36612\
        );

    \I__6849\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36609\
        );

    \I__6848\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36604\
        );

    \I__6847\ : InMux
    port map (
            O => \N__36628\,
            I => \N__36604\
        );

    \I__6846\ : InMux
    port map (
            O => \N__36627\,
            I => \N__36601\
        );

    \I__6845\ : InMux
    port map (
            O => \N__36626\,
            I => \N__36590\
        );

    \I__6844\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36590\
        );

    \I__6843\ : InMux
    port map (
            O => \N__36622\,
            I => \N__36590\
        );

    \I__6842\ : InMux
    port map (
            O => \N__36619\,
            I => \N__36590\
        );

    \I__6841\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36590\
        );

    \I__6840\ : Odrv4
    port map (
            O => \N__36615\,
            I => n1257
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__36612\,
            I => n1257
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__36609\,
            I => n1257
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__36604\,
            I => n1257
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__36601\,
            I => n1257
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__36590\,
            I => n1257
        );

    \I__6834\ : InMux
    port map (
            O => \N__36577\,
            I => n12572
        );

    \I__6833\ : InMux
    port map (
            O => \N__36574\,
            I => \N__36571\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__36571\,
            I => \N__36567\
        );

    \I__6831\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36564\
        );

    \I__6830\ : Span4Mux_h
    port map (
            O => \N__36567\,
            I => \N__36561\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__36564\,
            I => \N__36558\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__36561\,
            I => \N__36553\
        );

    \I__6827\ : Span4Mux_s1_v
    port map (
            O => \N__36558\,
            I => \N__36553\
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__36553\,
            I => n15224
        );

    \I__6825\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36547\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__36547\,
            I => \N__36542\
        );

    \I__6823\ : CascadeMux
    port map (
            O => \N__36546\,
            I => \N__36533\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__36545\,
            I => \N__36530\
        );

    \I__6821\ : Span12Mux_v
    port map (
            O => \N__36542\,
            I => \N__36526\
        );

    \I__6820\ : InMux
    port map (
            O => \N__36541\,
            I => \N__36523\
        );

    \I__6819\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36520\
        );

    \I__6818\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36515\
        );

    \I__6817\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36515\
        );

    \I__6816\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36512\
        );

    \I__6815\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36503\
        );

    \I__6814\ : InMux
    port map (
            O => \N__36533\,
            I => \N__36503\
        );

    \I__6813\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36503\
        );

    \I__6812\ : InMux
    port map (
            O => \N__36529\,
            I => \N__36503\
        );

    \I__6811\ : Odrv12
    port map (
            O => \N__36526\,
            I => n1158
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__36523\,
            I => n1158
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__36520\,
            I => n1158
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__36515\,
            I => n1158
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__36512\,
            I => n1158
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__36503\,
            I => n1158
        );

    \I__6805\ : InMux
    port map (
            O => \N__36490\,
            I => n12573
        );

    \I__6804\ : CascadeMux
    port map (
            O => \N__36487\,
            I => \N__36466\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__36486\,
            I => \N__36463\
        );

    \I__6802\ : CascadeMux
    port map (
            O => \N__36485\,
            I => \N__36459\
        );

    \I__6801\ : CascadeMux
    port map (
            O => \N__36484\,
            I => \N__36455\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__36483\,
            I => \N__36451\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__36482\,
            I => \N__36448\
        );

    \I__6798\ : CascadeMux
    port map (
            O => \N__36481\,
            I => \N__36445\
        );

    \I__6797\ : CascadeMux
    port map (
            O => \N__36480\,
            I => \N__36442\
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__36479\,
            I => \N__36439\
        );

    \I__6795\ : CascadeMux
    port map (
            O => \N__36478\,
            I => \N__36435\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__36477\,
            I => \N__36432\
        );

    \I__6793\ : CascadeMux
    port map (
            O => \N__36476\,
            I => \N__36429\
        );

    \I__6792\ : CascadeMux
    port map (
            O => \N__36475\,
            I => \N__36426\
        );

    \I__6791\ : CascadeMux
    port map (
            O => \N__36474\,
            I => \N__36423\
        );

    \I__6790\ : CascadeMux
    port map (
            O => \N__36473\,
            I => \N__36420\
        );

    \I__6789\ : CascadeMux
    port map (
            O => \N__36472\,
            I => \N__36417\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__36471\,
            I => \N__36413\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__36470\,
            I => \N__36410\
        );

    \I__6786\ : CascadeMux
    port map (
            O => \N__36469\,
            I => \N__36407\
        );

    \I__6785\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36403\
        );

    \I__6784\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36388\
        );

    \I__6783\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36388\
        );

    \I__6782\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36388\
        );

    \I__6781\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36388\
        );

    \I__6780\ : InMux
    port map (
            O => \N__36455\,
            I => \N__36388\
        );

    \I__6779\ : InMux
    port map (
            O => \N__36454\,
            I => \N__36388\
        );

    \I__6778\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36388\
        );

    \I__6777\ : InMux
    port map (
            O => \N__36448\,
            I => \N__36379\
        );

    \I__6776\ : InMux
    port map (
            O => \N__36445\,
            I => \N__36379\
        );

    \I__6775\ : InMux
    port map (
            O => \N__36442\,
            I => \N__36379\
        );

    \I__6774\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36379\
        );

    \I__6773\ : CascadeMux
    port map (
            O => \N__36438\,
            I => \N__36376\
        );

    \I__6772\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36367\
        );

    \I__6771\ : InMux
    port map (
            O => \N__36432\,
            I => \N__36367\
        );

    \I__6770\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36367\
        );

    \I__6769\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36367\
        );

    \I__6768\ : InMux
    port map (
            O => \N__36423\,
            I => \N__36362\
        );

    \I__6767\ : InMux
    port map (
            O => \N__36420\,
            I => \N__36362\
        );

    \I__6766\ : InMux
    port map (
            O => \N__36417\,
            I => \N__36349\
        );

    \I__6765\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36349\
        );

    \I__6764\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36349\
        );

    \I__6763\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36349\
        );

    \I__6762\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36349\
        );

    \I__6761\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36349\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__36403\,
            I => \N__36342\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__36388\,
            I => \N__36342\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__36379\,
            I => \N__36342\
        );

    \I__6757\ : InMux
    port map (
            O => \N__36376\,
            I => \N__36339\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__36367\,
            I => \N__36332\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__36362\,
            I => \N__36332\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__36349\,
            I => \N__36332\
        );

    \I__6753\ : Span4Mux_v
    port map (
            O => \N__36342\,
            I => \N__36327\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__36339\,
            I => \N__36327\
        );

    \I__6751\ : Span4Mux_v
    port map (
            O => \N__36332\,
            I => \N__36324\
        );

    \I__6750\ : Span4Mux_h
    port map (
            O => \N__36327\,
            I => \N__36321\
        );

    \I__6749\ : Odrv4
    port map (
            O => \N__36324\,
            I => n2_adj_626
        );

    \I__6748\ : Odrv4
    port map (
            O => \N__36321\,
            I => n2_adj_626
        );

    \I__6747\ : InMux
    port map (
            O => \N__36316\,
            I => n12574
        );

    \I__6746\ : InMux
    port map (
            O => \N__36313\,
            I => \N__36310\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__36310\,
            I => encoder0_position_scaled_17
        );

    \I__6744\ : InMux
    port map (
            O => \N__36307\,
            I => \N__36304\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__36304\,
            I => encoder0_position_scaled_20
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__36301\,
            I => \N__36298\
        );

    \I__6741\ : InMux
    port map (
            O => \N__36298\,
            I => \N__36294\
        );

    \I__6740\ : CascadeMux
    port map (
            O => \N__36297\,
            I => \N__36291\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__36294\,
            I => \N__36288\
        );

    \I__6738\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36284\
        );

    \I__6737\ : Span4Mux_h
    port map (
            O => \N__36288\,
            I => \N__36281\
        );

    \I__6736\ : InMux
    port map (
            O => \N__36287\,
            I => \N__36278\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__36284\,
            I => encoder0_position_25
        );

    \I__6734\ : Odrv4
    port map (
            O => \N__36281\,
            I => encoder0_position_25
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__36278\,
            I => encoder0_position_25
        );

    \I__6732\ : InMux
    port map (
            O => \N__36271\,
            I => \N__36268\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__36268\,
            I => \N__36265\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__36265\,
            I => n8
        );

    \I__6729\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36255\
        );

    \I__6728\ : InMux
    port map (
            O => \N__36261\,
            I => \N__36255\
        );

    \I__6727\ : InMux
    port map (
            O => \N__36260\,
            I => \N__36252\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__36255\,
            I => \N__36249\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__36252\,
            I => \N__36246\
        );

    \I__6724\ : Span4Mux_v
    port map (
            O => \N__36249\,
            I => \N__36243\
        );

    \I__6723\ : Span4Mux_h
    port map (
            O => \N__36246\,
            I => \N__36240\
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__36243\,
            I => n294
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__36240\,
            I => n294
        );

    \I__6720\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36232\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__36232\,
            I => \N__36229\
        );

    \I__6718\ : Span4Mux_v
    port map (
            O => \N__36229\,
            I => \N__36226\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__36226\,
            I => \N__36223\
        );

    \I__6716\ : Span4Mux_h
    port map (
            O => \N__36223\,
            I => \N__36219\
        );

    \I__6715\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36216\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__36219\,
            I => n15059
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__36216\,
            I => n15059
        );

    \I__6712\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36208\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__36208\,
            I => \N__36202\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__36207\,
            I => \N__36195\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__36206\,
            I => \N__36188\
        );

    \I__6708\ : InMux
    port map (
            O => \N__36205\,
            I => \N__36185\
        );

    \I__6707\ : Span4Mux_v
    port map (
            O => \N__36202\,
            I => \N__36182\
        );

    \I__6706\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36177\
        );

    \I__6705\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36177\
        );

    \I__6704\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36174\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__36198\,
            I => \N__36170\
        );

    \I__6702\ : InMux
    port map (
            O => \N__36195\,
            I => \N__36163\
        );

    \I__6701\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36163\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__36193\,
            I => \N__36160\
        );

    \I__6699\ : CascadeMux
    port map (
            O => \N__36192\,
            I => \N__36154\
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__36191\,
            I => \N__36151\
        );

    \I__6697\ : InMux
    port map (
            O => \N__36188\,
            I => \N__36146\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__36185\,
            I => \N__36143\
        );

    \I__6695\ : Span4Mux_h
    port map (
            O => \N__36182\,
            I => \N__36136\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36136\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__36174\,
            I => \N__36136\
        );

    \I__6692\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36129\
        );

    \I__6691\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36129\
        );

    \I__6690\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36129\
        );

    \I__6689\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36126\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36123\
        );

    \I__6687\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36118\
        );

    \I__6686\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36118\
        );

    \I__6685\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36113\
        );

    \I__6684\ : InMux
    port map (
            O => \N__36157\,
            I => \N__36113\
        );

    \I__6683\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36104\
        );

    \I__6682\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36104\
        );

    \I__6681\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36104\
        );

    \I__6680\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36104\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__36146\,
            I => \N__36097\
        );

    \I__6678\ : Span4Mux_v
    port map (
            O => \N__36143\,
            I => \N__36097\
        );

    \I__6677\ : Span4Mux_v
    port map (
            O => \N__36136\,
            I => \N__36097\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__36129\,
            I => \N__36094\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__36126\,
            I => \N__36089\
        );

    \I__6674\ : Span4Mux_h
    port map (
            O => \N__36123\,
            I => \N__36089\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__36118\,
            I => n2148
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__36113\,
            I => n2148
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__36104\,
            I => n2148
        );

    \I__6670\ : Odrv4
    port map (
            O => \N__36097\,
            I => n2148
        );

    \I__6669\ : Odrv12
    port map (
            O => \N__36094\,
            I => n2148
        );

    \I__6668\ : Odrv4
    port map (
            O => \N__36089\,
            I => n2148
        );

    \I__6667\ : InMux
    port map (
            O => \N__36076\,
            I => n12563
        );

    \I__6666\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36069\
        );

    \I__6665\ : CascadeMux
    port map (
            O => \N__36072\,
            I => \N__36066\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__36069\,
            I => \N__36063\
        );

    \I__6663\ : InMux
    port map (
            O => \N__36066\,
            I => \N__36060\
        );

    \I__6662\ : Span12Mux_h
    port map (
            O => \N__36063\,
            I => \N__36057\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__36060\,
            I => \N__36054\
        );

    \I__6660\ : Odrv12
    port map (
            O => \N__36057\,
            I => n15035
        );

    \I__6659\ : Odrv4
    port map (
            O => \N__36054\,
            I => n15035
        );

    \I__6658\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36046\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36041\
        );

    \I__6656\ : CascadeMux
    port map (
            O => \N__36045\,
            I => \N__36038\
        );

    \I__6655\ : InMux
    port map (
            O => \N__36044\,
            I => \N__36033\
        );

    \I__6654\ : Span4Mux_v
    port map (
            O => \N__36041\,
            I => \N__36028\
        );

    \I__6653\ : InMux
    port map (
            O => \N__36038\,
            I => \N__36025\
        );

    \I__6652\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36022\
        );

    \I__6651\ : InMux
    port map (
            O => \N__36036\,
            I => \N__36019\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__36033\,
            I => \N__36012\
        );

    \I__6649\ : InMux
    port map (
            O => \N__36032\,
            I => \N__36007\
        );

    \I__6648\ : InMux
    port map (
            O => \N__36031\,
            I => \N__36007\
        );

    \I__6647\ : Span4Mux_h
    port map (
            O => \N__36028\,
            I => \N__35998\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__36025\,
            I => \N__35998\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__36022\,
            I => \N__35998\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__36019\,
            I => \N__35998\
        );

    \I__6643\ : InMux
    port map (
            O => \N__36018\,
            I => \N__35995\
        );

    \I__6642\ : CascadeMux
    port map (
            O => \N__36017\,
            I => \N__35988\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__36016\,
            I => \N__35982\
        );

    \I__6640\ : CascadeMux
    port map (
            O => \N__36015\,
            I => \N__35979\
        );

    \I__6639\ : Span4Mux_h
    port map (
            O => \N__36012\,
            I => \N__35969\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__36007\,
            I => \N__35969\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__35998\,
            I => \N__35969\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__35995\,
            I => \N__35969\
        );

    \I__6635\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35966\
        );

    \I__6634\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35963\
        );

    \I__6633\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35960\
        );

    \I__6632\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35957\
        );

    \I__6631\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35950\
        );

    \I__6630\ : InMux
    port map (
            O => \N__35987\,
            I => \N__35950\
        );

    \I__6629\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35950\
        );

    \I__6628\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35941\
        );

    \I__6627\ : InMux
    port map (
            O => \N__35982\,
            I => \N__35941\
        );

    \I__6626\ : InMux
    port map (
            O => \N__35979\,
            I => \N__35941\
        );

    \I__6625\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35941\
        );

    \I__6624\ : Span4Mux_h
    port map (
            O => \N__35969\,
            I => \N__35938\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__35966\,
            I => n2049
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__35963\,
            I => n2049
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__35960\,
            I => n2049
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__35957\,
            I => n2049
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__35950\,
            I => n2049
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__35941\,
            I => n2049
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__35938\,
            I => n2049
        );

    \I__6616\ : InMux
    port map (
            O => \N__35923\,
            I => n12564
        );

    \I__6615\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35917\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__35917\,
            I => \N__35914\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__35914\,
            I => \N__35911\
        );

    \I__6612\ : Span4Mux_h
    port map (
            O => \N__35911\,
            I => \N__35907\
        );

    \I__6611\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35904\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__35907\,
            I => n15012
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__35904\,
            I => n15012
        );

    \I__6608\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35896\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35891\
        );

    \I__6606\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35885\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__35894\,
            I => \N__35882\
        );

    \I__6604\ : Span4Mux_h
    port map (
            O => \N__35891\,
            I => \N__35879\
        );

    \I__6603\ : CascadeMux
    port map (
            O => \N__35890\,
            I => \N__35876\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__35889\,
            I => \N__35864\
        );

    \I__6601\ : CascadeMux
    port map (
            O => \N__35888\,
            I => \N__35859\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__35885\,
            I => \N__35855\
        );

    \I__6599\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35852\
        );

    \I__6598\ : Span4Mux_v
    port map (
            O => \N__35879\,
            I => \N__35849\
        );

    \I__6597\ : InMux
    port map (
            O => \N__35876\,
            I => \N__35846\
        );

    \I__6596\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35843\
        );

    \I__6595\ : InMux
    port map (
            O => \N__35874\,
            I => \N__35838\
        );

    \I__6594\ : InMux
    port map (
            O => \N__35873\,
            I => \N__35838\
        );

    \I__6593\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35835\
        );

    \I__6592\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35832\
        );

    \I__6591\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35825\
        );

    \I__6590\ : InMux
    port map (
            O => \N__35869\,
            I => \N__35825\
        );

    \I__6589\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35825\
        );

    \I__6588\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35812\
        );

    \I__6587\ : InMux
    port map (
            O => \N__35864\,
            I => \N__35812\
        );

    \I__6586\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35812\
        );

    \I__6585\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35812\
        );

    \I__6584\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35812\
        );

    \I__6583\ : InMux
    port map (
            O => \N__35858\,
            I => \N__35812\
        );

    \I__6582\ : Span4Mux_s3_h
    port map (
            O => \N__35855\,
            I => \N__35807\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__35852\,
            I => \N__35807\
        );

    \I__6580\ : Odrv4
    port map (
            O => \N__35849\,
            I => n1950
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__35846\,
            I => n1950
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__35843\,
            I => n1950
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__35838\,
            I => n1950
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__35835\,
            I => n1950
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__35832\,
            I => n1950
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__35825\,
            I => n1950
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__35812\,
            I => n1950
        );

    \I__6572\ : Odrv4
    port map (
            O => \N__35807\,
            I => n1950
        );

    \I__6571\ : InMux
    port map (
            O => \N__35788\,
            I => n12565
        );

    \I__6570\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35782\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__35782\,
            I => \N__35779\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__35779\,
            I => \N__35776\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__35776\,
            I => \N__35773\
        );

    \I__6566\ : Odrv4
    port map (
            O => \N__35773\,
            I => n14990
        );

    \I__6565\ : InMux
    port map (
            O => \N__35770\,
            I => \N__35767\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__35767\,
            I => \N__35762\
        );

    \I__6563\ : InMux
    port map (
            O => \N__35766\,
            I => \N__35758\
        );

    \I__6562\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35755\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__35762\,
            I => \N__35748\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__35761\,
            I => \N__35744\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35741\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35738\
        );

    \I__6557\ : CascadeMux
    port map (
            O => \N__35754\,
            I => \N__35734\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__35753\,
            I => \N__35730\
        );

    \I__6555\ : CascadeMux
    port map (
            O => \N__35752\,
            I => \N__35722\
        );

    \I__6554\ : InMux
    port map (
            O => \N__35751\,
            I => \N__35717\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__35748\,
            I => \N__35714\
        );

    \I__6552\ : InMux
    port map (
            O => \N__35747\,
            I => \N__35711\
        );

    \I__6551\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35708\
        );

    \I__6550\ : Span4Mux_s3_h
    port map (
            O => \N__35741\,
            I => \N__35705\
        );

    \I__6549\ : Span4Mux_s3_h
    port map (
            O => \N__35738\,
            I => \N__35702\
        );

    \I__6548\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35689\
        );

    \I__6547\ : InMux
    port map (
            O => \N__35734\,
            I => \N__35689\
        );

    \I__6546\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35689\
        );

    \I__6545\ : InMux
    port map (
            O => \N__35730\,
            I => \N__35689\
        );

    \I__6544\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35689\
        );

    \I__6543\ : InMux
    port map (
            O => \N__35728\,
            I => \N__35689\
        );

    \I__6542\ : InMux
    port map (
            O => \N__35727\,
            I => \N__35680\
        );

    \I__6541\ : InMux
    port map (
            O => \N__35726\,
            I => \N__35680\
        );

    \I__6540\ : InMux
    port map (
            O => \N__35725\,
            I => \N__35680\
        );

    \I__6539\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35680\
        );

    \I__6538\ : InMux
    port map (
            O => \N__35721\,
            I => \N__35675\
        );

    \I__6537\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35675\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__35717\,
            I => n1851
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__35714\,
            I => n1851
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__35711\,
            I => n1851
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__35708\,
            I => n1851
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__35705\,
            I => n1851
        );

    \I__6531\ : Odrv4
    port map (
            O => \N__35702\,
            I => n1851
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__35689\,
            I => n1851
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__35680\,
            I => n1851
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__35675\,
            I => n1851
        );

    \I__6527\ : InMux
    port map (
            O => \N__35656\,
            I => n12566
        );

    \I__6526\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35650\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__35650\,
            I => \N__35647\
        );

    \I__6524\ : Span4Mux_v
    port map (
            O => \N__35647\,
            I => \N__35643\
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__35646\,
            I => \N__35640\
        );

    \I__6522\ : Span4Mux_h
    port map (
            O => \N__35643\,
            I => \N__35637\
        );

    \I__6521\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35634\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__35637\,
            I => n14969
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__35634\,
            I => n14969
        );

    \I__6518\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35625\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__35628\,
            I => \N__35616\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__35625\,
            I => \N__35612\
        );

    \I__6515\ : CascadeMux
    port map (
            O => \N__35624\,
            I => \N__35608\
        );

    \I__6514\ : InMux
    port map (
            O => \N__35623\,
            I => \N__35604\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__35622\,
            I => \N__35601\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__35621\,
            I => \N__35596\
        );

    \I__6511\ : InMux
    port map (
            O => \N__35620\,
            I => \N__35585\
        );

    \I__6510\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35585\
        );

    \I__6509\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35585\
        );

    \I__6508\ : InMux
    port map (
            O => \N__35615\,
            I => \N__35585\
        );

    \I__6507\ : Span4Mux_v
    port map (
            O => \N__35612\,
            I => \N__35581\
        );

    \I__6506\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35574\
        );

    \I__6505\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35574\
        );

    \I__6504\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35574\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__35604\,
            I => \N__35571\
        );

    \I__6502\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35566\
        );

    \I__6501\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35566\
        );

    \I__6500\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35559\
        );

    \I__6499\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35559\
        );

    \I__6498\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35559\
        );

    \I__6497\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35556\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__35585\,
            I => \N__35553\
        );

    \I__6495\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35550\
        );

    \I__6494\ : Span4Mux_h
    port map (
            O => \N__35581\,
            I => \N__35543\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__35574\,
            I => \N__35543\
        );

    \I__6492\ : Span4Mux_v
    port map (
            O => \N__35571\,
            I => \N__35543\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__35566\,
            I => n1752
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__35559\,
            I => n1752
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__35556\,
            I => n1752
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__35553\,
            I => n1752
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__35550\,
            I => n1752
        );

    \I__6486\ : Odrv4
    port map (
            O => \N__35543\,
            I => n1752
        );

    \I__6485\ : InMux
    port map (
            O => \N__35530\,
            I => \bfn_9_27_0_\
        );

    \I__6484\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35524\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__35524\,
            I => \N__35521\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__35521\,
            I => \N__35517\
        );

    \I__6481\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35514\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__35517\,
            I => \N__35511\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__35514\,
            I => \N__35508\
        );

    \I__6478\ : Odrv4
    port map (
            O => \N__35511\,
            I => n14949
        );

    \I__6477\ : Odrv4
    port map (
            O => \N__35508\,
            I => n14949
        );

    \I__6476\ : CascadeMux
    port map (
            O => \N__35503\,
            I => \N__35500\
        );

    \I__6475\ : InMux
    port map (
            O => \N__35500\,
            I => \N__35497\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__35497\,
            I => \N__35494\
        );

    \I__6473\ : Span4Mux_h
    port map (
            O => \N__35494\,
            I => \N__35488\
        );

    \I__6472\ : CascadeMux
    port map (
            O => \N__35493\,
            I => \N__35477\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__35492\,
            I => \N__35473\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__35491\,
            I => \N__35470\
        );

    \I__6469\ : Span4Mux_h
    port map (
            O => \N__35488\,
            I => \N__35465\
        );

    \I__6468\ : InMux
    port map (
            O => \N__35487\,
            I => \N__35462\
        );

    \I__6467\ : InMux
    port map (
            O => \N__35486\,
            I => \N__35455\
        );

    \I__6466\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35455\
        );

    \I__6465\ : InMux
    port map (
            O => \N__35484\,
            I => \N__35455\
        );

    \I__6464\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35446\
        );

    \I__6463\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35446\
        );

    \I__6462\ : InMux
    port map (
            O => \N__35481\,
            I => \N__35446\
        );

    \I__6461\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35446\
        );

    \I__6460\ : InMux
    port map (
            O => \N__35477\,
            I => \N__35433\
        );

    \I__6459\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35433\
        );

    \I__6458\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35433\
        );

    \I__6457\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35433\
        );

    \I__6456\ : InMux
    port map (
            O => \N__35469\,
            I => \N__35433\
        );

    \I__6455\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35433\
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__35465\,
            I => n1653
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__35462\,
            I => n1653
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__35455\,
            I => n1653
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__35446\,
            I => n1653
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__35433\,
            I => n1653
        );

    \I__6449\ : InMux
    port map (
            O => \N__35422\,
            I => n12568
        );

    \I__6448\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35416\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__35416\,
            I => \N__35413\
        );

    \I__6446\ : Span4Mux_v
    port map (
            O => \N__35413\,
            I => \N__35410\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__35410\,
            I => \N__35406\
        );

    \I__6444\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35403\
        );

    \I__6443\ : Odrv4
    port map (
            O => \N__35406\,
            I => n15292
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__35403\,
            I => n15292
        );

    \I__6441\ : InMux
    port map (
            O => \N__35398\,
            I => \N__35395\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__35395\,
            I => \N__35392\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__35392\,
            I => \N__35385\
        );

    \I__6438\ : CascadeMux
    port map (
            O => \N__35391\,
            I => \N__35379\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__35390\,
            I => \N__35375\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__35389\,
            I => \N__35369\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__35388\,
            I => \N__35366\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__35385\,
            I => \N__35361\
        );

    \I__6433\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35356\
        );

    \I__6432\ : InMux
    port map (
            O => \N__35383\,
            I => \N__35356\
        );

    \I__6431\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35353\
        );

    \I__6430\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35342\
        );

    \I__6429\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35342\
        );

    \I__6428\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35342\
        );

    \I__6427\ : InMux
    port map (
            O => \N__35374\,
            I => \N__35342\
        );

    \I__6426\ : InMux
    port map (
            O => \N__35373\,
            I => \N__35342\
        );

    \I__6425\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35331\
        );

    \I__6424\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35331\
        );

    \I__6423\ : InMux
    port map (
            O => \N__35366\,
            I => \N__35331\
        );

    \I__6422\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35331\
        );

    \I__6421\ : InMux
    port map (
            O => \N__35364\,
            I => \N__35331\
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__35361\,
            I => n1554
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__35356\,
            I => n1554
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__35353\,
            I => n1554
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__35342\,
            I => n1554
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__35331\,
            I => n1554
        );

    \I__6415\ : InMux
    port map (
            O => \N__35320\,
            I => n12569
        );

    \I__6414\ : InMux
    port map (
            O => \N__35317\,
            I => \N__35314\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__35314\,
            I => \N__35311\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__35311\,
            I => \N__35307\
        );

    \I__6411\ : CascadeMux
    port map (
            O => \N__35310\,
            I => \N__35304\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__35307\,
            I => \N__35301\
        );

    \I__6409\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35298\
        );

    \I__6408\ : Odrv4
    port map (
            O => \N__35301\,
            I => n15276
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__35298\,
            I => n15276
        );

    \I__6406\ : CascadeMux
    port map (
            O => \N__35293\,
            I => \N__35290\
        );

    \I__6405\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35287\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__35287\,
            I => \N__35283\
        );

    \I__6403\ : CascadeMux
    port map (
            O => \N__35286\,
            I => \N__35276\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__35283\,
            I => \N__35271\
        );

    \I__6401\ : InMux
    port map (
            O => \N__35282\,
            I => \N__35268\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__35281\,
            I => \N__35265\
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__35280\,
            I => \N__35262\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__35279\,
            I => \N__35259\
        );

    \I__6397\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35251\
        );

    \I__6396\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35251\
        );

    \I__6395\ : CascadeMux
    port map (
            O => \N__35274\,
            I => \N__35248\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__35271\,
            I => \N__35243\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__35268\,
            I => \N__35240\
        );

    \I__6392\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35231\
        );

    \I__6391\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35231\
        );

    \I__6390\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35231\
        );

    \I__6389\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35231\
        );

    \I__6388\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35228\
        );

    \I__6387\ : InMux
    port map (
            O => \N__35256\,
            I => \N__35225\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__35251\,
            I => \N__35222\
        );

    \I__6385\ : InMux
    port map (
            O => \N__35248\,
            I => \N__35215\
        );

    \I__6384\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35215\
        );

    \I__6383\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35215\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__35243\,
            I => n1455
        );

    \I__6381\ : Odrv4
    port map (
            O => \N__35240\,
            I => n1455
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__35231\,
            I => n1455
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__35228\,
            I => n1455
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__35225\,
            I => n1455
        );

    \I__6377\ : Odrv4
    port map (
            O => \N__35222\,
            I => n1455
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__35215\,
            I => n1455
        );

    \I__6375\ : InMux
    port map (
            O => \N__35200\,
            I => n12570
        );

    \I__6374\ : InMux
    port map (
            O => \N__35197\,
            I => n12555
        );

    \I__6373\ : InMux
    port map (
            O => \N__35194\,
            I => n12556
        );

    \I__6372\ : InMux
    port map (
            O => \N__35191\,
            I => n12557
        );

    \I__6371\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35185\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__35185\,
            I => \N__35181\
        );

    \I__6369\ : CascadeMux
    port map (
            O => \N__35184\,
            I => \N__35178\
        );

    \I__6368\ : Span4Mux_v
    port map (
            O => \N__35181\,
            I => \N__35175\
        );

    \I__6367\ : InMux
    port map (
            O => \N__35178\,
            I => \N__35172\
        );

    \I__6366\ : Odrv4
    port map (
            O => \N__35175\,
            I => n15437
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__35172\,
            I => n15437
        );

    \I__6364\ : InMux
    port map (
            O => \N__35167\,
            I => n12558
        );

    \I__6363\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35161\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__35161\,
            I => \N__35158\
        );

    \I__6361\ : Sp12to4
    port map (
            O => \N__35158\,
            I => \N__35154\
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__35157\,
            I => \N__35151\
        );

    \I__6359\ : Span12Mux_v
    port map (
            O => \N__35154\,
            I => \N__35148\
        );

    \I__6358\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35145\
        );

    \I__6357\ : Odrv12
    port map (
            O => \N__35148\,
            I => n15401
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__35145\,
            I => n15401
        );

    \I__6355\ : InMux
    port map (
            O => \N__35140\,
            I => \bfn_9_26_0_\
        );

    \I__6354\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35134\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__35134\,
            I => \N__35130\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__35133\,
            I => \N__35127\
        );

    \I__6351\ : Span4Mux_h
    port map (
            O => \N__35130\,
            I => \N__35124\
        );

    \I__6350\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35121\
        );

    \I__6349\ : Sp12to4
    port map (
            O => \N__35124\,
            I => \N__35116\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__35116\
        );

    \I__6347\ : Odrv12
    port map (
            O => \N__35116\,
            I => n15375
        );

    \I__6346\ : InMux
    port map (
            O => \N__35113\,
            I => \N__35110\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__35110\,
            I => \N__35098\
        );

    \I__6344\ : CascadeMux
    port map (
            O => \N__35109\,
            I => \N__35094\
        );

    \I__6343\ : CascadeMux
    port map (
            O => \N__35108\,
            I => \N__35089\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__35107\,
            I => \N__35086\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__35106\,
            I => \N__35081\
        );

    \I__6340\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35076\
        );

    \I__6339\ : InMux
    port map (
            O => \N__35104\,
            I => \N__35076\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__35103\,
            I => \N__35071\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__35102\,
            I => \N__35068\
        );

    \I__6336\ : InMux
    port map (
            O => \N__35101\,
            I => \N__35064\
        );

    \I__6335\ : Span4Mux_v
    port map (
            O => \N__35098\,
            I => \N__35061\
        );

    \I__6334\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35054\
        );

    \I__6333\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35054\
        );

    \I__6332\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35054\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__35092\,
            I => \N__35049\
        );

    \I__6330\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35039\
        );

    \I__6329\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35039\
        );

    \I__6328\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35039\
        );

    \I__6327\ : InMux
    port map (
            O => \N__35084\,
            I => \N__35034\
        );

    \I__6326\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35034\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35031\
        );

    \I__6324\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35026\
        );

    \I__6323\ : InMux
    port map (
            O => \N__35074\,
            I => \N__35026\
        );

    \I__6322\ : InMux
    port map (
            O => \N__35071\,
            I => \N__35023\
        );

    \I__6321\ : InMux
    port map (
            O => \N__35068\,
            I => \N__35018\
        );

    \I__6320\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35018\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__35064\,
            I => \N__35015\
        );

    \I__6318\ : Span4Mux_v
    port map (
            O => \N__35061\,
            I => \N__35010\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__35054\,
            I => \N__35010\
        );

    \I__6316\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35007\
        );

    \I__6315\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35004\
        );

    \I__6314\ : InMux
    port map (
            O => \N__35049\,
            I => \N__34997\
        );

    \I__6313\ : InMux
    port map (
            O => \N__35048\,
            I => \N__34997\
        );

    \I__6312\ : InMux
    port map (
            O => \N__35047\,
            I => \N__34997\
        );

    \I__6311\ : InMux
    port map (
            O => \N__35046\,
            I => \N__34994\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__35039\,
            I => \N__34989\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__35034\,
            I => \N__34989\
        );

    \I__6308\ : Span4Mux_v
    port map (
            O => \N__35031\,
            I => \N__34978\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__35026\,
            I => \N__34978\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__35023\,
            I => \N__34978\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__35018\,
            I => \N__34978\
        );

    \I__6304\ : Span4Mux_h
    port map (
            O => \N__35015\,
            I => \N__34978\
        );

    \I__6303\ : Span4Mux_h
    port map (
            O => \N__35010\,
            I => \N__34975\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__35007\,
            I => n2445
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__35004\,
            I => n2445
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__34997\,
            I => n2445
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__34994\,
            I => n2445
        );

    \I__6298\ : Odrv4
    port map (
            O => \N__34989\,
            I => n2445
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__34978\,
            I => n2445
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__34975\,
            I => n2445
        );

    \I__6295\ : InMux
    port map (
            O => \N__34960\,
            I => n12560
        );

    \I__6294\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34954\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__34954\,
            I => \N__34951\
        );

    \I__6292\ : Span12Mux_h
    port map (
            O => \N__34951\,
            I => \N__34947\
        );

    \I__6291\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34944\
        );

    \I__6290\ : Odrv12
    port map (
            O => \N__34947\,
            I => n15348
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__34944\,
            I => n15348
        );

    \I__6288\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34936\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__34936\,
            I => \N__34932\
        );

    \I__6286\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34921\
        );

    \I__6285\ : Span4Mux_h
    port map (
            O => \N__34932\,
            I => \N__34916\
        );

    \I__6284\ : InMux
    port map (
            O => \N__34931\,
            I => \N__34913\
        );

    \I__6283\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34910\
        );

    \I__6282\ : InMux
    port map (
            O => \N__34929\,
            I => \N__34907\
        );

    \I__6281\ : CascadeMux
    port map (
            O => \N__34928\,
            I => \N__34901\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__34927\,
            I => \N__34897\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__34926\,
            I => \N__34891\
        );

    \I__6278\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34885\
        );

    \I__6277\ : InMux
    port map (
            O => \N__34924\,
            I => \N__34885\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__34921\,
            I => \N__34882\
        );

    \I__6275\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34877\
        );

    \I__6274\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34877\
        );

    \I__6273\ : Span4Mux_v
    port map (
            O => \N__34916\,
            I => \N__34872\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__34913\,
            I => \N__34872\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__34910\,
            I => \N__34869\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__34907\,
            I => \N__34866\
        );

    \I__6269\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34861\
        );

    \I__6268\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34852\
        );

    \I__6267\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34852\
        );

    \I__6266\ : InMux
    port map (
            O => \N__34901\,
            I => \N__34852\
        );

    \I__6265\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34852\
        );

    \I__6264\ : InMux
    port map (
            O => \N__34897\,
            I => \N__34847\
        );

    \I__6263\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34847\
        );

    \I__6262\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34838\
        );

    \I__6261\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34838\
        );

    \I__6260\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34838\
        );

    \I__6259\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34838\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__34885\,
            I => \N__34835\
        );

    \I__6257\ : Span4Mux_s3_h
    port map (
            O => \N__34882\,
            I => \N__34830\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__34877\,
            I => \N__34830\
        );

    \I__6255\ : Span4Mux_h
    port map (
            O => \N__34872\,
            I => \N__34823\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__34869\,
            I => \N__34823\
        );

    \I__6253\ : Span4Mux_s3_h
    port map (
            O => \N__34866\,
            I => \N__34823\
        );

    \I__6252\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34818\
        );

    \I__6251\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34818\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__34861\,
            I => n2346
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__34852\,
            I => n2346
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__34847\,
            I => n2346
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__34838\,
            I => n2346
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__34835\,
            I => n2346
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__34830\,
            I => n2346
        );

    \I__6244\ : Odrv4
    port map (
            O => \N__34823\,
            I => n2346
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__34818\,
            I => n2346
        );

    \I__6242\ : InMux
    port map (
            O => \N__34801\,
            I => n12561
        );

    \I__6241\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34795\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__34795\,
            I => \N__34791\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__34794\,
            I => \N__34788\
        );

    \I__6238\ : Span4Mux_v
    port map (
            O => \N__34791\,
            I => \N__34785\
        );

    \I__6237\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34782\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__34785\,
            I => n15322
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__34782\,
            I => n15322
        );

    \I__6234\ : InMux
    port map (
            O => \N__34777\,
            I => n12562
        );

    \I__6233\ : CascadeMux
    port map (
            O => \N__34774\,
            I => \n3138_cascade_\
        );

    \I__6232\ : CascadeMux
    port map (
            O => \N__34771\,
            I => \n3229_cascade_\
        );

    \I__6231\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34765\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__34765\,
            I => n11658
        );

    \I__6229\ : InMux
    port map (
            O => \N__34762\,
            I => \bfn_9_25_0_\
        );

    \I__6228\ : InMux
    port map (
            O => \N__34759\,
            I => n12552
        );

    \I__6227\ : InMux
    port map (
            O => \N__34756\,
            I => n12553
        );

    \I__6226\ : InMux
    port map (
            O => \N__34753\,
            I => n12554
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__34750\,
            I => \n11750_cascade_\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__34747\,
            I => \n13900_cascade_\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__34744\,
            I => \n3232_cascade_\
        );

    \I__6222\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34738\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__34738\,
            I => n13906
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__34735\,
            I => \n13912_cascade_\
        );

    \I__6219\ : InMux
    port map (
            O => \N__34732\,
            I => n12381
        );

    \I__6218\ : InMux
    port map (
            O => \N__34729\,
            I => n12382
        );

    \I__6217\ : InMux
    port map (
            O => \N__34726\,
            I => n12383
        );

    \I__6216\ : InMux
    port map (
            O => \N__34723\,
            I => n12384
        );

    \I__6215\ : InMux
    port map (
            O => \N__34720\,
            I => \bfn_9_22_0_\
        );

    \I__6214\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34712\
        );

    \I__6213\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34709\
        );

    \I__6212\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34706\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34699\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__34709\,
            I => \N__34699\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__34706\,
            I => \N__34699\
        );

    \I__6208\ : Span4Mux_v
    port map (
            O => \N__34699\,
            I => \N__34696\
        );

    \I__6207\ : Odrv4
    port map (
            O => \N__34696\,
            I => n2622
        );

    \I__6206\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34690\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__34690\,
            I => \N__34687\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__34687\,
            I => n2689
        );

    \I__6203\ : InMux
    port map (
            O => \N__34684\,
            I => n12373
        );

    \I__6202\ : InMux
    port map (
            O => \N__34681\,
            I => n12374
        );

    \I__6201\ : InMux
    port map (
            O => \N__34678\,
            I => n12375
        );

    \I__6200\ : InMux
    port map (
            O => \N__34675\,
            I => n12376
        );

    \I__6199\ : InMux
    port map (
            O => \N__34672\,
            I => \bfn_9_21_0_\
        );

    \I__6198\ : InMux
    port map (
            O => \N__34669\,
            I => n12378
        );

    \I__6197\ : InMux
    port map (
            O => \N__34666\,
            I => n12379
        );

    \I__6196\ : InMux
    port map (
            O => \N__34663\,
            I => n12380
        );

    \I__6195\ : InMux
    port map (
            O => \N__34660\,
            I => n12364
        );

    \I__6194\ : InMux
    port map (
            O => \N__34657\,
            I => n12365
        );

    \I__6193\ : InMux
    port map (
            O => \N__34654\,
            I => n12366
        );

    \I__6192\ : InMux
    port map (
            O => \N__34651\,
            I => n12367
        );

    \I__6191\ : InMux
    port map (
            O => \N__34648\,
            I => n12368
        );

    \I__6190\ : InMux
    port map (
            O => \N__34645\,
            I => \bfn_9_20_0_\
        );

    \I__6189\ : InMux
    port map (
            O => \N__34642\,
            I => \N__34639\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__34639\,
            I => \N__34635\
        );

    \I__6187\ : InMux
    port map (
            O => \N__34638\,
            I => \N__34632\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__34635\,
            I => n2625
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__34632\,
            I => n2625
        );

    \I__6184\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34624\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__34624\,
            I => \N__34621\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__34621\,
            I => n2692
        );

    \I__6181\ : InMux
    port map (
            O => \N__34618\,
            I => n12370
        );

    \I__6180\ : InMux
    port map (
            O => \N__34615\,
            I => n12371
        );

    \I__6179\ : InMux
    port map (
            O => \N__34612\,
            I => n12372
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__34609\,
            I => \N__34605\
        );

    \I__6177\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34602\
        );

    \I__6176\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34599\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__34602\,
            I => \N__34595\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__34599\,
            I => \N__34592\
        );

    \I__6173\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34589\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__34595\,
            I => \N__34586\
        );

    \I__6171\ : Span4Mux_v
    port map (
            O => \N__34592\,
            I => \N__34581\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34581\
        );

    \I__6169\ : Odrv4
    port map (
            O => \N__34586\,
            I => n2520
        );

    \I__6168\ : Odrv4
    port map (
            O => \N__34581\,
            I => n2520
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__34576\,
            I => \N__34573\
        );

    \I__6166\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__6164\ : Span4Mux_h
    port map (
            O => \N__34567\,
            I => \N__34564\
        );

    \I__6163\ : Odrv4
    port map (
            O => \N__34564\,
            I => n2587
        );

    \I__6162\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34558\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34555\
        );

    \I__6160\ : Span4Mux_h
    port map (
            O => \N__34555\,
            I => \N__34552\
        );

    \I__6159\ : Odrv4
    port map (
            O => \N__34552\,
            I => n2580
        );

    \I__6158\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34544\
        );

    \I__6157\ : InMux
    port map (
            O => \N__34548\,
            I => \N__34541\
        );

    \I__6156\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34538\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34533\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34533\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34530\
        );

    \I__6152\ : Span4Mux_h
    port map (
            O => \N__34533\,
            I => \N__34527\
        );

    \I__6151\ : Odrv12
    port map (
            O => \N__34530\,
            I => n2513
        );

    \I__6150\ : Odrv4
    port map (
            O => \N__34527\,
            I => n2513
        );

    \I__6149\ : CascadeMux
    port map (
            O => \N__34522\,
            I => \n2721_cascade_\
        );

    \I__6148\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34515\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__34518\,
            I => \N__34512\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34508\
        );

    \I__6145\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34505\
        );

    \I__6144\ : CascadeMux
    port map (
            O => \N__34511\,
            I => \N__34502\
        );

    \I__6143\ : Span4Mux_h
    port map (
            O => \N__34508\,
            I => \N__34497\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34497\
        );

    \I__6141\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34494\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__34497\,
            I => n2526
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__34494\,
            I => n2526
        );

    \I__6138\ : CascadeMux
    port map (
            O => \N__34489\,
            I => \N__34486\
        );

    \I__6137\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34483\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34480\
        );

    \I__6135\ : Span4Mux_v
    port map (
            O => \N__34480\,
            I => \N__34477\
        );

    \I__6134\ : Odrv4
    port map (
            O => \N__34477\,
            I => n2593
        );

    \I__6133\ : CascadeMux
    port map (
            O => \N__34474\,
            I => \n2625_cascade_\
        );

    \I__6132\ : InMux
    port map (
            O => \N__34471\,
            I => \bfn_9_19_0_\
        );

    \I__6131\ : InMux
    port map (
            O => \N__34468\,
            I => n12362
        );

    \I__6130\ : InMux
    port map (
            O => \N__34465\,
            I => n12363
        );

    \I__6129\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34458\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__34461\,
            I => \N__34455\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__34458\,
            I => \N__34452\
        );

    \I__6126\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34449\
        );

    \I__6125\ : Span4Mux_h
    port map (
            O => \N__34452\,
            I => \N__34444\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__34449\,
            I => \N__34444\
        );

    \I__6123\ : Sp12to4
    port map (
            O => \N__34444\,
            I => \N__34440\
        );

    \I__6122\ : InMux
    port map (
            O => \N__34443\,
            I => \N__34437\
        );

    \I__6121\ : Odrv12
    port map (
            O => \N__34440\,
            I => n2531
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__34437\,
            I => n2531
        );

    \I__6119\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34429\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__34429\,
            I => \N__34426\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__34426\,
            I => \N__34423\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__34423\,
            I => n2598
        );

    \I__6115\ : CascadeMux
    port map (
            O => \N__34420\,
            I => \n2630_cascade_\
        );

    \I__6114\ : CascadeMux
    port map (
            O => \N__34417\,
            I => \n14288_cascade_\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__34414\,
            I => \N__34410\
        );

    \I__6112\ : InMux
    port map (
            O => \N__34413\,
            I => \N__34407\
        );

    \I__6111\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34404\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__34407\,
            I => \N__34401\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__34404\,
            I => \N__34398\
        );

    \I__6108\ : Odrv12
    port map (
            O => \N__34401\,
            I => n2527
        );

    \I__6107\ : Odrv4
    port map (
            O => \N__34398\,
            I => n2527
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__34393\,
            I => \N__34390\
        );

    \I__6105\ : InMux
    port map (
            O => \N__34390\,
            I => \N__34387\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34384\
        );

    \I__6103\ : Span4Mux_v
    port map (
            O => \N__34384\,
            I => \N__34381\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__34381\,
            I => n2594
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__34378\,
            I => \n2626_cascade_\
        );

    \I__6100\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34372\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__34372\,
            I => \N__34369\
        );

    \I__6098\ : Odrv4
    port map (
            O => \N__34369\,
            I => n14278
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__34366\,
            I => \n14280_cascade_\
        );

    \I__6096\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34360\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__34360\,
            I => n14286
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__34357\,
            I => \N__34354\
        );

    \I__6093\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34350\
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__34353\,
            I => \N__34347\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__34350\,
            I => \N__34343\
        );

    \I__6090\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34340\
        );

    \I__6089\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34337\
        );

    \I__6088\ : Span4Mux_h
    port map (
            O => \N__34343\,
            I => \N__34334\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__34340\,
            I => \N__34331\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__34337\,
            I => \N__34328\
        );

    \I__6085\ : Odrv4
    port map (
            O => \N__34334\,
            I => n2522
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__34331\,
            I => n2522
        );

    \I__6083\ : Odrv4
    port map (
            O => \N__34328\,
            I => n2522
        );

    \I__6082\ : InMux
    port map (
            O => \N__34321\,
            I => \N__34318\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__34318\,
            I => \N__34315\
        );

    \I__6080\ : Span4Mux_h
    port map (
            O => \N__34315\,
            I => \N__34312\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__34312\,
            I => n2589
        );

    \I__6078\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34306\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__34306\,
            I => \N__34303\
        );

    \I__6076\ : Span4Mux_v
    port map (
            O => \N__34303\,
            I => \N__34300\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__34300\,
            I => n2597
        );

    \I__6074\ : CascadeMux
    port map (
            O => \N__34297\,
            I => \N__34293\
        );

    \I__6073\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34290\
        );

    \I__6072\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34287\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__34290\,
            I => \N__34284\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34281\
        );

    \I__6069\ : Span4Mux_h
    port map (
            O => \N__34284\,
            I => \N__34277\
        );

    \I__6068\ : Span4Mux_v
    port map (
            O => \N__34281\,
            I => \N__34274\
        );

    \I__6067\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34271\
        );

    \I__6066\ : Odrv4
    port map (
            O => \N__34277\,
            I => n2530
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__34274\,
            I => n2530
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__34271\,
            I => n2530
        );

    \I__6063\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34261\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__34261\,
            I => \N__34258\
        );

    \I__6061\ : Odrv4
    port map (
            O => \N__34258\,
            I => n898
        );

    \I__6060\ : CascadeMux
    port map (
            O => \N__34255\,
            I => \N__34252\
        );

    \I__6059\ : InMux
    port map (
            O => \N__34252\,
            I => \N__34247\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__34251\,
            I => \N__34244\
        );

    \I__6057\ : CascadeMux
    port map (
            O => \N__34250\,
            I => \N__34241\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__34247\,
            I => \N__34238\
        );

    \I__6055\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34235\
        );

    \I__6054\ : InMux
    port map (
            O => \N__34241\,
            I => \N__34232\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__34238\,
            I => n831
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__34235\,
            I => n831
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__34232\,
            I => n831
        );

    \I__6050\ : CascadeMux
    port map (
            O => \N__34225\,
            I => \N__34220\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__34224\,
            I => \N__34216\
        );

    \I__6048\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34211\
        );

    \I__6047\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34206\
        );

    \I__6046\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34206\
        );

    \I__6045\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34199\
        );

    \I__6044\ : InMux
    port map (
            O => \N__34215\,
            I => \N__34199\
        );

    \I__6043\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34199\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__34211\,
            I => n861
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__34206\,
            I => n861
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__34199\,
            I => n861
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__34192\,
            I => \N__34188\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__34191\,
            I => \N__34185\
        );

    \I__6037\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34182\
        );

    \I__6036\ : InMux
    port map (
            O => \N__34185\,
            I => \N__34179\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__34182\,
            I => n930
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__34179\,
            I => n930
        );

    \I__6033\ : CascadeMux
    port map (
            O => \N__34174\,
            I => \n930_cascade_\
        );

    \I__6032\ : InMux
    port map (
            O => \N__34171\,
            I => \N__34167\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__34170\,
            I => \N__34164\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34160\
        );

    \I__6029\ : InMux
    port map (
            O => \N__34164\,
            I => \N__34157\
        );

    \I__6028\ : InMux
    port map (
            O => \N__34163\,
            I => \N__34154\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__34160\,
            I => n929
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__34157\,
            I => n929
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__34154\,
            I => n929
        );

    \I__6024\ : CascadeMux
    port map (
            O => \N__34147\,
            I => \N__34143\
        );

    \I__6023\ : InMux
    port map (
            O => \N__34146\,
            I => \N__34140\
        );

    \I__6022\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34137\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__34140\,
            I => \N__34134\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__34137\,
            I => n927
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__34134\,
            I => n927
        );

    \I__6018\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34125\
        );

    \I__6017\ : CascadeMux
    port map (
            O => \N__34128\,
            I => \N__34122\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__34125\,
            I => \N__34118\
        );

    \I__6015\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34115\
        );

    \I__6014\ : InMux
    port map (
            O => \N__34121\,
            I => \N__34112\
        );

    \I__6013\ : Odrv4
    port map (
            O => \N__34118\,
            I => n928
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__34115\,
            I => n928
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__34112\,
            I => n928
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__34105\,
            I => \n13726_cascade_\
        );

    \I__6009\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34099\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__34099\,
            I => n11710
        );

    \I__6007\ : InMux
    port map (
            O => \N__34096\,
            I => \N__34093\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__34093\,
            I => n1000
        );

    \I__6005\ : CascadeMux
    port map (
            O => \N__34090\,
            I => \n960_cascade_\
        );

    \I__6004\ : CascadeMux
    port map (
            O => \N__34087\,
            I => \N__34083\
        );

    \I__6003\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34079\
        );

    \I__6002\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34076\
        );

    \I__6001\ : InMux
    port map (
            O => \N__34082\,
            I => \N__34073\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__34079\,
            I => n933
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__34076\,
            I => n933
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__34073\,
            I => n933
        );

    \I__5997\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34061\
        );

    \I__5996\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34058\
        );

    \I__5995\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34055\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__34061\,
            I => n295
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__34058\,
            I => n295
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__34055\,
            I => n295
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__34048\,
            I => \N__34045\
        );

    \I__5990\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34042\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__34042\,
            I => n1001
        );

    \I__5988\ : CascadeMux
    port map (
            O => \N__34039\,
            I => \N__34035\
        );

    \I__5987\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34031\
        );

    \I__5986\ : InMux
    port map (
            O => \N__34035\,
            I => \N__34028\
        );

    \I__5985\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34025\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__34031\,
            I => n931
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__34028\,
            I => n931
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__34025\,
            I => n931
        );

    \I__5981\ : InMux
    port map (
            O => \N__34018\,
            I => \N__34011\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__34017\,
            I => \N__34008\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__34016\,
            I => \N__34005\
        );

    \I__5978\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34000\
        );

    \I__5977\ : InMux
    port map (
            O => \N__34014\,
            I => \N__33997\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__34011\,
            I => \N__33994\
        );

    \I__5975\ : InMux
    port map (
            O => \N__34008\,
            I => \N__33985\
        );

    \I__5974\ : InMux
    port map (
            O => \N__34005\,
            I => \N__33985\
        );

    \I__5973\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33985\
        );

    \I__5972\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33985\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__34000\,
            I => n960
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__33997\,
            I => n960
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__33994\,
            I => n960
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__33985\,
            I => n960
        );

    \I__5967\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__33973\,
            I => n998
        );

    \I__5965\ : CascadeMux
    port map (
            O => \N__33970\,
            I => \N__33966\
        );

    \I__5964\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33962\
        );

    \I__5963\ : InMux
    port map (
            O => \N__33966\,
            I => \N__33959\
        );

    \I__5962\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33956\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__33962\,
            I => n1032
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__33959\,
            I => n1032
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__33956\,
            I => n1032
        );

    \I__5958\ : CascadeMux
    port map (
            O => \N__33949\,
            I => \N__33944\
        );

    \I__5957\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33941\
        );

    \I__5956\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33938\
        );

    \I__5955\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33935\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__33941\,
            I => n296
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__33938\,
            I => n296
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__33935\,
            I => n296
        );

    \I__5951\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33924\
        );

    \I__5950\ : CascadeMux
    port map (
            O => \N__33927\,
            I => \N__33921\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__33924\,
            I => \N__33917\
        );

    \I__5948\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33914\
        );

    \I__5947\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33911\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__33917\,
            I => n1033
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__33914\,
            I => n1033
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__33911\,
            I => n1033
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__33904\,
            I => \N__33901\
        );

    \I__5942\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33898\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33894\
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__33897\,
            I => \N__33891\
        );

    \I__5939\ : Span4Mux_s1_v
    port map (
            O => \N__33894\,
            I => \N__33887\
        );

    \I__5938\ : InMux
    port map (
            O => \N__33891\,
            I => \N__33884\
        );

    \I__5937\ : InMux
    port map (
            O => \N__33890\,
            I => \N__33881\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__33887\,
            I => n1031
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__33884\,
            I => n1031
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__33881\,
            I => n1031
        );

    \I__5933\ : CascadeMux
    port map (
            O => \N__33874\,
            I => \N__33870\
        );

    \I__5932\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33866\
        );

    \I__5931\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33863\
        );

    \I__5930\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33860\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__33866\,
            I => n1029
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__33863\,
            I => n1029
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__33860\,
            I => n1029
        );

    \I__5926\ : CascadeMux
    port map (
            O => \N__33853\,
            I => \n11646_cascade_\
        );

    \I__5925\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33846\
        );

    \I__5924\ : CascadeMux
    port map (
            O => \N__33849\,
            I => \N__33843\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__33846\,
            I => \N__33839\
        );

    \I__5922\ : InMux
    port map (
            O => \N__33843\,
            I => \N__33836\
        );

    \I__5921\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33833\
        );

    \I__5920\ : Odrv12
    port map (
            O => \N__33839\,
            I => n1030
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__33836\,
            I => n1030
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__33833\,
            I => n1030
        );

    \I__5917\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33823\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__33823\,
            I => n13323
        );

    \I__5915\ : InMux
    port map (
            O => \N__33820\,
            I => n12107
        );

    \I__5914\ : InMux
    port map (
            O => \N__33817\,
            I => n12108
        );

    \I__5913\ : InMux
    port map (
            O => \N__33814\,
            I => n12109
        );

    \I__5912\ : InMux
    port map (
            O => \N__33811\,
            I => n12110
        );

    \I__5911\ : CascadeMux
    port map (
            O => \N__33808\,
            I => \N__33805\
        );

    \I__5910\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33802\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__33802\,
            I => \N__33799\
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__33799\,
            I => n996
        );

    \I__5907\ : InMux
    port map (
            O => \N__33796\,
            I => n12111
        );

    \I__5906\ : CascadeMux
    port map (
            O => \N__33793\,
            I => \N__33790\
        );

    \I__5905\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33787\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__33787\,
            I => n995
        );

    \I__5903\ : InMux
    port map (
            O => \N__33784\,
            I => n12112
        );

    \I__5902\ : InMux
    port map (
            O => \N__33781\,
            I => n12113
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__33778\,
            I => \N__33775\
        );

    \I__5900\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33772\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__33772\,
            I => \N__33767\
        );

    \I__5898\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33762\
        );

    \I__5897\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33762\
        );

    \I__5896\ : Span4Mux_s2_v
    port map (
            O => \N__33767\,
            I => \N__33759\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33756\
        );

    \I__5894\ : Odrv4
    port map (
            O => \N__33759\,
            I => n1026
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__33756\,
            I => n1026
        );

    \I__5892\ : InMux
    port map (
            O => \N__33751\,
            I => \N__33748\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__33748\,
            I => n997
        );

    \I__5890\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33742\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__33742\,
            I => n999
        );

    \I__5888\ : InMux
    port map (
            O => \N__33739\,
            I => \N__33734\
        );

    \I__5887\ : CascadeMux
    port map (
            O => \N__33738\,
            I => \N__33731\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__33737\,
            I => \N__33728\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__33734\,
            I => \N__33725\
        );

    \I__5884\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33722\
        );

    \I__5883\ : InMux
    port map (
            O => \N__33728\,
            I => \N__33719\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__33725\,
            I => n932
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__33722\,
            I => n932
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__33719\,
            I => n932
        );

    \I__5879\ : InMux
    port map (
            O => \N__33712\,
            I => n12101
        );

    \I__5878\ : CascadeMux
    port map (
            O => \N__33709\,
            I => \N__33704\
        );

    \I__5877\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33699\
        );

    \I__5876\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33699\
        );

    \I__5875\ : InMux
    port map (
            O => \N__33704\,
            I => \N__33696\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__33699\,
            I => \N__33693\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__33696\,
            I => \N__33690\
        );

    \I__5872\ : Span4Mux_s3_v
    port map (
            O => \N__33693\,
            I => \N__33687\
        );

    \I__5871\ : Span4Mux_h
    port map (
            O => \N__33690\,
            I => \N__33684\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__33687\,
            I => n832
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__33684\,
            I => n832
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__33679\,
            I => \N__33676\
        );

    \I__5867\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33673\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__33673\,
            I => n899
        );

    \I__5865\ : InMux
    port map (
            O => \N__33670\,
            I => n12102
        );

    \I__5864\ : InMux
    port map (
            O => \N__33667\,
            I => n12103
        );

    \I__5863\ : CascadeMux
    port map (
            O => \N__33664\,
            I => \N__33661\
        );

    \I__5862\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33658\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__33658\,
            I => \N__33653\
        );

    \I__5860\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33648\
        );

    \I__5859\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33648\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__33653\,
            I => \N__33645\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__33648\,
            I => \N__33642\
        );

    \I__5856\ : Odrv4
    port map (
            O => \N__33645\,
            I => n830
        );

    \I__5855\ : Odrv4
    port map (
            O => \N__33642\,
            I => n830
        );

    \I__5854\ : CascadeMux
    port map (
            O => \N__33637\,
            I => \N__33634\
        );

    \I__5853\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33631\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__33631\,
            I => n897
        );

    \I__5851\ : InMux
    port map (
            O => \N__33628\,
            I => n12104
        );

    \I__5850\ : CascadeMux
    port map (
            O => \N__33625\,
            I => \N__33622\
        );

    \I__5849\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33617\
        );

    \I__5848\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33612\
        );

    \I__5847\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33612\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__33617\,
            I => n829
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__33612\,
            I => n829
        );

    \I__5844\ : InMux
    port map (
            O => \N__33607\,
            I => \N__33604\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__33604\,
            I => n896
        );

    \I__5842\ : InMux
    port map (
            O => \N__33601\,
            I => n12105
        );

    \I__5841\ : InMux
    port map (
            O => \N__33598\,
            I => \N__33594\
        );

    \I__5840\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33591\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__33594\,
            I => \N__33588\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__33591\,
            I => n828
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__33588\,
            I => n828
        );

    \I__5836\ : InMux
    port map (
            O => \N__33583\,
            I => n12106
        );

    \I__5835\ : InMux
    port map (
            O => \N__33580\,
            I => \N__33577\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__33577\,
            I => n900
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__33574\,
            I => \N__33569\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__33573\,
            I => \N__33566\
        );

    \I__5831\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33563\
        );

    \I__5830\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33558\
        );

    \I__5829\ : InMux
    port map (
            O => \N__33566\,
            I => \N__33558\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__33563\,
            I => n833
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__33558\,
            I => n833
        );

    \I__5826\ : InMux
    port map (
            O => \N__33553\,
            I => \bfn_7_30_0_\
        );

    \I__5825\ : CascadeMux
    port map (
            O => \N__33550\,
            I => \N__33547\
        );

    \I__5824\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33544\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33541\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__33541\,
            I => \N__33538\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__33538\,
            I => n8_adj_632
        );

    \I__5820\ : InMux
    port map (
            O => \N__33535\,
            I => n12599
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__33532\,
            I => \N__33529\
        );

    \I__5818\ : InMux
    port map (
            O => \N__33529\,
            I => \N__33526\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__33526\,
            I => n7_adj_631
        );

    \I__5816\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33517\
        );

    \I__5815\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33517\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__33517\,
            I => n7
        );

    \I__5813\ : InMux
    port map (
            O => \N__33514\,
            I => n12600
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__33511\,
            I => \N__33508\
        );

    \I__5811\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33505\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__33505\,
            I => \N__33502\
        );

    \I__5809\ : Span4Mux_h
    port map (
            O => \N__33502\,
            I => \N__33499\
        );

    \I__5808\ : Odrv4
    port map (
            O => \N__33499\,
            I => n6_adj_630
        );

    \I__5807\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__33493\,
            I => \N__33488\
        );

    \I__5805\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33485\
        );

    \I__5804\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33482\
        );

    \I__5803\ : Odrv4
    port map (
            O => \N__33488\,
            I => n6
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__33485\,
            I => n6
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__33482\,
            I => n6
        );

    \I__5800\ : InMux
    port map (
            O => \N__33475\,
            I => n12601
        );

    \I__5799\ : CascadeMux
    port map (
            O => \N__33472\,
            I => \N__33469\
        );

    \I__5798\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33466\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33463\
        );

    \I__5796\ : Span4Mux_v
    port map (
            O => \N__33463\,
            I => \N__33458\
        );

    \I__5795\ : InMux
    port map (
            O => \N__33462\,
            I => \N__33455\
        );

    \I__5794\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33452\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__33458\,
            I => n5
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__33455\,
            I => n5
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__33452\,
            I => n5
        );

    \I__5790\ : InMux
    port map (
            O => \N__33445\,
            I => n12602
        );

    \I__5789\ : CascadeMux
    port map (
            O => \N__33442\,
            I => \N__33439\
        );

    \I__5788\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33436\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33433\
        );

    \I__5786\ : Span4Mux_h
    port map (
            O => \N__33433\,
            I => \N__33430\
        );

    \I__5785\ : Odrv4
    port map (
            O => \N__33430\,
            I => n4_adj_628
        );

    \I__5784\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33424\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__33424\,
            I => \N__33421\
        );

    \I__5782\ : Span4Mux_h
    port map (
            O => \N__33421\,
            I => \N__33416\
        );

    \I__5781\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33411\
        );

    \I__5780\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33411\
        );

    \I__5779\ : Odrv4
    port map (
            O => \N__33416\,
            I => n4
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__33411\,
            I => n4
        );

    \I__5777\ : InMux
    port map (
            O => \N__33406\,
            I => n12603
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__33403\,
            I => \N__33400\
        );

    \I__5775\ : InMux
    port map (
            O => \N__33400\,
            I => \N__33397\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__33397\,
            I => n3_adj_627
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__33394\,
            I => \N__33389\
        );

    \I__5772\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33383\
        );

    \I__5771\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33383\
        );

    \I__5770\ : InMux
    port map (
            O => \N__33389\,
            I => \N__33378\
        );

    \I__5769\ : InMux
    port map (
            O => \N__33388\,
            I => \N__33378\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__33383\,
            I => n3_adj_567
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__33378\,
            I => n3_adj_567
        );

    \I__5766\ : InMux
    port map (
            O => \N__33373\,
            I => n12604
        );

    \I__5765\ : InMux
    port map (
            O => \N__33370\,
            I => n12605
        );

    \I__5764\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33364\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__33364\,
            I => \N__33359\
        );

    \I__5762\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33354\
        );

    \I__5761\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33354\
        );

    \I__5760\ : Span4Mux_h
    port map (
            O => \N__33359\,
            I => \N__33351\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__33354\,
            I => n2_adj_568
        );

    \I__5758\ : Odrv4
    port map (
            O => \N__33351\,
            I => n2_adj_568
        );

    \I__5757\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33343\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__33343\,
            I => n901
        );

    \I__5755\ : InMux
    port map (
            O => \N__33340\,
            I => \bfn_7_29_0_\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__33337\,
            I => \N__33334\
        );

    \I__5753\ : InMux
    port map (
            O => \N__33334\,
            I => \N__33331\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__33331\,
            I => \N__33328\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__33328\,
            I => n16_adj_640
        );

    \I__5750\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33322\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33319\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__33319\,
            I => n16
        );

    \I__5747\ : InMux
    port map (
            O => \N__33316\,
            I => n12591
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__33313\,
            I => \N__33310\
        );

    \I__5745\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33307\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__33307\,
            I => \N__33304\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__33304\,
            I => n15_adj_639
        );

    \I__5742\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33298\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__33298\,
            I => \N__33295\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__33295\,
            I => \N__33292\
        );

    \I__5739\ : Span4Mux_h
    port map (
            O => \N__33292\,
            I => \N__33289\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__33289\,
            I => n15
        );

    \I__5737\ : InMux
    port map (
            O => \N__33286\,
            I => n12592
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__33283\,
            I => \N__33280\
        );

    \I__5735\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33277\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__33277\,
            I => \N__33274\
        );

    \I__5733\ : Odrv12
    port map (
            O => \N__33274\,
            I => n14_adj_638
        );

    \I__5732\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33268\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__33268\,
            I => \N__33265\
        );

    \I__5730\ : Odrv12
    port map (
            O => \N__33265\,
            I => n14
        );

    \I__5729\ : InMux
    port map (
            O => \N__33262\,
            I => n12593
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__33259\,
            I => \N__33256\
        );

    \I__5727\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33253\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__33253\,
            I => \N__33250\
        );

    \I__5725\ : Span4Mux_h
    port map (
            O => \N__33250\,
            I => \N__33247\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__33247\,
            I => n13_adj_637
        );

    \I__5723\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33241\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33238\
        );

    \I__5721\ : Span4Mux_h
    port map (
            O => \N__33238\,
            I => \N__33235\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__33235\,
            I => n13
        );

    \I__5719\ : InMux
    port map (
            O => \N__33232\,
            I => n12594
        );

    \I__5718\ : CascadeMux
    port map (
            O => \N__33229\,
            I => \N__33226\
        );

    \I__5717\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33223\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__33223\,
            I => \N__33220\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__33220\,
            I => \N__33217\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__33217\,
            I => n12_adj_636
        );

    \I__5713\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33211\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__33211\,
            I => \N__33208\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__33208\,
            I => \N__33205\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__33205\,
            I => n12
        );

    \I__5709\ : InMux
    port map (
            O => \N__33202\,
            I => n12595
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__33199\,
            I => \N__33196\
        );

    \I__5707\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33193\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__33193\,
            I => \N__33190\
        );

    \I__5705\ : Span4Mux_h
    port map (
            O => \N__33190\,
            I => \N__33187\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__33187\,
            I => n11_adj_635
        );

    \I__5703\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33181\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__33181\,
            I => \N__33178\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__33178\,
            I => \N__33175\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__33175\,
            I => n11
        );

    \I__5699\ : InMux
    port map (
            O => \N__33172\,
            I => n12596
        );

    \I__5698\ : CascadeMux
    port map (
            O => \N__33169\,
            I => \N__33166\
        );

    \I__5697\ : InMux
    port map (
            O => \N__33166\,
            I => \N__33163\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__33163\,
            I => \N__33160\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__33160\,
            I => \N__33157\
        );

    \I__5694\ : Span4Mux_v
    port map (
            O => \N__33157\,
            I => \N__33154\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__33154\,
            I => n10_adj_634
        );

    \I__5692\ : CascadeMux
    port map (
            O => \N__33151\,
            I => \N__33148\
        );

    \I__5691\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33145\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__5689\ : Span4Mux_s2_v
    port map (
            O => \N__33142\,
            I => \N__33139\
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__33139\,
            I => n10
        );

    \I__5687\ : InMux
    port map (
            O => \N__33136\,
            I => n12597
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__33133\,
            I => \N__33130\
        );

    \I__5685\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33127\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__33127\,
            I => \N__33124\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__33124\,
            I => \N__33121\
        );

    \I__5682\ : Odrv4
    port map (
            O => \N__33121\,
            I => n9_adj_633
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__33118\,
            I => \N__33115\
        );

    \I__5680\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33112\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__33109\
        );

    \I__5678\ : Odrv4
    port map (
            O => \N__33109\,
            I => n9
        );

    \I__5677\ : InMux
    port map (
            O => \N__33106\,
            I => \bfn_7_28_0_\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__33103\,
            I => \N__33100\
        );

    \I__5675\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__33097\,
            I => n24_adj_648
        );

    \I__5673\ : InMux
    port map (
            O => \N__33094\,
            I => n12583
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__33091\,
            I => \N__33088\
        );

    \I__5671\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33085\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__33085\,
            I => \N__33082\
        );

    \I__5669\ : Span12Mux_v
    port map (
            O => \N__33082\,
            I => \N__33079\
        );

    \I__5668\ : Odrv12
    port map (
            O => \N__33079\,
            I => n23_adj_647
        );

    \I__5667\ : InMux
    port map (
            O => \N__33076\,
            I => n12584
        );

    \I__5666\ : CascadeMux
    port map (
            O => \N__33073\,
            I => \N__33070\
        );

    \I__5665\ : InMux
    port map (
            O => \N__33070\,
            I => \N__33067\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__33067\,
            I => \N__33064\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__33064\,
            I => n22_adj_646
        );

    \I__5662\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33058\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__33058\,
            I => \N__33055\
        );

    \I__5660\ : Odrv4
    port map (
            O => \N__33055\,
            I => n22
        );

    \I__5659\ : InMux
    port map (
            O => \N__33052\,
            I => n12585
        );

    \I__5658\ : CascadeMux
    port map (
            O => \N__33049\,
            I => \N__33046\
        );

    \I__5657\ : InMux
    port map (
            O => \N__33046\,
            I => \N__33043\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__33043\,
            I => \N__33040\
        );

    \I__5655\ : Span4Mux_h
    port map (
            O => \N__33040\,
            I => \N__33037\
        );

    \I__5654\ : Odrv4
    port map (
            O => \N__33037\,
            I => n21_adj_645
        );

    \I__5653\ : InMux
    port map (
            O => \N__33034\,
            I => \N__33031\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__33031\,
            I => \N__33028\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__33028\,
            I => n21
        );

    \I__5650\ : InMux
    port map (
            O => \N__33025\,
            I => n12586
        );

    \I__5649\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33019\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__33019\,
            I => \N__33016\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__33016\,
            I => n20
        );

    \I__5646\ : InMux
    port map (
            O => \N__33013\,
            I => n12587
        );

    \I__5645\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33007\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__33007\,
            I => n19_adj_643
        );

    \I__5643\ : InMux
    port map (
            O => \N__33004\,
            I => n12588
        );

    \I__5642\ : CascadeMux
    port map (
            O => \N__33001\,
            I => \N__32998\
        );

    \I__5641\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32995\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__32995\,
            I => n18_adj_642
        );

    \I__5639\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32989\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__32989\,
            I => \N__32986\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__32986\,
            I => n18
        );

    \I__5636\ : InMux
    port map (
            O => \N__32983\,
            I => n12589
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__32980\,
            I => \N__32977\
        );

    \I__5634\ : InMux
    port map (
            O => \N__32977\,
            I => \N__32974\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__32974\,
            I => n17_adj_641
        );

    \I__5632\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32968\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__32968\,
            I => \N__32965\
        );

    \I__5630\ : Span4Mux_h
    port map (
            O => \N__32965\,
            I => \N__32962\
        );

    \I__5629\ : Odrv4
    port map (
            O => \N__32962\,
            I => n17
        );

    \I__5628\ : InMux
    port map (
            O => \N__32959\,
            I => \bfn_7_27_0_\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__32956\,
            I => \N__32953\
        );

    \I__5626\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32950\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__32950\,
            I => n32_adj_656
        );

    \I__5624\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__32944\,
            I => n32
        );

    \I__5622\ : InMux
    port map (
            O => \N__32941\,
            I => n12575
        );

    \I__5621\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32935\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__32935\,
            I => \N__32932\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__32932\,
            I => n31_adj_655
        );

    \I__5618\ : InMux
    port map (
            O => \N__32929\,
            I => \N__32926\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__32926\,
            I => \N__32923\
        );

    \I__5616\ : Span4Mux_v
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__5615\ : Span4Mux_h
    port map (
            O => \N__32920\,
            I => \N__32917\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__32917\,
            I => n31
        );

    \I__5613\ : InMux
    port map (
            O => \N__32914\,
            I => n12576
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__32911\,
            I => \N__32908\
        );

    \I__5611\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32905\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32902\
        );

    \I__5609\ : Span4Mux_h
    port map (
            O => \N__32902\,
            I => \N__32899\
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__32899\,
            I => n30_adj_654
        );

    \I__5607\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32893\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__32893\,
            I => \N__32890\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__32890\,
            I => n30
        );

    \I__5604\ : InMux
    port map (
            O => \N__32887\,
            I => n12577
        );

    \I__5603\ : CascadeMux
    port map (
            O => \N__32884\,
            I => \N__32881\
        );

    \I__5602\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32878\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__32878\,
            I => \N__32875\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__32875\,
            I => n29_adj_653
        );

    \I__5599\ : InMux
    port map (
            O => \N__32872\,
            I => n12578
        );

    \I__5598\ : CascadeMux
    port map (
            O => \N__32869\,
            I => \N__32866\
        );

    \I__5597\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32863\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__32863\,
            I => n28_adj_652
        );

    \I__5595\ : InMux
    port map (
            O => \N__32860\,
            I => \N__32857\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__32857\,
            I => \N__32854\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__32854\,
            I => \N__32851\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__32851\,
            I => n28
        );

    \I__5591\ : InMux
    port map (
            O => \N__32848\,
            I => n12579
        );

    \I__5590\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32842\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__32842\,
            I => \N__32839\
        );

    \I__5588\ : Odrv12
    port map (
            O => \N__32839\,
            I => n27
        );

    \I__5587\ : InMux
    port map (
            O => \N__32836\,
            I => n12580
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__32833\,
            I => \N__32830\
        );

    \I__5585\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32827\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__32827\,
            I => n26_adj_650
        );

    \I__5583\ : InMux
    port map (
            O => \N__32824\,
            I => n12581
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__32821\,
            I => \N__32818\
        );

    \I__5581\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32815\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__32815\,
            I => n25_adj_649
        );

    \I__5579\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32809\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__32809\,
            I => \N__32806\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__32806\,
            I => n25
        );

    \I__5576\ : InMux
    port map (
            O => \N__32803\,
            I => \bfn_7_26_0_\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__32800\,
            I => \N__32796\
        );

    \I__5574\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32792\
        );

    \I__5573\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32789\
        );

    \I__5572\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32786\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__32792\,
            I => \N__32783\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__32789\,
            I => encoder0_position_8
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__32786\,
            I => encoder0_position_8
        );

    \I__5568\ : Odrv12
    port map (
            O => \N__32783\,
            I => encoder0_position_8
        );

    \I__5567\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32772\
        );

    \I__5566\ : InMux
    port map (
            O => \N__32775\,
            I => \N__32768\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32765\
        );

    \I__5564\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32762\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__32768\,
            I => \N__32759\
        );

    \I__5562\ : Sp12to4
    port map (
            O => \N__32765\,
            I => \N__32756\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__32762\,
            I => \N__32753\
        );

    \I__5560\ : Span4Mux_v
    port map (
            O => \N__32759\,
            I => \N__32750\
        );

    \I__5559\ : Span12Mux_v
    port map (
            O => \N__32756\,
            I => \N__32747\
        );

    \I__5558\ : Span4Mux_h
    port map (
            O => \N__32753\,
            I => \N__32744\
        );

    \I__5557\ : Odrv4
    port map (
            O => \N__32750\,
            I => n311
        );

    \I__5556\ : Odrv12
    port map (
            O => \N__32747\,
            I => n311
        );

    \I__5555\ : Odrv4
    port map (
            O => \N__32744\,
            I => n311
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__32737\,
            I => \N__32734\
        );

    \I__5553\ : InMux
    port map (
            O => \N__32734\,
            I => \N__32729\
        );

    \I__5552\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32726\
        );

    \I__5551\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32723\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__32729\,
            I => encoder0_position_5
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__32726\,
            I => encoder0_position_5
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__32723\,
            I => encoder0_position_5
        );

    \I__5547\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32711\
        );

    \I__5546\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32708\
        );

    \I__5545\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32705\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__32711\,
            I => \N__32702\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__32708\,
            I => encoder0_position_15
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__32705\,
            I => encoder0_position_15
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__32702\,
            I => encoder0_position_15
        );

    \I__5540\ : InMux
    port map (
            O => \N__32695\,
            I => \N__32691\
        );

    \I__5539\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32687\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__32691\,
            I => \N__32684\
        );

    \I__5537\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32681\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__32687\,
            I => \N__32678\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__32684\,
            I => \N__32675\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32672\
        );

    \I__5533\ : Span12Mux_s6_h
    port map (
            O => \N__32678\,
            I => \N__32669\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__32675\,
            I => n304
        );

    \I__5531\ : Odrv12
    port map (
            O => \N__32672\,
            I => n304
        );

    \I__5530\ : Odrv12
    port map (
            O => \N__32669\,
            I => n304
        );

    \I__5529\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32659\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__32659\,
            I => \N__32656\
        );

    \I__5527\ : Span4Mux_v
    port map (
            O => \N__32656\,
            I => \N__32652\
        );

    \I__5526\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32649\
        );

    \I__5525\ : Span4Mux_h
    port map (
            O => \N__32652\,
            I => \N__32646\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__32649\,
            I => n2320
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__32646\,
            I => n2320
        );

    \I__5522\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32637\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__32640\,
            I => \N__32634\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__32637\,
            I => \N__32631\
        );

    \I__5519\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32628\
        );

    \I__5518\ : Span12Mux_v
    port map (
            O => \N__32631\,
            I => \N__32625\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__32628\,
            I => n2319
        );

    \I__5516\ : Odrv12
    port map (
            O => \N__32625\,
            I => n2319
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__32620\,
            I => \N__32617\
        );

    \I__5514\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32614\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__32614\,
            I => n14008
        );

    \I__5512\ : InMux
    port map (
            O => \N__32611\,
            I => \N__32608\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__32608\,
            I => n14006
        );

    \I__5510\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32602\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__32602\,
            I => \N__32599\
        );

    \I__5508\ : Span4Mux_h
    port map (
            O => \N__32599\,
            I => \N__32596\
        );

    \I__5507\ : Span4Mux_v
    port map (
            O => \N__32596\,
            I => \N__32593\
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__32593\,
            I => n14014
        );

    \I__5505\ : CascadeMux
    port map (
            O => \N__32590\,
            I => \N__32587\
        );

    \I__5504\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32582\
        );

    \I__5503\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32577\
        );

    \I__5502\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32577\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__32582\,
            I => encoder0_position_1
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__32577\,
            I => encoder0_position_1
        );

    \I__5499\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32569\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__32569\,
            I => \N__32565\
        );

    \I__5497\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32561\
        );

    \I__5496\ : Span4Mux_v
    port map (
            O => \N__32565\,
            I => \N__32558\
        );

    \I__5495\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32555\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__32561\,
            I => encoder0_position_0
        );

    \I__5493\ : Odrv4
    port map (
            O => \N__32558\,
            I => encoder0_position_0
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__32555\,
            I => encoder0_position_0
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__32548\,
            I => \N__32545\
        );

    \I__5490\ : InMux
    port map (
            O => \N__32545\,
            I => \N__32542\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__32542\,
            I => n33_adj_657
        );

    \I__5488\ : CascadeMux
    port map (
            O => \N__32539\,
            I => \N__32536\
        );

    \I__5487\ : InMux
    port map (
            O => \N__32536\,
            I => \N__32533\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__32533\,
            I => \N__32530\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__32530\,
            I => \N__32527\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__32527\,
            I => n33
        );

    \I__5483\ : InMux
    port map (
            O => \N__32524\,
            I => \bfn_7_25_0_\
        );

    \I__5482\ : InMux
    port map (
            O => \N__32521\,
            I => \N__32518\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32515\
        );

    \I__5480\ : Odrv4
    port map (
            O => \N__32515\,
            I => n2295
        );

    \I__5479\ : CascadeMux
    port map (
            O => \N__32512\,
            I => \N__32508\
        );

    \I__5478\ : CascadeMux
    port map (
            O => \N__32511\,
            I => \N__32505\
        );

    \I__5477\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32502\
        );

    \I__5476\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32499\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__32502\,
            I => \N__32495\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__32499\,
            I => \N__32492\
        );

    \I__5473\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32489\
        );

    \I__5472\ : Span4Mux_v
    port map (
            O => \N__32495\,
            I => \N__32482\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__32492\,
            I => \N__32482\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__32489\,
            I => \N__32482\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__32482\,
            I => n2228
        );

    \I__5468\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32476\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__32476\,
            I => \N__32472\
        );

    \I__5466\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32468\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__32472\,
            I => \N__32465\
        );

    \I__5464\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32462\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__32468\,
            I => encoder0_position_2
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__32465\,
            I => encoder0_position_2
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__32462\,
            I => encoder0_position_2
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__32455\,
            I => \N__32452\
        );

    \I__5459\ : InMux
    port map (
            O => \N__32452\,
            I => \N__32448\
        );

    \I__5458\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32444\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32441\
        );

    \I__5456\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32438\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__32444\,
            I => \N__32433\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__32441\,
            I => \N__32433\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__32438\,
            I => \N__32430\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__32433\,
            I => n2321
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__32430\,
            I => n2321
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__32425\,
            I => \N__32422\
        );

    \I__5449\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32418\
        );

    \I__5448\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32415\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32412\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__32415\,
            I => \N__32408\
        );

    \I__5445\ : Span4Mux_h
    port map (
            O => \N__32412\,
            I => \N__32405\
        );

    \I__5444\ : InMux
    port map (
            O => \N__32411\,
            I => \N__32402\
        );

    \I__5443\ : Odrv12
    port map (
            O => \N__32408\,
            I => n2324
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__32405\,
            I => n2324
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__32402\,
            I => n2324
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__32395\,
            I => \N__32391\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__32394\,
            I => \N__32388\
        );

    \I__5438\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32385\
        );

    \I__5437\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32381\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__32385\,
            I => \N__32378\
        );

    \I__5435\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32375\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32372\
        );

    \I__5433\ : Span4Mux_h
    port map (
            O => \N__32378\,
            I => \N__32369\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__32375\,
            I => n2328
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__32372\,
            I => n2328
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__32369\,
            I => n2328
        );

    \I__5429\ : CascadeMux
    port map (
            O => \N__32362\,
            I => \N__32359\
        );

    \I__5428\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32355\
        );

    \I__5427\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32352\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__32355\,
            I => \N__32349\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__32352\,
            I => \N__32343\
        );

    \I__5424\ : Span12Mux_s6_h
    port map (
            O => \N__32349\,
            I => \N__32343\
        );

    \I__5423\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32340\
        );

    \I__5422\ : Odrv12
    port map (
            O => \N__32343\,
            I => n2327
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__32340\,
            I => n2327
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__32335\,
            I => \N__32331\
        );

    \I__5419\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32328\
        );

    \I__5418\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32325\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__32328\,
            I => \N__32322\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__32325\,
            I => \N__32319\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__32322\,
            I => \N__32315\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__32319\,
            I => \N__32312\
        );

    \I__5413\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32309\
        );

    \I__5412\ : Odrv4
    port map (
            O => \N__32315\,
            I => n2322
        );

    \I__5411\ : Odrv4
    port map (
            O => \N__32312\,
            I => n2322
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__32309\,
            I => n2322
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__32302\,
            I => \N__32299\
        );

    \I__5408\ : InMux
    port map (
            O => \N__32299\,
            I => \N__32295\
        );

    \I__5407\ : InMux
    port map (
            O => \N__32298\,
            I => \N__32292\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__32295\,
            I => \N__32289\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__32292\,
            I => \N__32286\
        );

    \I__5404\ : Span4Mux_v
    port map (
            O => \N__32289\,
            I => \N__32281\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__32286\,
            I => \N__32281\
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__32281\,
            I => n2326
        );

    \I__5401\ : CascadeMux
    port map (
            O => \N__32278\,
            I => \N__32273\
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__32277\,
            I => \N__32270\
        );

    \I__5399\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32267\
        );

    \I__5398\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32264\
        );

    \I__5397\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32261\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__32267\,
            I => \N__32256\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__32264\,
            I => \N__32256\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__32261\,
            I => \N__32253\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__32256\,
            I => \N__32248\
        );

    \I__5392\ : Span4Mux_v
    port map (
            O => \N__32253\,
            I => \N__32248\
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__32248\,
            I => n2325
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__32245\,
            I => \N__32242\
        );

    \I__5389\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32238\
        );

    \I__5388\ : InMux
    port map (
            O => \N__32241\,
            I => \N__32235\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__32238\,
            I => \N__32232\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__32235\,
            I => \N__32229\
        );

    \I__5385\ : Span4Mux_s3_h
    port map (
            O => \N__32232\,
            I => \N__32226\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__32229\,
            I => \N__32222\
        );

    \I__5383\ : Span4Mux_v
    port map (
            O => \N__32226\,
            I => \N__32219\
        );

    \I__5382\ : InMux
    port map (
            O => \N__32225\,
            I => \N__32216\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__32222\,
            I => n2323
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__32219\,
            I => n2323
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__32216\,
            I => n2323
        );

    \I__5378\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32205\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__32208\,
            I => \N__32202\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32198\
        );

    \I__5375\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32195\
        );

    \I__5374\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32192\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__32198\,
            I => \N__32189\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__32195\,
            I => encoder0_position_3
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__32192\,
            I => encoder0_position_3
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__32189\,
            I => encoder0_position_3
        );

    \I__5369\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32177\
        );

    \I__5368\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32174\
        );

    \I__5367\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32171\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__32177\,
            I => \N__32168\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__32174\,
            I => encoder0_position_11
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__32171\,
            I => encoder0_position_11
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__32168\,
            I => encoder0_position_11
        );

    \I__5362\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32157\
        );

    \I__5361\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32154\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__32157\,
            I => \N__32149\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__32154\,
            I => \N__32149\
        );

    \I__5358\ : Span4Mux_h
    port map (
            O => \N__32149\,
            I => \N__32145\
        );

    \I__5357\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32142\
        );

    \I__5356\ : Span4Mux_s3_h
    port map (
            O => \N__32145\,
            I => \N__32137\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__32142\,
            I => \N__32137\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__32137\,
            I => \N__32134\
        );

    \I__5353\ : Odrv4
    port map (
            O => \N__32134\,
            I => n308
        );

    \I__5352\ : InMux
    port map (
            O => \N__32131\,
            I => n12289
        );

    \I__5351\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32125\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__32125\,
            I => \N__32122\
        );

    \I__5349\ : Span4Mux_v
    port map (
            O => \N__32122\,
            I => \N__32118\
        );

    \I__5348\ : InMux
    port map (
            O => \N__32121\,
            I => \N__32115\
        );

    \I__5347\ : Odrv4
    port map (
            O => \N__32118\,
            I => n2219
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__32115\,
            I => n2219
        );

    \I__5345\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32107\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__32107\,
            I => \N__32104\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__32104\,
            I => \N__32101\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__32101\,
            I => n2286_adj_600
        );

    \I__5341\ : InMux
    port map (
            O => \N__32098\,
            I => n12290
        );

    \I__5340\ : InMux
    port map (
            O => \N__32095\,
            I => \N__32092\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__32092\,
            I => \N__32089\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__32089\,
            I => \N__32084\
        );

    \I__5337\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32079\
        );

    \I__5336\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32079\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__32084\,
            I => n2218
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__32079\,
            I => n2218
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__32074\,
            I => \N__32071\
        );

    \I__5332\ : InMux
    port map (
            O => \N__32071\,
            I => \N__32068\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__32068\,
            I => \N__32065\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__32065\,
            I => \N__32062\
        );

    \I__5329\ : Span4Mux_h
    port map (
            O => \N__32062\,
            I => \N__32059\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__32059\,
            I => n2285_adj_599
        );

    \I__5327\ : InMux
    port map (
            O => \N__32056\,
            I => \bfn_7_22_0_\
        );

    \I__5326\ : InMux
    port map (
            O => \N__32053\,
            I => n12292
        );

    \I__5325\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32047\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32043\
        );

    \I__5323\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32040\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__32043\,
            I => \N__32036\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__32033\
        );

    \I__5320\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32030\
        );

    \I__5319\ : Span4Mux_h
    port map (
            O => \N__32036\,
            I => \N__32027\
        );

    \I__5318\ : Span4Mux_v
    port map (
            O => \N__32033\,
            I => \N__32022\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__32022\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__32027\,
            I => n2216
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__32022\,
            I => n2216
        );

    \I__5314\ : InMux
    port map (
            O => \N__32017\,
            I => \N__32014\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__32014\,
            I => n2283
        );

    \I__5312\ : InMux
    port map (
            O => \N__32011\,
            I => n12293
        );

    \I__5311\ : CascadeMux
    port map (
            O => \N__32008\,
            I => \N__32004\
        );

    \I__5310\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32001\
        );

    \I__5309\ : InMux
    port map (
            O => \N__32004\,
            I => \N__31998\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31995\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__31998\,
            I => \N__31992\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__31995\,
            I => \N__31988\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__31992\,
            I => \N__31985\
        );

    \I__5304\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31982\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__31988\,
            I => \N__31979\
        );

    \I__5302\ : Span4Mux_h
    port map (
            O => \N__31985\,
            I => \N__31974\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31974\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__31979\,
            I => n2215
        );

    \I__5299\ : Odrv4
    port map (
            O => \N__31974\,
            I => n2215
        );

    \I__5298\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31966\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__31966\,
            I => \N__31963\
        );

    \I__5296\ : Span4Mux_v
    port map (
            O => \N__31963\,
            I => \N__31960\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__31960\,
            I => n2282
        );

    \I__5294\ : InMux
    port map (
            O => \N__31957\,
            I => n12294
        );

    \I__5293\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31950\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__31953\,
            I => \N__31947\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31944\
        );

    \I__5290\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31941\
        );

    \I__5289\ : Span4Mux_h
    port map (
            O => \N__31944\,
            I => \N__31938\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__31941\,
            I => \N__31935\
        );

    \I__5287\ : Span4Mux_h
    port map (
            O => \N__31938\,
            I => \N__31932\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__31935\,
            I => \N__31929\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__31932\,
            I => n2214
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__31929\,
            I => n2214
        );

    \I__5283\ : InMux
    port map (
            O => \N__31924\,
            I => n12295
        );

    \I__5282\ : CascadeMux
    port map (
            O => \N__31921\,
            I => \N__31918\
        );

    \I__5281\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31914\
        );

    \I__5280\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31911\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__31914\,
            I => \N__31906\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__31911\,
            I => \N__31906\
        );

    \I__5277\ : Span4Mux_v
    port map (
            O => \N__31906\,
            I => \N__31903\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__31903\,
            I => n2313
        );

    \I__5275\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31896\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__31899\,
            I => \N__31893\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__31896\,
            I => \N__31889\
        );

    \I__5272\ : InMux
    port map (
            O => \N__31893\,
            I => \N__31886\
        );

    \I__5271\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31883\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__31889\,
            I => n2225
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__31886\,
            I => n2225
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__31883\,
            I => n2225
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__31876\,
            I => \N__31873\
        );

    \I__5266\ : InMux
    port map (
            O => \N__31873\,
            I => \N__31870\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__31870\,
            I => n2292
        );

    \I__5264\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31863\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__31866\,
            I => \N__31860\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31857\
        );

    \I__5261\ : InMux
    port map (
            O => \N__31860\,
            I => \N__31854\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__31857\,
            I => n2224
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__31854\,
            I => n2224
        );

    \I__5258\ : InMux
    port map (
            O => \N__31849\,
            I => \N__31846\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__31846\,
            I => n2291
        );

    \I__5256\ : InMux
    port map (
            O => \N__31843\,
            I => n12281
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__31840\,
            I => \N__31836\
        );

    \I__5254\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31832\
        );

    \I__5253\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31829\
        );

    \I__5252\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31826\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__31832\,
            I => \N__31819\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31819\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__31826\,
            I => \N__31819\
        );

    \I__5248\ : Odrv12
    port map (
            O => \N__31819\,
            I => n2227
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__31816\,
            I => \N__31813\
        );

    \I__5246\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31810\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__31810\,
            I => \N__31807\
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__31807\,
            I => n2294
        );

    \I__5243\ : InMux
    port map (
            O => \N__31804\,
            I => n12282
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__31801\,
            I => \N__31797\
        );

    \I__5241\ : CascadeMux
    port map (
            O => \N__31800\,
            I => \N__31794\
        );

    \I__5240\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31790\
        );

    \I__5239\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31787\
        );

    \I__5238\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31784\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__31790\,
            I => n2226
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__31787\,
            I => n2226
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__31784\,
            I => n2226
        );

    \I__5234\ : InMux
    port map (
            O => \N__31777\,
            I => \N__31774\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__31774\,
            I => n2293
        );

    \I__5232\ : InMux
    port map (
            O => \N__31771\,
            I => \bfn_7_21_0_\
        );

    \I__5231\ : InMux
    port map (
            O => \N__31768\,
            I => n12284
        );

    \I__5230\ : InMux
    port map (
            O => \N__31765\,
            I => n12285
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__31762\,
            I => \N__31758\
        );

    \I__5228\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31755\
        );

    \I__5227\ : InMux
    port map (
            O => \N__31758\,
            I => \N__31752\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__31755\,
            I => \N__31749\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__31752\,
            I => n2223
        );

    \I__5224\ : Odrv4
    port map (
            O => \N__31749\,
            I => n2223
        );

    \I__5223\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31741\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__31741\,
            I => n2290_adj_604
        );

    \I__5221\ : InMux
    port map (
            O => \N__31738\,
            I => n12286
        );

    \I__5220\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31731\
        );

    \I__5219\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31727\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31724\
        );

    \I__5217\ : InMux
    port map (
            O => \N__31730\,
            I => \N__31721\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__31727\,
            I => n2222
        );

    \I__5215\ : Odrv12
    port map (
            O => \N__31724\,
            I => n2222
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__31721\,
            I => n2222
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__31714\,
            I => \N__31711\
        );

    \I__5212\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31708\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__31708\,
            I => n2289_adj_603
        );

    \I__5210\ : InMux
    port map (
            O => \N__31705\,
            I => n12287
        );

    \I__5209\ : InMux
    port map (
            O => \N__31702\,
            I => \N__31698\
        );

    \I__5208\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31695\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__31698\,
            I => \N__31692\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__31695\,
            I => \N__31689\
        );

    \I__5205\ : Span4Mux_v
    port map (
            O => \N__31692\,
            I => \N__31686\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__31689\,
            I => \N__31683\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__31686\,
            I => n2221
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__31683\,
            I => n2221
        );

    \I__5201\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31675\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__31675\,
            I => \N__31672\
        );

    \I__5199\ : Span4Mux_h
    port map (
            O => \N__31672\,
            I => \N__31669\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__31669\,
            I => n2288_adj_602
        );

    \I__5197\ : InMux
    port map (
            O => \N__31666\,
            I => n12288
        );

    \I__5196\ : InMux
    port map (
            O => \N__31663\,
            I => \N__31660\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__31660\,
            I => \N__31656\
        );

    \I__5194\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31653\
        );

    \I__5193\ : Span4Mux_v
    port map (
            O => \N__31656\,
            I => \N__31648\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__31653\,
            I => \N__31648\
        );

    \I__5191\ : Span4Mux_h
    port map (
            O => \N__31648\,
            I => \N__31645\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__31645\,
            I => n2220
        );

    \I__5189\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31639\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__31639\,
            I => \N__31636\
        );

    \I__5187\ : Span4Mux_s2_h
    port map (
            O => \N__31636\,
            I => \N__31633\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__31633\,
            I => \N__31630\
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__31630\,
            I => n2287_adj_601
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__31627\,
            I => \N__31624\
        );

    \I__5183\ : InMux
    port map (
            O => \N__31624\,
            I => \N__31620\
        );

    \I__5182\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31616\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__31620\,
            I => \N__31613\
        );

    \I__5180\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31610\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__31616\,
            I => n2532
        );

    \I__5178\ : Odrv12
    port map (
            O => \N__31613\,
            I => n2532
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__31610\,
            I => n2532
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__5175\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31597\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__31597\,
            I => \N__31594\
        );

    \I__5173\ : Span4Mux_v
    port map (
            O => \N__31594\,
            I => \N__31591\
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__31591\,
            I => n2599
        );

    \I__5171\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31585\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__31585\,
            I => n2483
        );

    \I__5169\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31579\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__31579\,
            I => \N__31575\
        );

    \I__5167\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31572\
        );

    \I__5166\ : Span4Mux_h
    port map (
            O => \N__31575\,
            I => \N__31568\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__31572\,
            I => \N__31565\
        );

    \I__5164\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31562\
        );

    \I__5163\ : Odrv4
    port map (
            O => \N__31568\,
            I => n2416
        );

    \I__5162\ : Odrv4
    port map (
            O => \N__31565\,
            I => n2416
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__31562\,
            I => n2416
        );

    \I__5160\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31552\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__31552\,
            I => \N__31549\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__31549\,
            I => \N__31544\
        );

    \I__5157\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31539\
        );

    \I__5156\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31539\
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__31544\,
            I => n2515
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__31539\,
            I => n2515
        );

    \I__5153\ : InMux
    port map (
            O => \N__31534\,
            I => \N__31531\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__31531\,
            I => \N__31528\
        );

    \I__5151\ : Odrv12
    port map (
            O => \N__31528\,
            I => n2301
        );

    \I__5150\ : InMux
    port map (
            O => \N__31525\,
            I => \bfn_7_20_0_\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__31522\,
            I => \N__31518\
        );

    \I__5148\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31514\
        );

    \I__5147\ : InMux
    port map (
            O => \N__31518\,
            I => \N__31511\
        );

    \I__5146\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31508\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__31514\,
            I => \N__31503\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31503\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__31508\,
            I => n2233
        );

    \I__5142\ : Odrv12
    port map (
            O => \N__31503\,
            I => n2233
        );

    \I__5141\ : CascadeMux
    port map (
            O => \N__31498\,
            I => \N__31495\
        );

    \I__5140\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31492\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__31492\,
            I => \N__31489\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__31489\,
            I => \N__31486\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__31486\,
            I => n2300
        );

    \I__5136\ : InMux
    port map (
            O => \N__31483\,
            I => n12276
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__31480\,
            I => \N__31477\
        );

    \I__5134\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31473\
        );

    \I__5133\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31470\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__31473\,
            I => \N__31467\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__31470\,
            I => \N__31462\
        );

    \I__5130\ : Span4Mux_h
    port map (
            O => \N__31467\,
            I => \N__31462\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__31462\,
            I => \N__31459\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__31459\,
            I => n2232
        );

    \I__5127\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31453\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__31453\,
            I => \N__31450\
        );

    \I__5125\ : Span12Mux_s6_h
    port map (
            O => \N__31450\,
            I => \N__31447\
        );

    \I__5124\ : Odrv12
    port map (
            O => \N__31447\,
            I => n2299
        );

    \I__5123\ : InMux
    port map (
            O => \N__31444\,
            I => n12277
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__31441\,
            I => \N__31438\
        );

    \I__5121\ : InMux
    port map (
            O => \N__31438\,
            I => \N__31434\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__31437\,
            I => \N__31430\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__31434\,
            I => \N__31427\
        );

    \I__5118\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31422\
        );

    \I__5117\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31422\
        );

    \I__5116\ : Span4Mux_h
    port map (
            O => \N__31427\,
            I => \N__31419\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__31422\,
            I => n2231
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__31419\,
            I => n2231
        );

    \I__5113\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31411\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__31411\,
            I => \N__31408\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__31408\,
            I => n2298
        );

    \I__5110\ : InMux
    port map (
            O => \N__31405\,
            I => n12278
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__31402\,
            I => \N__31399\
        );

    \I__5108\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31396\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__31396\,
            I => \N__31392\
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__31395\,
            I => \N__31389\
        );

    \I__5105\ : Span4Mux_v
    port map (
            O => \N__31392\,
            I => \N__31386\
        );

    \I__5104\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31383\
        );

    \I__5103\ : Odrv4
    port map (
            O => \N__31386\,
            I => n2230
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__31383\,
            I => n2230
        );

    \I__5101\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31375\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__5099\ : Span4Mux_v
    port map (
            O => \N__31372\,
            I => \N__31369\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__31369\,
            I => n2297
        );

    \I__5097\ : InMux
    port map (
            O => \N__31366\,
            I => n12279
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__31363\,
            I => \N__31359\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__31362\,
            I => \N__31355\
        );

    \I__5094\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31352\
        );

    \I__5093\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31349\
        );

    \I__5092\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31346\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__31352\,
            I => \N__31343\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31340\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__31346\,
            I => n2229
        );

    \I__5088\ : Odrv12
    port map (
            O => \N__31343\,
            I => n2229
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__31340\,
            I => n2229
        );

    \I__5086\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31330\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__31330\,
            I => \N__31327\
        );

    \I__5084\ : Odrv12
    port map (
            O => \N__31327\,
            I => n2296
        );

    \I__5083\ : InMux
    port map (
            O => \N__31324\,
            I => n12280
        );

    \I__5082\ : InMux
    port map (
            O => \N__31321\,
            I => \N__31318\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__31318\,
            I => \N__31315\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__31315\,
            I => n2591
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__31312\,
            I => \n2524_cascade_\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__31309\,
            I => \N__31306\
        );

    \I__5077\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31303\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__31303\,
            I => \N__31300\
        );

    \I__5075\ : Odrv12
    port map (
            O => \N__31300\,
            I => n2391
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__31297\,
            I => \N__31293\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__31296\,
            I => \N__31289\
        );

    \I__5072\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31286\
        );

    \I__5071\ : InMux
    port map (
            O => \N__31292\,
            I => \N__31283\
        );

    \I__5070\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31280\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__31286\,
            I => \N__31275\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__31283\,
            I => \N__31275\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__31280\,
            I => n2423
        );

    \I__5066\ : Odrv4
    port map (
            O => \N__31275\,
            I => n2423
        );

    \I__5065\ : InMux
    port map (
            O => \N__31270\,
            I => \N__31267\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__31267\,
            I => \N__31264\
        );

    \I__5063\ : Span4Mux_v
    port map (
            O => \N__31264\,
            I => \N__31261\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__31261\,
            I => n2601
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__31258\,
            I => \N__31255\
        );

    \I__5060\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31252\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31249\
        );

    \I__5058\ : Span4Mux_h
    port map (
            O => \N__31249\,
            I => \N__31246\
        );

    \I__5057\ : Span4Mux_h
    port map (
            O => \N__31246\,
            I => \N__31243\
        );

    \I__5056\ : Odrv4
    port map (
            O => \N__31243\,
            I => n2394
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__31240\,
            I => \N__31236\
        );

    \I__5054\ : CascadeMux
    port map (
            O => \N__31239\,
            I => \N__31233\
        );

    \I__5053\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31229\
        );

    \I__5052\ : InMux
    port map (
            O => \N__31233\,
            I => \N__31226\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__31232\,
            I => \N__31223\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__31229\,
            I => \N__31218\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__31226\,
            I => \N__31218\
        );

    \I__5048\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31215\
        );

    \I__5047\ : Span4Mux_v
    port map (
            O => \N__31218\,
            I => \N__31212\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__31215\,
            I => n2426
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__31212\,
            I => n2426
        );

    \I__5044\ : InMux
    port map (
            O => \N__31207\,
            I => \N__31204\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__31204\,
            I => n2480
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__31201\,
            I => \N__31198\
        );

    \I__5041\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31195\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__31195\,
            I => \N__31190\
        );

    \I__5039\ : InMux
    port map (
            O => \N__31194\,
            I => \N__31187\
        );

    \I__5038\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31184\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__31190\,
            I => n2413
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__31187\,
            I => n2413
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__31184\,
            I => n2413
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__31177\,
            I => \N__31174\
        );

    \I__5033\ : InMux
    port map (
            O => \N__31174\,
            I => \N__31171\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__31171\,
            I => \N__31166\
        );

    \I__5031\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31161\
        );

    \I__5030\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31161\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__31166\,
            I => n2512
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__31161\,
            I => n2512
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__31156\,
            I => \N__31153\
        );

    \I__5026\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31150\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__31150\,
            I => \N__31147\
        );

    \I__5024\ : Span4Mux_v
    port map (
            O => \N__31147\,
            I => \N__31144\
        );

    \I__5023\ : Span4Mux_h
    port map (
            O => \N__31144\,
            I => \N__31141\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__31141\,
            I => n2388
        );

    \I__5021\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31134\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__31137\,
            I => \N__31131\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31128\
        );

    \I__5018\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31125\
        );

    \I__5017\ : Span4Mux_h
    port map (
            O => \N__31128\,
            I => \N__31122\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__31125\,
            I => n2420
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__31122\,
            I => n2420
        );

    \I__5014\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31114\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__31114\,
            I => n2487
        );

    \I__5012\ : CascadeMux
    port map (
            O => \N__31111\,
            I => \n2420_cascade_\
        );

    \I__5011\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31104\
        );

    \I__5010\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31101\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__31104\,
            I => \N__31098\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__31101\,
            I => \N__31095\
        );

    \I__5007\ : Span4Mux_h
    port map (
            O => \N__31098\,
            I => \N__31092\
        );

    \I__5006\ : Span4Mux_h
    port map (
            O => \N__31095\,
            I => \N__31089\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__31092\,
            I => n2519
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__31089\,
            I => n2519
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__31084\,
            I => \n2519_cascade_\
        );

    \I__5002\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31078\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__31078\,
            I => \N__31075\
        );

    \I__5000\ : Span4Mux_v
    port map (
            O => \N__31075\,
            I => \N__31072\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__31072\,
            I => n2586
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__31069\,
            I => \n2628_cascade_\
        );

    \I__4997\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31063\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__31063\,
            I => n2585
        );

    \I__4995\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31057\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__31057\,
            I => \N__31053\
        );

    \I__4993\ : InMux
    port map (
            O => \N__31056\,
            I => \N__31050\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__31053\,
            I => \N__31046\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__31050\,
            I => \N__31043\
        );

    \I__4990\ : InMux
    port map (
            O => \N__31049\,
            I => \N__31040\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__31046\,
            I => n2518
        );

    \I__4988\ : Odrv4
    port map (
            O => \N__31043\,
            I => n2518
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__31040\,
            I => n2518
        );

    \I__4986\ : InMux
    port map (
            O => \N__31033\,
            I => \N__31029\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31026\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__31029\,
            I => \N__31023\
        );

    \I__4983\ : InMux
    port map (
            O => \N__31026\,
            I => \N__31020\
        );

    \I__4982\ : Span4Mux_v
    port map (
            O => \N__31023\,
            I => \N__31014\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__31020\,
            I => \N__31014\
        );

    \I__4980\ : InMux
    port map (
            O => \N__31019\,
            I => \N__31011\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__31014\,
            I => n2417
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__31011\,
            I => n2417
        );

    \I__4977\ : InMux
    port map (
            O => \N__31006\,
            I => \N__31003\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__31003\,
            I => n2484
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__31000\,
            I => \N__30997\
        );

    \I__4974\ : InMux
    port map (
            O => \N__30997\,
            I => \N__30994\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__30994\,
            I => \N__30990\
        );

    \I__4972\ : InMux
    port map (
            O => \N__30993\,
            I => \N__30987\
        );

    \I__4971\ : Span4Mux_v
    port map (
            O => \N__30990\,
            I => \N__30984\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__30987\,
            I => \N__30981\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__30984\,
            I => \N__30976\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__30981\,
            I => \N__30976\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__30976\,
            I => n2516
        );

    \I__4966\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30968\
        );

    \I__4965\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30965\
        );

    \I__4964\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30962\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__30968\,
            I => \N__30959\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__30965\,
            I => \N__30954\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__30962\,
            I => \N__30954\
        );

    \I__4960\ : Span4Mux_v
    port map (
            O => \N__30959\,
            I => \N__30951\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__30954\,
            I => n2514
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__30951\,
            I => n2514
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__30946\,
            I => \n2516_cascade_\
        );

    \I__4956\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30940\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__30940\,
            I => \N__30937\
        );

    \I__4954\ : Odrv4
    port map (
            O => \N__30937\,
            I => n13810
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__30934\,
            I => \n13816_cascade_\
        );

    \I__4952\ : InMux
    port map (
            O => \N__30931\,
            I => \N__30928\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__30928\,
            I => \N__30924\
        );

    \I__4950\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30921\
        );

    \I__4949\ : Odrv12
    port map (
            O => \N__30924\,
            I => n2511
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__30921\,
            I => n2511
        );

    \I__4947\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30913\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30910\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__30910\,
            I => n2582
        );

    \I__4944\ : CascadeMux
    port map (
            O => \N__30907\,
            I => \n2544_cascade_\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__30904\,
            I => \N__30901\
        );

    \I__4942\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30898\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__30898\,
            I => \N__30895\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__30895\,
            I => n2579
        );

    \I__4939\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30888\
        );

    \I__4938\ : CascadeMux
    port map (
            O => \N__30891\,
            I => \N__30885\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__30888\,
            I => \N__30881\
        );

    \I__4936\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30878\
        );

    \I__4935\ : InMux
    port map (
            O => \N__30884\,
            I => \N__30875\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__30881\,
            I => \N__30872\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__30878\,
            I => \N__30869\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__30875\,
            I => \N__30866\
        );

    \I__4931\ : Odrv4
    port map (
            O => \N__30872\,
            I => n2425
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__30869\,
            I => n2425
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__30866\,
            I => n2425
        );

    \I__4928\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__30856\,
            I => n2492
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__30853\,
            I => \N__30849\
        );

    \I__4925\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30846\
        );

    \I__4924\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30843\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__30846\,
            I => \N__30840\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__30843\,
            I => \N__30837\
        );

    \I__4921\ : Span4Mux_h
    port map (
            O => \N__30840\,
            I => \N__30834\
        );

    \I__4920\ : Odrv4
    port map (
            O => \N__30837\,
            I => n2524
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__30834\,
            I => n2524
        );

    \I__4918\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30826\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__30826\,
            I => n2590
        );

    \I__4916\ : InMux
    port map (
            O => \N__30823\,
            I => \N__30820\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__30820\,
            I => \N__30817\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__30817\,
            I => n2592
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__30814\,
            I => \N__30810\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__30813\,
            I => \N__30807\
        );

    \I__4911\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30804\
        );

    \I__4910\ : InMux
    port map (
            O => \N__30807\,
            I => \N__30801\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__30804\,
            I => \N__30797\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30794\
        );

    \I__4907\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30791\
        );

    \I__4906\ : Odrv4
    port map (
            O => \N__30797\,
            I => n2525
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__30794\,
            I => n2525
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__30791\,
            I => n2525
        );

    \I__4903\ : InMux
    port map (
            O => \N__30784\,
            I => \N__30780\
        );

    \I__4902\ : CascadeMux
    port map (
            O => \N__30783\,
            I => \N__30777\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__30780\,
            I => \N__30774\
        );

    \I__4900\ : InMux
    port map (
            O => \N__30777\,
            I => \N__30771\
        );

    \I__4899\ : Span4Mux_v
    port map (
            O => \N__30774\,
            I => \N__30768\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__30771\,
            I => \N__30765\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__30768\,
            I => n2517
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__30765\,
            I => n2517
        );

    \I__4895\ : InMux
    port map (
            O => \N__30760\,
            I => \N__30757\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__30757\,
            I => n2584
        );

    \I__4893\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30751\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__30751\,
            I => \N__30748\
        );

    \I__4891\ : Odrv4
    port map (
            O => \N__30748\,
            I => n2595
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__30745\,
            I => \N__30741\
        );

    \I__4889\ : CascadeMux
    port map (
            O => \N__30744\,
            I => \N__30738\
        );

    \I__4888\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30735\
        );

    \I__4887\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30732\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__30735\,
            I => \N__30729\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__30732\,
            I => \N__30725\
        );

    \I__4884\ : Span4Mux_h
    port map (
            O => \N__30729\,
            I => \N__30722\
        );

    \I__4883\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30719\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__30725\,
            I => n2528
        );

    \I__4881\ : Odrv4
    port map (
            O => \N__30722\,
            I => n2528
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__30719\,
            I => n2528
        );

    \I__4879\ : InMux
    port map (
            O => \N__30712\,
            I => \N__30709\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__30709\,
            I => n2491
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__30706\,
            I => \N__30703\
        );

    \I__4876\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30700\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__30700\,
            I => \N__30696\
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__30699\,
            I => \N__30693\
        );

    \I__4873\ : Span4Mux_v
    port map (
            O => \N__30696\,
            I => \N__30690\
        );

    \I__4872\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30687\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__30690\,
            I => \N__30682\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__30687\,
            I => \N__30682\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__30682\,
            I => \N__30678\
        );

    \I__4868\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30675\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__30678\,
            I => n2424
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__30675\,
            I => n2424
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__30670\,
            I => \N__30666\
        );

    \I__4864\ : CascadeMux
    port map (
            O => \N__30669\,
            I => \N__30662\
        );

    \I__4863\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30659\
        );

    \I__4862\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30656\
        );

    \I__4861\ : InMux
    port map (
            O => \N__30662\,
            I => \N__30653\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__30659\,
            I => \N__30650\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__30656\,
            I => \N__30647\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__30653\,
            I => n2523
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__30650\,
            I => n2523
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__30647\,
            I => n2523
        );

    \I__4855\ : InMux
    port map (
            O => \N__30640\,
            I => \N__30637\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__30637\,
            I => \N__30634\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__30634\,
            I => \N__30631\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__30631\,
            I => n2583
        );

    \I__4851\ : InMux
    port map (
            O => \N__30628\,
            I => \N__30625\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__30625\,
            I => \N__30622\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__30622\,
            I => n2596
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__30619\,
            I => \N__30615\
        );

    \I__4847\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30612\
        );

    \I__4846\ : InMux
    port map (
            O => \N__30615\,
            I => \N__30609\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__30612\,
            I => \N__30606\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__30609\,
            I => \N__30603\
        );

    \I__4843\ : Span4Mux_h
    port map (
            O => \N__30606\,
            I => \N__30597\
        );

    \I__4842\ : Span4Mux_v
    port map (
            O => \N__30603\,
            I => \N__30597\
        );

    \I__4841\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30594\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__30597\,
            I => n2529
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__30594\,
            I => n2529
        );

    \I__4838\ : InMux
    port map (
            O => \N__30589\,
            I => n12118
        );

    \I__4837\ : InMux
    port map (
            O => \N__30586\,
            I => \N__30583\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__30583\,
            I => n1095
        );

    \I__4835\ : InMux
    port map (
            O => \N__30580\,
            I => n12119
        );

    \I__4834\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30574\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__30574\,
            I => n1094
        );

    \I__4832\ : InMux
    port map (
            O => \N__30571\,
            I => n12120
        );

    \I__4831\ : InMux
    port map (
            O => \N__30568\,
            I => \bfn_6_32_0_\
        );

    \I__4830\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30562\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__30562\,
            I => n1093
        );

    \I__4828\ : CascadeMux
    port map (
            O => \N__30559\,
            I => \N__30556\
        );

    \I__4827\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30553\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__30553\,
            I => n1096
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__30550\,
            I => \N__30547\
        );

    \I__4824\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30544\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__30544\,
            I => \N__30540\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__30543\,
            I => \N__30537\
        );

    \I__4821\ : Span4Mux_s2_h
    port map (
            O => \N__30540\,
            I => \N__30533\
        );

    \I__4820\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30530\
        );

    \I__4819\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30527\
        );

    \I__4818\ : Span4Mux_h
    port map (
            O => \N__30533\,
            I => \N__30524\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__30530\,
            I => n1128
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__30527\,
            I => n1128
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__30524\,
            I => n1128
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__30517\,
            I => \N__30513\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__30516\,
            I => \N__30510\
        );

    \I__4812\ : InMux
    port map (
            O => \N__30513\,
            I => \N__30506\
        );

    \I__4811\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30503\
        );

    \I__4810\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30500\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__30506\,
            I => n1028
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__30503\,
            I => n1028
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__30500\,
            I => n1028
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__30493\,
            I => \N__30489\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__30492\,
            I => \N__30485\
        );

    \I__4804\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30482\
        );

    \I__4803\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30479\
        );

    \I__4802\ : InMux
    port map (
            O => \N__30485\,
            I => \N__30476\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__30482\,
            I => \N__30469\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__30479\,
            I => \N__30469\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__30476\,
            I => \N__30469\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__30469\,
            I => n1027
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__30466\,
            I => \n1059_cascade_\
        );

    \I__4796\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30460\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__30460\,
            I => n1099
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__30457\,
            I => \N__30454\
        );

    \I__4793\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30450\
        );

    \I__4792\ : CascadeMux
    port map (
            O => \N__30453\,
            I => \N__30446\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__30450\,
            I => \N__30443\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__30449\,
            I => \N__30440\
        );

    \I__4789\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30437\
        );

    \I__4788\ : Span4Mux_s1_h
    port map (
            O => \N__30443\,
            I => \N__30434\
        );

    \I__4787\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30431\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__30437\,
            I => \N__30428\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__30434\,
            I => \N__30425\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__30431\,
            I => n1131
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__30428\,
            I => n1131
        );

    \I__4782\ : Odrv4
    port map (
            O => \N__30425\,
            I => n1131
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__30418\,
            I => \N__30414\
        );

    \I__4780\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30411\
        );

    \I__4779\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30408\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30402\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__30408\,
            I => \N__30402\
        );

    \I__4776\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30399\
        );

    \I__4775\ : Span4Mux_v
    port map (
            O => \N__30402\,
            I => \N__30396\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__30399\,
            I => encoder0_position_23
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__30396\,
            I => encoder0_position_23
        );

    \I__4772\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30386\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__30390\,
            I => \N__30383\
        );

    \I__4770\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30380\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__30386\,
            I => \N__30377\
        );

    \I__4768\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30374\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__30380\,
            I => encoder0_position_24
        );

    \I__4766\ : Odrv12
    port map (
            O => \N__30377\,
            I => encoder0_position_24
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__30374\,
            I => encoder0_position_24
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__30367\,
            I => \N__30364\
        );

    \I__4763\ : InMux
    port map (
            O => \N__30364\,
            I => \N__30361\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__30361\,
            I => n1101
        );

    \I__4761\ : InMux
    port map (
            O => \N__30358\,
            I => \bfn_6_31_0_\
        );

    \I__4760\ : InMux
    port map (
            O => \N__30355\,
            I => \N__30352\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__30352\,
            I => n1100
        );

    \I__4758\ : InMux
    port map (
            O => \N__30349\,
            I => n12114
        );

    \I__4757\ : InMux
    port map (
            O => \N__30346\,
            I => n12115
        );

    \I__4756\ : InMux
    port map (
            O => \N__30343\,
            I => \N__30340\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__30340\,
            I => \N__30337\
        );

    \I__4754\ : Span4Mux_s1_v
    port map (
            O => \N__30337\,
            I => \N__30334\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__30334\,
            I => n1098
        );

    \I__4752\ : InMux
    port map (
            O => \N__30331\,
            I => n12116
        );

    \I__4751\ : InMux
    port map (
            O => \N__30328\,
            I => \N__30325\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__30325\,
            I => n1097
        );

    \I__4749\ : InMux
    port map (
            O => \N__30322\,
            I => n12117
        );

    \I__4748\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30314\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__30318\,
            I => \N__30311\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__30317\,
            I => \N__30308\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__30314\,
            I => \N__30304\
        );

    \I__4744\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30301\
        );

    \I__4743\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30298\
        );

    \I__4742\ : InMux
    port map (
            O => \N__30307\,
            I => \N__30295\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__30304\,
            I => n13254
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__30301\,
            I => n13254
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__30298\,
            I => n13254
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__30295\,
            I => n13254
        );

    \I__4737\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30283\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__30283\,
            I => n2286
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__30280\,
            I => \n13255_cascade_\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__30277\,
            I => \N__30273\
        );

    \I__4733\ : InMux
    port map (
            O => \N__30276\,
            I => \N__30268\
        );

    \I__4732\ : InMux
    port map (
            O => \N__30273\,
            I => \N__30263\
        );

    \I__4731\ : InMux
    port map (
            O => \N__30272\,
            I => \N__30263\
        );

    \I__4730\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30260\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30255\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__30263\,
            I => \N__30255\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__30260\,
            I => encoder0_position_26
        );

    \I__4726\ : Odrv4
    port map (
            O => \N__30255\,
            I => encoder0_position_26
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__30250\,
            I => \N__30246\
        );

    \I__4724\ : InMux
    port map (
            O => \N__30249\,
            I => \N__30240\
        );

    \I__4723\ : InMux
    port map (
            O => \N__30246\,
            I => \N__30240\
        );

    \I__4722\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30236\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__30240\,
            I => \N__30233\
        );

    \I__4720\ : InMux
    port map (
            O => \N__30239\,
            I => \N__30230\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__30236\,
            I => encoder0_position_30
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__30233\,
            I => encoder0_position_30
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__30230\,
            I => encoder0_position_30
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__4715\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30217\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__30217\,
            I => n403
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__30214\,
            I => \n11712_cascade_\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__30211\,
            I => \n861_cascade_\
        );

    \I__4711\ : CascadeMux
    port map (
            O => \N__30208\,
            I => \n14170_cascade_\
        );

    \I__4710\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__30202\,
            I => n2285
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__30199\,
            I => \N__30196\
        );

    \I__4707\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__30193\,
            I => n293
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__30190\,
            I => \n293_cascade_\
        );

    \I__4704\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30184\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__30184\,
            I => n5_adj_697
        );

    \I__4702\ : CascadeMux
    port map (
            O => \N__30181\,
            I => \n5_adj_697_cascade_\
        );

    \I__4701\ : InMux
    port map (
            O => \N__30178\,
            I => \N__30175\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__30175\,
            I => n2290
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__30172\,
            I => \n13254_cascade_\
        );

    \I__4698\ : InMux
    port map (
            O => \N__30169\,
            I => \N__30166\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__30166\,
            I => n13259
        );

    \I__4696\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30160\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__30160\,
            I => n13263
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__4693\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30151\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__30151\,
            I => n174
        );

    \I__4691\ : InMux
    port map (
            O => \N__30148\,
            I => \quad_counter0.n12653\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__30145\,
            I => \N__30141\
        );

    \I__4689\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30137\
        );

    \I__4688\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30134\
        );

    \I__4687\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30131\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__30137\,
            I => \N__30128\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__30134\,
            I => encoder0_position_16
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__30131\,
            I => encoder0_position_16
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__30128\,
            I => encoder0_position_16
        );

    \I__4682\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30117\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__30120\,
            I => \N__30113\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__30117\,
            I => \N__30110\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__30116\,
            I => \N__30107\
        );

    \I__4678\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30103\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__30110\,
            I => \N__30100\
        );

    \I__4676\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30097\
        );

    \I__4675\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30094\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__30103\,
            I => encoder0_position_27
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__30100\,
            I => encoder0_position_27
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__30097\,
            I => encoder0_position_27
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__30094\,
            I => encoder0_position_27
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__30085\,
            I => \N__30082\
        );

    \I__4669\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30079\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__30079\,
            I => n175
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__30076\,
            I => \N__30072\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__30075\,
            I => \N__30069\
        );

    \I__4665\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30065\
        );

    \I__4664\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30061\
        );

    \I__4663\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30058\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__30065\,
            I => \N__30055\
        );

    \I__4661\ : InMux
    port map (
            O => \N__30064\,
            I => \N__30052\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__30061\,
            I => encoder0_position_29
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__30058\,
            I => encoder0_position_29
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__30055\,
            I => encoder0_position_29
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__30052\,
            I => encoder0_position_29
        );

    \I__4656\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30040\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__30040\,
            I => n404
        );

    \I__4654\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30030\
        );

    \I__4653\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30030\
        );

    \I__4652\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30027\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__30030\,
            I => \N__30024\
        );

    \I__4650\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30021\
        );

    \I__4649\ : Span4Mux_v
    port map (
            O => \N__30024\,
            I => \N__30018\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__30021\,
            I => encoder0_position_22
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__30018\,
            I => encoder0_position_22
        );

    \I__4646\ : InMux
    port map (
            O => \N__30013\,
            I => \quad_counter0.n12644\
        );

    \I__4645\ : InMux
    port map (
            O => \N__30010\,
            I => \quad_counter0.n12645\
        );

    \I__4644\ : InMux
    port map (
            O => \N__30007\,
            I => \bfn_6_26_0_\
        );

    \I__4643\ : InMux
    port map (
            O => \N__30004\,
            I => \quad_counter0.n12647\
        );

    \I__4642\ : InMux
    port map (
            O => \N__30001\,
            I => \quad_counter0.n12648\
        );

    \I__4641\ : InMux
    port map (
            O => \N__29998\,
            I => \quad_counter0.n12649\
        );

    \I__4640\ : InMux
    port map (
            O => \N__29995\,
            I => \quad_counter0.n12650\
        );

    \I__4639\ : InMux
    port map (
            O => \N__29992\,
            I => \quad_counter0.n12651\
        );

    \I__4638\ : InMux
    port map (
            O => \N__29989\,
            I => \quad_counter0.n12652\
        );

    \I__4637\ : InMux
    port map (
            O => \N__29986\,
            I => \quad_counter0.n12636\
        );

    \I__4636\ : InMux
    port map (
            O => \N__29983\,
            I => \quad_counter0.n12637\
        );

    \I__4635\ : InMux
    port map (
            O => \N__29980\,
            I => \bfn_6_25_0_\
        );

    \I__4634\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29970\
        );

    \I__4633\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29970\
        );

    \I__4632\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29967\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29964\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__29967\,
            I => encoder0_position_17
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__29964\,
            I => encoder0_position_17
        );

    \I__4628\ : InMux
    port map (
            O => \N__29959\,
            I => \quad_counter0.n12639\
        );

    \I__4627\ : CascadeMux
    port map (
            O => \N__29956\,
            I => \N__29952\
        );

    \I__4626\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29948\
        );

    \I__4625\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29945\
        );

    \I__4624\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29942\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__29948\,
            I => \N__29939\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__29945\,
            I => encoder0_position_18
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__29942\,
            I => encoder0_position_18
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__29939\,
            I => encoder0_position_18
        );

    \I__4619\ : InMux
    port map (
            O => \N__29932\,
            I => \quad_counter0.n12640\
        );

    \I__4618\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29923\
        );

    \I__4617\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29923\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__29923\,
            I => \N__29919\
        );

    \I__4615\ : InMux
    port map (
            O => \N__29922\,
            I => \N__29916\
        );

    \I__4614\ : Span4Mux_v
    port map (
            O => \N__29919\,
            I => \N__29913\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__29916\,
            I => encoder0_position_19
        );

    \I__4612\ : Odrv4
    port map (
            O => \N__29913\,
            I => encoder0_position_19
        );

    \I__4611\ : InMux
    port map (
            O => \N__29908\,
            I => \quad_counter0.n12641\
        );

    \I__4610\ : InMux
    port map (
            O => \N__29905\,
            I => \N__29902\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__29902\,
            I => \N__29898\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__29901\,
            I => \N__29894\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__29898\,
            I => \N__29891\
        );

    \I__4606\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29888\
        );

    \I__4605\ : InMux
    port map (
            O => \N__29894\,
            I => \N__29885\
        );

    \I__4604\ : Span4Mux_v
    port map (
            O => \N__29891\,
            I => \N__29880\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29880\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__29885\,
            I => encoder0_position_20
        );

    \I__4601\ : Odrv4
    port map (
            O => \N__29880\,
            I => encoder0_position_20
        );

    \I__4600\ : InMux
    port map (
            O => \N__29875\,
            I => \quad_counter0.n12642\
        );

    \I__4599\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29866\
        );

    \I__4598\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29866\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__29866\,
            I => \N__29862\
        );

    \I__4596\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29859\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__29862\,
            I => \N__29856\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__29859\,
            I => encoder0_position_21
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__29856\,
            I => encoder0_position_21
        );

    \I__4592\ : InMux
    port map (
            O => \N__29851\,
            I => \quad_counter0.n12643\
        );

    \I__4591\ : InMux
    port map (
            O => \N__29848\,
            I => \quad_counter0.n12627\
        );

    \I__4590\ : InMux
    port map (
            O => \N__29845\,
            I => \quad_counter0.n12628\
        );

    \I__4589\ : InMux
    port map (
            O => \N__29842\,
            I => \quad_counter0.n12629\
        );

    \I__4588\ : InMux
    port map (
            O => \N__29839\,
            I => \bfn_6_24_0_\
        );

    \I__4587\ : InMux
    port map (
            O => \N__29836\,
            I => \quad_counter0.n12631\
        );

    \I__4586\ : InMux
    port map (
            O => \N__29833\,
            I => \quad_counter0.n12632\
        );

    \I__4585\ : InMux
    port map (
            O => \N__29830\,
            I => \quad_counter0.n12633\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__29827\,
            I => \N__29823\
        );

    \I__4583\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29820\
        );

    \I__4582\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29816\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29813\
        );

    \I__4580\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29810\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__29816\,
            I => encoder0_position_12
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__29813\,
            I => encoder0_position_12
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__29810\,
            I => encoder0_position_12
        );

    \I__4576\ : InMux
    port map (
            O => \N__29803\,
            I => \quad_counter0.n12634\
        );

    \I__4575\ : InMux
    port map (
            O => \N__29800\,
            I => \quad_counter0.n12635\
        );

    \I__4574\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29794\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__29794\,
            I => \N__29791\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__29791\,
            I => \N__29788\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__29788\,
            I => n2382
        );

    \I__4570\ : CascadeMux
    port map (
            O => \N__29785\,
            I => \n2315_cascade_\
        );

    \I__4569\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29778\
        );

    \I__4568\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29775\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__29778\,
            I => \N__29772\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29767\
        );

    \I__4565\ : Span4Mux_h
    port map (
            O => \N__29772\,
            I => \N__29767\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__29767\,
            I => n2414
        );

    \I__4563\ : CascadeMux
    port map (
            O => \N__29764\,
            I => \n2414_cascade_\
        );

    \I__4562\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29758\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__29758\,
            I => \N__29755\
        );

    \I__4560\ : Odrv4
    port map (
            O => \N__29755\,
            I => n2481
        );

    \I__4559\ : InMux
    port map (
            O => \N__29752\,
            I => \bfn_6_23_0_\
        );

    \I__4558\ : InMux
    port map (
            O => \N__29749\,
            I => \quad_counter0.n12623\
        );

    \I__4557\ : InMux
    port map (
            O => \N__29746\,
            I => \quad_counter0.n12624\
        );

    \I__4556\ : InMux
    port map (
            O => \N__29743\,
            I => \quad_counter0.n12625\
        );

    \I__4555\ : InMux
    port map (
            O => \N__29740\,
            I => \quad_counter0.n12626\
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__29737\,
            I => \n11682_cascade_\
        );

    \I__4553\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29731\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29728\
        );

    \I__4551\ : Odrv4
    port map (
            O => \N__29728\,
            I => n13397
        );

    \I__4550\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29722\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29719\
        );

    \I__4548\ : Odrv12
    port map (
            O => \N__29719\,
            I => n2086
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__29716\,
            I => \N__29713\
        );

    \I__4546\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29709\
        );

    \I__4545\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29706\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__29709\,
            I => \N__29700\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__29706\,
            I => \N__29700\
        );

    \I__4542\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29697\
        );

    \I__4541\ : Odrv12
    port map (
            O => \N__29700\,
            I => n2019
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__29697\,
            I => n2019
        );

    \I__4539\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29688\
        );

    \I__4538\ : InMux
    port map (
            O => \N__29691\,
            I => \N__29685\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__29688\,
            I => \N__29682\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__29685\,
            I => \N__29677\
        );

    \I__4535\ : Span4Mux_s1_h
    port map (
            O => \N__29682\,
            I => \N__29677\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__29677\,
            I => \N__29673\
        );

    \I__4533\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29670\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__29673\,
            I => n2118
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__29670\,
            I => n2118
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__29665\,
            I => \N__29662\
        );

    \I__4529\ : InMux
    port map (
            O => \N__29662\,
            I => \N__29658\
        );

    \I__4528\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29654\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__29658\,
            I => \N__29651\
        );

    \I__4526\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29648\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__29654\,
            I => n2432
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__29651\,
            I => n2432
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__29648\,
            I => n2432
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__29641\,
            I => \N__29638\
        );

    \I__4521\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29635\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__29635\,
            I => \N__29632\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__29632\,
            I => \N__29629\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__29629\,
            I => n2499
        );

    \I__4517\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29622\
        );

    \I__4516\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29619\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__29622\,
            I => \N__29616\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__29619\,
            I => \N__29612\
        );

    \I__4513\ : Span4Mux_v
    port map (
            O => \N__29616\,
            I => \N__29609\
        );

    \I__4512\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29606\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__29612\,
            I => n2025
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__29609\,
            I => n2025
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__29606\,
            I => n2025
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__29599\,
            I => \N__29596\
        );

    \I__4507\ : InMux
    port map (
            O => \N__29596\,
            I => \N__29593\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__29593\,
            I => \N__29590\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__29590\,
            I => \N__29587\
        );

    \I__4504\ : Span4Mux_h
    port map (
            O => \N__29587\,
            I => \N__29584\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__29584\,
            I => n2092
        );

    \I__4502\ : CascadeMux
    port map (
            O => \N__29581\,
            I => \N__29578\
        );

    \I__4501\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29575\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__29575\,
            I => \N__29572\
        );

    \I__4499\ : Span12Mux_s5_h
    port map (
            O => \N__29572\,
            I => \N__29568\
        );

    \I__4498\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29565\
        );

    \I__4497\ : Odrv12
    port map (
            O => \N__29568\,
            I => n2124
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__29565\,
            I => n2124
        );

    \I__4495\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29557\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__29557\,
            I => \N__29554\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__29554\,
            I => \N__29551\
        );

    \I__4492\ : Span4Mux_v
    port map (
            O => \N__29551\,
            I => \N__29548\
        );

    \I__4491\ : Odrv4
    port map (
            O => \N__29548\,
            I => n2191
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__29545\,
            I => \n2124_cascade_\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__29542\,
            I => \n2223_cascade_\
        );

    \I__4488\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29535\
        );

    \I__4487\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29532\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__29535\,
            I => \N__29527\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__29532\,
            I => \N__29527\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__29527\,
            I => \N__29524\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__29524\,
            I => n2315
        );

    \I__4482\ : InMux
    port map (
            O => \N__29521\,
            I => \N__29518\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__29518\,
            I => \N__29515\
        );

    \I__4480\ : Span4Mux_h
    port map (
            O => \N__29515\,
            I => \N__29512\
        );

    \I__4479\ : Span4Mux_h
    port map (
            O => \N__29512\,
            I => \N__29509\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__29509\,
            I => n2192
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__29506\,
            I => \N__29502\
        );

    \I__4476\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29498\
        );

    \I__4475\ : InMux
    port map (
            O => \N__29502\,
            I => \N__29495\
        );

    \I__4474\ : InMux
    port map (
            O => \N__29501\,
            I => \N__29492\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__29498\,
            I => \N__29489\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29486\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__29492\,
            I => \N__29483\
        );

    \I__4470\ : Span4Mux_h
    port map (
            O => \N__29489\,
            I => \N__29480\
        );

    \I__4469\ : Odrv12
    port map (
            O => \N__29486\,
            I => n2125
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__29483\,
            I => n2125
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__29480\,
            I => n2125
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__29473\,
            I => \n2224_cascade_\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__29470\,
            I => \n14174_cascade_\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__29467\,
            I => \n14178_cascade_\
        );

    \I__4463\ : InMux
    port map (
            O => \N__29464\,
            I => \N__29461\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__29461\,
            I => \N__29458\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__29458\,
            I => n14184
        );

    \I__4460\ : InMux
    port map (
            O => \N__29455\,
            I => \N__29452\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__29452\,
            I => \N__29449\
        );

    \I__4458\ : Odrv12
    port map (
            O => \N__29449\,
            I => n2500
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__29446\,
            I => \N__29442\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__29445\,
            I => \N__29439\
        );

    \I__4455\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29436\
        );

    \I__4454\ : InMux
    port map (
            O => \N__29439\,
            I => \N__29433\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__29436\,
            I => \N__29430\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__29433\,
            I => n2433
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__29430\,
            I => n2433
        );

    \I__4450\ : InMux
    port map (
            O => \N__29425\,
            I => \N__29421\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__29424\,
            I => \N__29418\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__29421\,
            I => \N__29415\
        );

    \I__4447\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29412\
        );

    \I__4446\ : Span4Mux_v
    port map (
            O => \N__29415\,
            I => \N__29406\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__29412\,
            I => \N__29406\
        );

    \I__4444\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29403\
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__29406\,
            I => n2431
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__29403\,
            I => n2431
        );

    \I__4441\ : InMux
    port map (
            O => \N__29398\,
            I => \N__29395\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__29395\,
            I => \N__29392\
        );

    \I__4439\ : Odrv4
    port map (
            O => \N__29392\,
            I => n2498
        );

    \I__4438\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29386\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__29386\,
            I => \N__29383\
        );

    \I__4436\ : Span4Mux_h
    port map (
            O => \N__29383\,
            I => \N__29380\
        );

    \I__4435\ : Span4Mux_h
    port map (
            O => \N__29380\,
            I => \N__29377\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__29377\,
            I => n2194
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__29374\,
            I => \N__29371\
        );

    \I__4432\ : InMux
    port map (
            O => \N__29371\,
            I => \N__29367\
        );

    \I__4431\ : InMux
    port map (
            O => \N__29370\,
            I => \N__29363\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__29367\,
            I => \N__29360\
        );

    \I__4429\ : CascadeMux
    port map (
            O => \N__29366\,
            I => \N__29357\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__29363\,
            I => \N__29354\
        );

    \I__4427\ : Span4Mux_h
    port map (
            O => \N__29360\,
            I => \N__29351\
        );

    \I__4426\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29348\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__29354\,
            I => \N__29345\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__29351\,
            I => n2127
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__29348\,
            I => n2127
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__29345\,
            I => n2127
        );

    \I__4421\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29335\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__29335\,
            I => \N__29332\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__29332\,
            I => \N__29329\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__29329\,
            I => n2501
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__29326\,
            I => \n2533_cascade_\
        );

    \I__4416\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29316\
        );

    \I__4415\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29316\
        );

    \I__4414\ : InMux
    port map (
            O => \N__29321\,
            I => \N__29313\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29310\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__29313\,
            I => \N__29307\
        );

    \I__4411\ : Span4Mux_h
    port map (
            O => \N__29310\,
            I => \N__29304\
        );

    \I__4410\ : Odrv12
    port map (
            O => \N__29307\,
            I => n2418
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__29304\,
            I => n2418
        );

    \I__4408\ : InMux
    port map (
            O => \N__29299\,
            I => \N__29296\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__29296\,
            I => n2485
        );

    \I__4406\ : InMux
    port map (
            O => \N__29293\,
            I => \bfn_6_19_0_\
        );

    \I__4405\ : InMux
    port map (
            O => \N__29290\,
            I => n12333
        );

    \I__4404\ : InMux
    port map (
            O => \N__29287\,
            I => n12334
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__29284\,
            I => \N__29281\
        );

    \I__4402\ : InMux
    port map (
            O => \N__29281\,
            I => \N__29276\
        );

    \I__4401\ : InMux
    port map (
            O => \N__29280\,
            I => \N__29273\
        );

    \I__4400\ : InMux
    port map (
            O => \N__29279\,
            I => \N__29270\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__29276\,
            I => n2415
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__29273\,
            I => n2415
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__29270\,
            I => n2415
        );

    \I__4396\ : InMux
    port map (
            O => \N__29263\,
            I => \N__29260\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__29260\,
            I => n2482
        );

    \I__4394\ : InMux
    port map (
            O => \N__29257\,
            I => n12335
        );

    \I__4393\ : InMux
    port map (
            O => \N__29254\,
            I => n12336
        );

    \I__4392\ : InMux
    port map (
            O => \N__29251\,
            I => n12337
        );

    \I__4391\ : InMux
    port map (
            O => \N__29248\,
            I => \N__29244\
        );

    \I__4390\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29241\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__29244\,
            I => \N__29238\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__29241\,
            I => \N__29235\
        );

    \I__4387\ : Span4Mux_h
    port map (
            O => \N__29238\,
            I => \N__29232\
        );

    \I__4386\ : Odrv12
    port map (
            O => \N__29235\,
            I => n2412
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__29232\,
            I => n2412
        );

    \I__4384\ : InMux
    port map (
            O => \N__29227\,
            I => n12338
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__29224\,
            I => \N__29220\
        );

    \I__4382\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29217\
        );

    \I__4381\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29214\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__29217\,
            I => \N__29211\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29208\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__29211\,
            I => \N__29204\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__29208\,
            I => \N__29201\
        );

    \I__4376\ : InMux
    port map (
            O => \N__29207\,
            I => \N__29198\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__29204\,
            I => n2421
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__29201\,
            I => n2421
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__29198\,
            I => n2421
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__29191\,
            I => \N__29188\
        );

    \I__4371\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29185\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__29185\,
            I => n2488
        );

    \I__4369\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29178\
        );

    \I__4368\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29174\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__29178\,
            I => \N__29171\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__29177\,
            I => \N__29168\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29165\
        );

    \I__4364\ : Span4Mux_h
    port map (
            O => \N__29171\,
            I => \N__29162\
        );

    \I__4363\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29159\
        );

    \I__4362\ : Span4Mux_v
    port map (
            O => \N__29165\,
            I => \N__29156\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__29162\,
            I => n2126
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__29159\,
            I => n2126
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__29156\,
            I => n2126
        );

    \I__4358\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29146\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__29146\,
            I => \N__29143\
        );

    \I__4356\ : Span4Mux_h
    port map (
            O => \N__29143\,
            I => \N__29140\
        );

    \I__4355\ : Span4Mux_h
    port map (
            O => \N__29140\,
            I => \N__29137\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__29137\,
            I => n2193
        );

    \I__4353\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29131\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__29131\,
            I => n2493
        );

    \I__4351\ : InMux
    port map (
            O => \N__29128\,
            I => \bfn_6_18_0_\
        );

    \I__4350\ : InMux
    port map (
            O => \N__29125\,
            I => n12325
        );

    \I__4349\ : InMux
    port map (
            O => \N__29122\,
            I => n12326
        );

    \I__4348\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29116\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__29116\,
            I => n2490
        );

    \I__4346\ : InMux
    port map (
            O => \N__29113\,
            I => n12327
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__29110\,
            I => \N__29107\
        );

    \I__4344\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29102\
        );

    \I__4343\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29097\
        );

    \I__4342\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29097\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__29102\,
            I => n2422
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__29097\,
            I => n2422
        );

    \I__4339\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29089\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__29089\,
            I => n2489
        );

    \I__4337\ : InMux
    port map (
            O => \N__29086\,
            I => n12328
        );

    \I__4336\ : InMux
    port map (
            O => \N__29083\,
            I => n12329
        );

    \I__4335\ : InMux
    port map (
            O => \N__29080\,
            I => n12330
        );

    \I__4334\ : InMux
    port map (
            O => \N__29077\,
            I => \N__29074\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__29074\,
            I => \N__29070\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__29073\,
            I => \N__29066\
        );

    \I__4331\ : Span4Mux_h
    port map (
            O => \N__29070\,
            I => \N__29063\
        );

    \I__4330\ : InMux
    port map (
            O => \N__29069\,
            I => \N__29058\
        );

    \I__4329\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29058\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__29063\,
            I => n2419
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__29058\,
            I => n2419
        );

    \I__4326\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29050\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__29050\,
            I => n2486
        );

    \I__4324\ : InMux
    port map (
            O => \N__29047\,
            I => n12331
        );

    \I__4323\ : InMux
    port map (
            O => \N__29044\,
            I => n12361
        );

    \I__4322\ : InMux
    port map (
            O => \N__29041\,
            I => \bfn_6_17_0_\
        );

    \I__4321\ : InMux
    port map (
            O => \N__29038\,
            I => n12317
        );

    \I__4320\ : InMux
    port map (
            O => \N__29035\,
            I => n12318
        );

    \I__4319\ : InMux
    port map (
            O => \N__29032\,
            I => n12319
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__29029\,
            I => \N__29026\
        );

    \I__4317\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29022\
        );

    \I__4316\ : InMux
    port map (
            O => \N__29025\,
            I => \N__29019\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__29015\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__29019\,
            I => \N__29012\
        );

    \I__4313\ : InMux
    port map (
            O => \N__29018\,
            I => \N__29009\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__29015\,
            I => \N__29006\
        );

    \I__4311\ : Span4Mux_v
    port map (
            O => \N__29012\,
            I => \N__29001\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__29009\,
            I => \N__29001\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__29006\,
            I => n2430
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__29001\,
            I => n2430
        );

    \I__4307\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__4305\ : Odrv4
    port map (
            O => \N__28990\,
            I => n2497
        );

    \I__4304\ : InMux
    port map (
            O => \N__28987\,
            I => n12320
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__28984\,
            I => \N__28981\
        );

    \I__4302\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28977\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__28980\,
            I => \N__28974\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__28977\,
            I => \N__28971\
        );

    \I__4299\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28968\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__28971\,
            I => \N__28965\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__28968\,
            I => n2429
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__28965\,
            I => n2429
        );

    \I__4295\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28957\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__28957\,
            I => \N__28954\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__28954\,
            I => n2496
        );

    \I__4292\ : InMux
    port map (
            O => \N__28951\,
            I => n12321
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__28948\,
            I => \N__28945\
        );

    \I__4290\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28942\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28938\
        );

    \I__4288\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28934\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__28938\,
            I => \N__28931\
        );

    \I__4286\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28928\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__28934\,
            I => n2428
        );

    \I__4284\ : Odrv4
    port map (
            O => \N__28931\,
            I => n2428
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__28928\,
            I => n2428
        );

    \I__4282\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28918\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__28918\,
            I => n2495
        );

    \I__4280\ : InMux
    port map (
            O => \N__28915\,
            I => n12322
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__28912\,
            I => \N__28908\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__28911\,
            I => \N__28905\
        );

    \I__4277\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28902\
        );

    \I__4276\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28899\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__28902\,
            I => \N__28896\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__28899\,
            I => \N__28892\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__28896\,
            I => \N__28889\
        );

    \I__4272\ : InMux
    port map (
            O => \N__28895\,
            I => \N__28886\
        );

    \I__4271\ : Span4Mux_v
    port map (
            O => \N__28892\,
            I => \N__28883\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__28889\,
            I => n2427
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__28886\,
            I => n2427
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__28883\,
            I => n2427
        );

    \I__4267\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28873\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__28873\,
            I => n2494
        );

    \I__4265\ : InMux
    port map (
            O => \N__28870\,
            I => n12323
        );

    \I__4264\ : InMux
    port map (
            O => \N__28867\,
            I => n12352
        );

    \I__4263\ : InMux
    port map (
            O => \N__28864\,
            I => n12353
        );

    \I__4262\ : InMux
    port map (
            O => \N__28861\,
            I => \bfn_6_16_0_\
        );

    \I__4261\ : InMux
    port map (
            O => \N__28858\,
            I => n12355
        );

    \I__4260\ : InMux
    port map (
            O => \N__28855\,
            I => n12356
        );

    \I__4259\ : InMux
    port map (
            O => \N__28852\,
            I => n12357
        );

    \I__4258\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__28846\,
            I => n2581
        );

    \I__4256\ : InMux
    port map (
            O => \N__28843\,
            I => n12358
        );

    \I__4255\ : InMux
    port map (
            O => \N__28840\,
            I => n12359
        );

    \I__4254\ : InMux
    port map (
            O => \N__28837\,
            I => n12360
        );

    \I__4253\ : InMux
    port map (
            O => \N__28834\,
            I => n12343
        );

    \I__4252\ : InMux
    port map (
            O => \N__28831\,
            I => n12344
        );

    \I__4251\ : InMux
    port map (
            O => \N__28828\,
            I => n12345
        );

    \I__4250\ : InMux
    port map (
            O => \N__28825\,
            I => \bfn_6_15_0_\
        );

    \I__4249\ : InMux
    port map (
            O => \N__28822\,
            I => n12347
        );

    \I__4248\ : InMux
    port map (
            O => \N__28819\,
            I => n12348
        );

    \I__4247\ : InMux
    port map (
            O => \N__28816\,
            I => n12349
        );

    \I__4246\ : InMux
    port map (
            O => \N__28813\,
            I => n12350
        );

    \I__4245\ : InMux
    port map (
            O => \N__28810\,
            I => n12351
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__28807\,
            I => \N__28804\
        );

    \I__4243\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28801\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28797\
        );

    \I__4241\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28794\
        );

    \I__4240\ : Odrv12
    port map (
            O => \N__28797\,
            I => n1125
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__28794\,
            I => n1125
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__28789\,
            I => \N__28785\
        );

    \I__4237\ : CascadeMux
    port map (
            O => \N__28788\,
            I => \N__28782\
        );

    \I__4236\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28779\
        );

    \I__4235\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28776\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__28779\,
            I => \N__28771\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__28776\,
            I => \N__28771\
        );

    \I__4232\ : Odrv12
    port map (
            O => \N__28771\,
            I => n1126
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__28768\,
            I => \n1126_cascade_\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__28765\,
            I => \N__28762\
        );

    \I__4229\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28759\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__28759\,
            I => \N__28755\
        );

    \I__4227\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28751\
        );

    \I__4226\ : Span4Mux_h
    port map (
            O => \N__28755\,
            I => \N__28748\
        );

    \I__4225\ : InMux
    port map (
            O => \N__28754\,
            I => \N__28745\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__28751\,
            I => n1127
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__28748\,
            I => n1127
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__28745\,
            I => n1127
        );

    \I__4221\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28735\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__28735\,
            I => n13994
        );

    \I__4219\ : InMux
    port map (
            O => \N__28732\,
            I => \bfn_6_14_0_\
        );

    \I__4218\ : InMux
    port map (
            O => \N__28729\,
            I => n12339
        );

    \I__4217\ : InMux
    port map (
            O => \N__28726\,
            I => n12340
        );

    \I__4216\ : InMux
    port map (
            O => \N__28723\,
            I => n12341
        );

    \I__4215\ : InMux
    port map (
            O => \N__28720\,
            I => n12342
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__28717\,
            I => \n1228_cascade_\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__28714\,
            I => \N__28710\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__28713\,
            I => \N__28707\
        );

    \I__4211\ : InMux
    port map (
            O => \N__28710\,
            I => \N__28703\
        );

    \I__4210\ : InMux
    port map (
            O => \N__28707\,
            I => \N__28698\
        );

    \I__4209\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28698\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__28703\,
            I => n1226
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__28698\,
            I => n1226
        );

    \I__4206\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__28690\,
            I => n14078
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__28687\,
            I => \N__28684\
        );

    \I__4203\ : InMux
    port map (
            O => \N__28684\,
            I => \N__28679\
        );

    \I__4202\ : InMux
    port map (
            O => \N__28683\,
            I => \N__28676\
        );

    \I__4201\ : InMux
    port map (
            O => \N__28682\,
            I => \N__28673\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__28679\,
            I => \N__28670\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__28676\,
            I => n1132
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__28673\,
            I => n1132
        );

    \I__4197\ : Odrv12
    port map (
            O => \N__28670\,
            I => n1132
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__28663\,
            I => \N__28660\
        );

    \I__4195\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28656\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__28659\,
            I => \N__28653\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__28656\,
            I => \N__28650\
        );

    \I__4192\ : InMux
    port map (
            O => \N__28653\,
            I => \N__28646\
        );

    \I__4191\ : Span4Mux_s1_h
    port map (
            O => \N__28650\,
            I => \N__28643\
        );

    \I__4190\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28640\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__28646\,
            I => n1129
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__28643\,
            I => n1129
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__28640\,
            I => n1129
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__28633\,
            I => \N__28630\
        );

    \I__4185\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28626\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__28629\,
            I => \N__28623\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__28626\,
            I => \N__28619\
        );

    \I__4182\ : InMux
    port map (
            O => \N__28623\,
            I => \N__28616\
        );

    \I__4181\ : InMux
    port map (
            O => \N__28622\,
            I => \N__28613\
        );

    \I__4180\ : Span4Mux_s1_h
    port map (
            O => \N__28619\,
            I => \N__28610\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__28616\,
            I => n1133
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__28613\,
            I => n1133
        );

    \I__4177\ : Odrv4
    port map (
            O => \N__28610\,
            I => n1133
        );

    \I__4176\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28600\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__28600\,
            I => \N__28597\
        );

    \I__4174\ : Odrv12
    port map (
            O => \N__28597\,
            I => n1195
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__28594\,
            I => \N__28590\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__28593\,
            I => \N__28587\
        );

    \I__4171\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28584\
        );

    \I__4170\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28580\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__28584\,
            I => \N__28577\
        );

    \I__4168\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28574\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__28580\,
            I => n1227
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__28577\,
            I => n1227
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__28574\,
            I => n1227
        );

    \I__4164\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28564\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__28564\,
            I => \N__28561\
        );

    \I__4162\ : Odrv12
    port map (
            O => \N__28561\,
            I => n1198
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__28558\,
            I => \N__28554\
        );

    \I__4160\ : CascadeMux
    port map (
            O => \N__28557\,
            I => \N__28551\
        );

    \I__4159\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28548\
        );

    \I__4158\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28545\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__28548\,
            I => \N__28542\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__28545\,
            I => n1230
        );

    \I__4155\ : Odrv4
    port map (
            O => \N__28542\,
            I => n1230
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__28537\,
            I => \N__28533\
        );

    \I__4153\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28529\
        );

    \I__4152\ : InMux
    port map (
            O => \N__28533\,
            I => \N__28526\
        );

    \I__4151\ : InMux
    port map (
            O => \N__28532\,
            I => \N__28523\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__28529\,
            I => n1229
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__28526\,
            I => n1229
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__28523\,
            I => n1229
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__28516\,
            I => \N__28512\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__28515\,
            I => \N__28508\
        );

    \I__4145\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28505\
        );

    \I__4144\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28502\
        );

    \I__4143\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28499\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__28505\,
            I => n1231
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__28502\,
            I => n1231
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__28499\,
            I => n1231
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__28492\,
            I => \n1230_cascade_\
        );

    \I__4138\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__28486\,
            I => n11642
        );

    \I__4136\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28480\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__28480\,
            I => n13318
        );

    \I__4134\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28474\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28470\
        );

    \I__4132\ : InMux
    port map (
            O => \N__28473\,
            I => \N__28467\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__28470\,
            I => \N__28464\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__28467\,
            I => \N__28461\
        );

    \I__4129\ : IoSpan4Mux
    port map (
            O => \N__28464\,
            I => \N__28458\
        );

    \I__4128\ : Span4Mux_v
    port map (
            O => \N__28461\,
            I => \N__28455\
        );

    \I__4127\ : Odrv4
    port map (
            O => \N__28458\,
            I => \debounce.reg_A_0\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__28455\,
            I => \debounce.reg_A_0\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__28450\,
            I => \N__28447\
        );

    \I__4124\ : InMux
    port map (
            O => \N__28447\,
            I => \N__28443\
        );

    \I__4123\ : InMux
    port map (
            O => \N__28446\,
            I => \N__28440\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__28443\,
            I => \N__28437\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__28440\,
            I => \N__28434\
        );

    \I__4120\ : Span4Mux_s3_v
    port map (
            O => \N__28437\,
            I => \N__28431\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__28434\,
            I => \reg_B_0\
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__28431\,
            I => \reg_B_0\
        );

    \I__4117\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28423\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__28423\,
            I => n2288
        );

    \I__4115\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28417\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__28417\,
            I => \N__28414\
        );

    \I__4113\ : Span4Mux_h
    port map (
            O => \N__28414\,
            I => \N__28411\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__28411\,
            I => n1293
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__28408\,
            I => \N__28405\
        );

    \I__4110\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28401\
        );

    \I__4109\ : InMux
    port map (
            O => \N__28404\,
            I => \N__28398\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__28401\,
            I => \N__28395\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__28398\,
            I => n1325
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__28395\,
            I => n1325
        );

    \I__4105\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28386\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__28389\,
            I => \N__28383\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__28386\,
            I => \N__28379\
        );

    \I__4102\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28376\
        );

    \I__4101\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28373\
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__28379\,
            I => n1326
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__28376\,
            I => n1326
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__28373\,
            I => n1326
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__28366\,
            I => \N__28363\
        );

    \I__4096\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28359\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__28362\,
            I => \N__28356\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__28359\,
            I => \N__28352\
        );

    \I__4093\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28349\
        );

    \I__4092\ : InMux
    port map (
            O => \N__28355\,
            I => \N__28346\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__28352\,
            I => n1327
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__28349\,
            I => n1327
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__28346\,
            I => n1327
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__28339\,
            I => \n1325_cascade_\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__4086\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28330\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__28330\,
            I => \N__28326\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__28329\,
            I => \N__28323\
        );

    \I__4083\ : Span4Mux_s3_h
    port map (
            O => \N__28326\,
            I => \N__28319\
        );

    \I__4082\ : InMux
    port map (
            O => \N__28323\,
            I => \N__28316\
        );

    \I__4081\ : InMux
    port map (
            O => \N__28322\,
            I => \N__28313\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__28319\,
            I => n1328
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__28316\,
            I => n1328
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__28313\,
            I => n1328
        );

    \I__4077\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28303\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__28303\,
            I => n13734
        );

    \I__4075\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28297\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28293\
        );

    \I__4073\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28290\
        );

    \I__4072\ : Span4Mux_s2_v
    port map (
            O => \N__28293\,
            I => \N__28287\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__28290\,
            I => n298
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__28287\,
            I => n298
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__28282\,
            I => \N__28279\
        );

    \I__4068\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28275\
        );

    \I__4067\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28272\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__28275\,
            I => n1233
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__28272\,
            I => n1233
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__28267\,
            I => \n298_cascade_\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__28264\,
            I => \N__28260\
        );

    \I__4062\ : InMux
    port map (
            O => \N__28263\,
            I => \N__28256\
        );

    \I__4061\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28253\
        );

    \I__4060\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28250\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__28256\,
            I => n1232
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__28253\,
            I => n1232
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__28250\,
            I => n1232
        );

    \I__4056\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28240\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28237\
        );

    \I__4054\ : Span4Mux_h
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__28234\,
            I => n1196
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__4051\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28224\
        );

    \I__4050\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28221\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__28224\,
            I => \N__28218\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__28221\,
            I => \N__28213\
        );

    \I__4047\ : Span4Mux_s2_v
    port map (
            O => \N__28218\,
            I => \N__28213\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__28213\,
            I => n1228
        );

    \I__4045\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__28207\,
            I => n2287
        );

    \I__4043\ : InMux
    port map (
            O => \N__28204\,
            I => n12098
        );

    \I__4042\ : InMux
    port map (
            O => \N__28201\,
            I => n12099
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__28198\,
            I => \N__28195\
        );

    \I__4040\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28192\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__28192\,
            I => n402
        );

    \I__4038\ : InMux
    port map (
            O => \N__28189\,
            I => n12100
        );

    \I__4037\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28183\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__28183\,
            I => n2289
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__28180\,
            I => \n13261_cascade_\
        );

    \I__4034\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28173\
        );

    \I__4033\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28170\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__28173\,
            I => \N__28166\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28163\
        );

    \I__4030\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28160\
        );

    \I__4029\ : Span4Mux_s2_v
    port map (
            O => \N__28166\,
            I => \N__28157\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__28163\,
            I => \N__28154\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__28160\,
            I => n297
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__28157\,
            I => n297
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__28154\,
            I => n297
        );

    \I__4024\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28144\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__28144\,
            I => \N__28140\
        );

    \I__4022\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28137\
        );

    \I__4021\ : Span4Mux_v
    port map (
            O => \N__28140\,
            I => \N__28134\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__28137\,
            I => \N__28131\
        );

    \I__4019\ : Span4Mux_h
    port map (
            O => \N__28134\,
            I => \N__28128\
        );

    \I__4018\ : IoSpan4Mux
    port map (
            O => \N__28131\,
            I => \N__28125\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__28128\,
            I => \debounce.reg_A_1\
        );

    \I__4016\ : Odrv4
    port map (
            O => \N__28125\,
            I => \debounce.reg_A_1\
        );

    \I__4015\ : InMux
    port map (
            O => \N__28120\,
            I => \N__28116\
        );

    \I__4014\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28113\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__28116\,
            I => \N__28108\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__28113\,
            I => \N__28108\
        );

    \I__4011\ : Span4Mux_s3_v
    port map (
            O => \N__28108\,
            I => \N__28105\
        );

    \I__4010\ : Odrv4
    port map (
            O => \N__28105\,
            I => \reg_B_1\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__28102\,
            I => \n13257_cascade_\
        );

    \I__4008\ : InMux
    port map (
            O => \N__28099\,
            I => \N__28094\
        );

    \I__4007\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28091\
        );

    \I__4006\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28088\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28085\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__28091\,
            I => \N__28080\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__28088\,
            I => \N__28080\
        );

    \I__4002\ : Span4Mux_v
    port map (
            O => \N__28085\,
            I => \N__28077\
        );

    \I__4001\ : Span4Mux_h
    port map (
            O => \N__28080\,
            I => \N__28074\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__28077\,
            I => n302
        );

    \I__3999\ : Odrv4
    port map (
            O => \N__28074\,
            I => n302
        );

    \I__3998\ : InMux
    port map (
            O => \N__28069\,
            I => \bfn_5_28_0_\
        );

    \I__3997\ : InMux
    port map (
            O => \N__28066\,
            I => n12096
        );

    \I__3996\ : InMux
    port map (
            O => \N__28063\,
            I => n12097
        );

    \I__3995\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28057\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28054\
        );

    \I__3993\ : Span4Mux_v
    port map (
            O => \N__28054\,
            I => \N__28051\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__28051\,
            I => n1801
        );

    \I__3991\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28045\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__28045\,
            I => \N__28040\
        );

    \I__3989\ : InMux
    port map (
            O => \N__28044\,
            I => \N__28037\
        );

    \I__3988\ : InMux
    port map (
            O => \N__28043\,
            I => \N__28034\
        );

    \I__3987\ : Span4Mux_v
    port map (
            O => \N__28040\,
            I => \N__28031\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__28037\,
            I => n303
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__28034\,
            I => n303
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__28031\,
            I => n303
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__28024\,
            I => \N__28021\
        );

    \I__3982\ : InMux
    port map (
            O => \N__28021\,
            I => \N__28016\
        );

    \I__3981\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28013\
        );

    \I__3980\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28010\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__28007\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__28013\,
            I => \N__28004\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__28010\,
            I => \N__27999\
        );

    \I__3976\ : Span4Mux_h
    port map (
            O => \N__28007\,
            I => \N__27999\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__28004\,
            I => n1833
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__27999\,
            I => n1833
        );

    \I__3973\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27990\
        );

    \I__3972\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27987\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__27990\,
            I => \N__27984\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__27987\,
            I => \N__27981\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__27984\,
            I => \N__27978\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__27981\,
            I => \N__27974\
        );

    \I__3967\ : Span4Mux_v
    port map (
            O => \N__27978\,
            I => \N__27971\
        );

    \I__3966\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27968\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__27974\,
            I => \N__27965\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__27971\,
            I => \N__27962\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27959\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__27965\,
            I => n307
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__27962\,
            I => n307
        );

    \I__3960\ : Odrv12
    port map (
            O => \N__27959\,
            I => n307
        );

    \I__3959\ : InMux
    port map (
            O => \N__27952\,
            I => \N__27949\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__27949\,
            I => \N__27946\
        );

    \I__3957\ : Span4Mux_v
    port map (
            O => \N__27946\,
            I => \N__27940\
        );

    \I__3956\ : InMux
    port map (
            O => \N__27945\,
            I => \N__27937\
        );

    \I__3955\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27932\
        );

    \I__3954\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27932\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__27940\,
            I => \N__27925\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27925\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__27932\,
            I => \N__27925\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__27925\,
            I => n13490
        );

    \I__3949\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27918\
        );

    \I__3948\ : InMux
    port map (
            O => \N__27921\,
            I => \N__27915\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__27918\,
            I => \N__27911\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__27915\,
            I => \N__27908\
        );

    \I__3945\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27905\
        );

    \I__3944\ : Span4Mux_v
    port map (
            O => \N__27911\,
            I => \N__27902\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__27908\,
            I => \N__27897\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__27905\,
            I => \N__27897\
        );

    \I__3941\ : Span4Mux_v
    port map (
            O => \N__27902\,
            I => \N__27894\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__27897\,
            I => \N__27891\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__27894\,
            I => n306
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__27891\,
            I => n306
        );

    \I__3937\ : InMux
    port map (
            O => \N__27886\,
            I => \N__27882\
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__27885\,
            I => \N__27879\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__27882\,
            I => \N__27876\
        );

    \I__3934\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27873\
        );

    \I__3933\ : Span4Mux_v
    port map (
            O => \N__27876\,
            I => \N__27867\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__27873\,
            I => \N__27867\
        );

    \I__3931\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27864\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__27867\,
            I => n1726
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__27864\,
            I => n1726
        );

    \I__3928\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27855\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__27858\,
            I => \N__27852\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27849\
        );

    \I__3925\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27846\
        );

    \I__3924\ : Span4Mux_v
    port map (
            O => \N__27849\,
            I => \N__27843\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__27846\,
            I => \N__27840\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__27843\,
            I => n1825
        );

    \I__3921\ : Odrv12
    port map (
            O => \N__27840\,
            I => n1825
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__27835\,
            I => \N__27831\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__27834\,
            I => \N__27828\
        );

    \I__3918\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27825\
        );

    \I__3917\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27822\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__27825\,
            I => \N__27816\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__27822\,
            I => \N__27816\
        );

    \I__3914\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27813\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__27816\,
            I => n1827
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__27813\,
            I => n1827
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__3910\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27802\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__27802\,
            I => \N__27798\
        );

    \I__3908\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27794\
        );

    \I__3907\ : Span4Mux_s3_h
    port map (
            O => \N__27798\,
            I => \N__27791\
        );

    \I__3906\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27788\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__27794\,
            I => n1826
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__27791\,
            I => n1826
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__27788\,
            I => n1826
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__27781\,
            I => \n1825_cascade_\
        );

    \I__3901\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27775\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__27775\,
            I => n14122
        );

    \I__3899\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27768\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__27771\,
            I => \N__27765\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__27768\,
            I => \N__27762\
        );

    \I__3896\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27759\
        );

    \I__3895\ : Span4Mux_h
    port map (
            O => \N__27762\,
            I => \N__27754\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__27759\,
            I => \N__27754\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__27754\,
            I => n1729
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__27751\,
            I => \N__27748\
        );

    \I__3891\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27745\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__27745\,
            I => n1796
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__27742\,
            I => \N__27738\
        );

    \I__3888\ : InMux
    port map (
            O => \N__27741\,
            I => \N__27735\
        );

    \I__3887\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27732\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27729\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__27732\,
            I => \N__27726\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__27729\,
            I => \N__27720\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__27726\,
            I => \N__27720\
        );

    \I__3882\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27717\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__27720\,
            I => n1828
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__27717\,
            I => n1828
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__27712\,
            I => \N__27707\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__27711\,
            I => \N__27704\
        );

    \I__3877\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27701\
        );

    \I__3876\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27698\
        );

    \I__3875\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27695\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__27701\,
            I => \N__27692\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__27698\,
            I => n1832
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__27695\,
            I => n1832
        );

    \I__3871\ : Odrv12
    port map (
            O => \N__27692\,
            I => n1832
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__27685\,
            I => \N__27682\
        );

    \I__3869\ : InMux
    port map (
            O => \N__27682\,
            I => \N__27677\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__27681\,
            I => \N__27674\
        );

    \I__3867\ : InMux
    port map (
            O => \N__27680\,
            I => \N__27671\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__27677\,
            I => \N__27668\
        );

    \I__3865\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27665\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__27671\,
            I => n1831
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__27668\,
            I => n1831
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__27665\,
            I => n1831
        );

    \I__3861\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27655\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__27655\,
            I => n11688
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__27652\,
            I => \N__27648\
        );

    \I__3858\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27645\
        );

    \I__3857\ : InMux
    port map (
            O => \N__27648\,
            I => \N__27642\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__27645\,
            I => \N__27639\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27636\
        );

    \I__3854\ : Span4Mux_v
    port map (
            O => \N__27639\,
            I => \N__27630\
        );

    \I__3853\ : Span4Mux_s1_h
    port map (
            O => \N__27636\,
            I => \N__27630\
        );

    \I__3852\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27627\
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__27630\,
            I => n2021
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__27627\,
            I => n2021
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__27622\,
            I => \N__27619\
        );

    \I__3848\ : InMux
    port map (
            O => \N__27619\,
            I => \N__27616\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__27616\,
            I => \N__27613\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__27613\,
            I => \N__27610\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__27610\,
            I => n2088
        );

    \I__3844\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27603\
        );

    \I__3843\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27600\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__27603\,
            I => \N__27597\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27593\
        );

    \I__3840\ : Span4Mux_v
    port map (
            O => \N__27597\,
            I => \N__27590\
        );

    \I__3839\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27587\
        );

    \I__3838\ : Span4Mux_v
    port map (
            O => \N__27593\,
            I => \N__27582\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__27590\,
            I => \N__27582\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__27587\,
            I => \N__27579\
        );

    \I__3835\ : Odrv4
    port map (
            O => \N__27582\,
            I => n2120
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__27579\,
            I => n2120
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__27574\,
            I => \N__27571\
        );

    \I__3832\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27567\
        );

    \I__3831\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27564\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__27567\,
            I => \N__27558\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__27564\,
            I => \N__27558\
        );

    \I__3828\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27555\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__27558\,
            I => \N__27552\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__27555\,
            I => n301
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__27552\,
            I => n301
        );

    \I__3824\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27544\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27541\
        );

    \I__3822\ : Odrv12
    port map (
            O => \N__27541\,
            I => n1897
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__27538\,
            I => \N__27534\
        );

    \I__3820\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27531\
        );

    \I__3819\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27528\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__27531\,
            I => \N__27525\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27522\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__27525\,
            I => \N__27519\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__27522\,
            I => \N__27516\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__27519\,
            I => n1929
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__27516\,
            I => n1929
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__27511\,
            I => \n1929_cascade_\
        );

    \I__3811\ : InMux
    port map (
            O => \N__27508\,
            I => \N__27505\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__27505\,
            I => n14136
        );

    \I__3809\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27499\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__27499\,
            I => \N__27496\
        );

    \I__3807\ : Odrv12
    port map (
            O => \N__27496\,
            I => n1901
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__27493\,
            I => \N__27490\
        );

    \I__3805\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27486\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__27489\,
            I => \N__27483\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__27486\,
            I => \N__27479\
        );

    \I__3802\ : InMux
    port map (
            O => \N__27483\,
            I => \N__27476\
        );

    \I__3801\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27473\
        );

    \I__3800\ : Span4Mux_h
    port map (
            O => \N__27479\,
            I => \N__27470\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__27476\,
            I => n1933
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__27473\,
            I => n1933
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__27470\,
            I => n1933
        );

    \I__3796\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27460\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__27460\,
            I => \N__27457\
        );

    \I__3794\ : Odrv12
    port map (
            O => \N__27457\,
            I => n1898
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__27454\,
            I => \N__27450\
        );

    \I__3792\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27447\
        );

    \I__3791\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27444\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__27447\,
            I => \N__27439\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27439\
        );

    \I__3788\ : Span4Mux_h
    port map (
            O => \N__27439\,
            I => \N__27435\
        );

    \I__3787\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27432\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__27435\,
            I => n1930
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__27432\,
            I => n1930
        );

    \I__3784\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27424\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__27424\,
            I => \N__27421\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__27418\,
            I => n1885
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__27415\,
            I => \N__27410\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__27414\,
            I => \N__27407\
        );

    \I__3778\ : InMux
    port map (
            O => \N__27413\,
            I => \N__27404\
        );

    \I__3777\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27401\
        );

    \I__3776\ : InMux
    port map (
            O => \N__27407\,
            I => \N__27398\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__27404\,
            I => \N__27395\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__27401\,
            I => \N__27392\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__27398\,
            I => \N__27389\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__27395\,
            I => \N__27386\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__27392\,
            I => n1818
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__27389\,
            I => n1818
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__27386\,
            I => n1818
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__27379\,
            I => \N__27376\
        );

    \I__3767\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27373\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__27373\,
            I => \N__27369\
        );

    \I__3765\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27366\
        );

    \I__3764\ : Odrv4
    port map (
            O => \N__27369\,
            I => n1917
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__27366\,
            I => n1917
        );

    \I__3762\ : InMux
    port map (
            O => \N__27361\,
            I => \N__27358\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__27358\,
            I => n1791
        );

    \I__3760\ : CascadeMux
    port map (
            O => \N__27355\,
            I => \N__27352\
        );

    \I__3759\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27349\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__27349\,
            I => \N__27345\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__27348\,
            I => \N__27342\
        );

    \I__3756\ : Span4Mux_h
    port map (
            O => \N__27345\,
            I => \N__27338\
        );

    \I__3755\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27335\
        );

    \I__3754\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27332\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__27338\,
            I => n1724
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__27335\,
            I => n1724
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__27332\,
            I => n1724
        );

    \I__3750\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27321\
        );

    \I__3749\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27318\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__27321\,
            I => \N__27315\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__27318\,
            I => n1823
        );

    \I__3746\ : Odrv12
    port map (
            O => \N__27315\,
            I => n1823
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__27310\,
            I => \N__27307\
        );

    \I__3744\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27303\
        );

    \I__3743\ : InMux
    port map (
            O => \N__27306\,
            I => \N__27299\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__27303\,
            I => \N__27296\
        );

    \I__3741\ : InMux
    port map (
            O => \N__27302\,
            I => \N__27293\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__27299\,
            I => \N__27290\
        );

    \I__3739\ : Span4Mux_s1_h
    port map (
            O => \N__27296\,
            I => \N__27285\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__27293\,
            I => \N__27285\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__27290\,
            I => n1824
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__27285\,
            I => n1824
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__27280\,
            I => \n1823_cascade_\
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__27277\,
            I => \N__27273\
        );

    \I__3733\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27269\
        );

    \I__3732\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27266\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__27272\,
            I => \N__27263\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__27269\,
            I => \N__27260\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27257\
        );

    \I__3728\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27254\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__27260\,
            I => \N__27251\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__27257\,
            I => n1830
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__27254\,
            I => n1830
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__27251\,
            I => n1830
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__27244\,
            I => \N__27241\
        );

    \I__3722\ : InMux
    port map (
            O => \N__27241\,
            I => \N__27237\
        );

    \I__3721\ : InMux
    port map (
            O => \N__27240\,
            I => \N__27233\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__27237\,
            I => \N__27230\
        );

    \I__3719\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27227\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__27233\,
            I => \N__27224\
        );

    \I__3717\ : Span4Mux_s1_h
    port map (
            O => \N__27230\,
            I => \N__27221\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__27227\,
            I => n1829
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__27224\,
            I => n1829
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__27221\,
            I => n1829
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__27214\,
            I => \n14126_cascade_\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__27211\,
            I => \N__27208\
        );

    \I__3711\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27205\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__27205\,
            I => \N__27202\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__27202\,
            I => n14128
        );

    \I__3708\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27196\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__27196\,
            I => n1793
        );

    \I__3706\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27190\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__27190\,
            I => \N__27187\
        );

    \I__3704\ : Span4Mux_h
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__3703\ : Odrv4
    port map (
            O => \N__27184\,
            I => n2000
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__27181\,
            I => \N__27177\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27174\
        );

    \I__3700\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27171\
        );

    \I__3699\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27168\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__27171\,
            I => \N__27165\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__27168\,
            I => \N__27159\
        );

    \I__3696\ : Span4Mux_h
    port map (
            O => \N__27165\,
            I => \N__27159\
        );

    \I__3695\ : InMux
    port map (
            O => \N__27164\,
            I => \N__27156\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__27159\,
            I => n2032
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__27156\,
            I => n2032
        );

    \I__3692\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27148\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__27148\,
            I => \N__27145\
        );

    \I__3690\ : Span4Mux_h
    port map (
            O => \N__27145\,
            I => \N__27142\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__27142\,
            I => n2091
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__27139\,
            I => \N__27136\
        );

    \I__3687\ : InMux
    port map (
            O => \N__27136\,
            I => \N__27133\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__27133\,
            I => \N__27129\
        );

    \I__3685\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27125\
        );

    \I__3684\ : Span4Mux_s3_h
    port map (
            O => \N__27129\,
            I => \N__27122\
        );

    \I__3683\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27119\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__27125\,
            I => n2024
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__27122\,
            I => n2024
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__27119\,
            I => n2024
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__27112\,
            I => \N__27109\
        );

    \I__3678\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27106\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__27106\,
            I => \N__27102\
        );

    \I__3676\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27099\
        );

    \I__3675\ : Span4Mux_h
    port map (
            O => \N__27102\,
            I => \N__27096\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__27099\,
            I => n2123
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__27096\,
            I => n2123
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__27091\,
            I => \n2123_cascade_\
        );

    \I__3671\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27084\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__27087\,
            I => \N__27081\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__27084\,
            I => \N__27078\
        );

    \I__3668\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27075\
        );

    \I__3667\ : Span4Mux_v
    port map (
            O => \N__27078\,
            I => \N__27072\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__27075\,
            I => n2121
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__27072\,
            I => n2121
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__27067\,
            I => \n13746_cascade_\
        );

    \I__3663\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__27061\,
            I => n13748
        );

    \I__3661\ : InMux
    port map (
            O => \N__27058\,
            I => \N__27054\
        );

    \I__3660\ : InMux
    port map (
            O => \N__27057\,
            I => \N__27050\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__27054\,
            I => \N__27047\
        );

    \I__3658\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27044\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__27050\,
            I => \N__27041\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__27047\,
            I => \N__27038\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__27044\,
            I => n2119
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__27041\,
            I => n2119
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__27038\,
            I => n2119
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__27031\,
            I => \n13754_cascade_\
        );

    \I__3651\ : InMux
    port map (
            O => \N__27028\,
            I => \N__27025\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__27025\,
            I => n13382
        );

    \I__3649\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27019\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__27019\,
            I => \N__27016\
        );

    \I__3647\ : Span4Mux_h
    port map (
            O => \N__27016\,
            I => \N__27013\
        );

    \I__3646\ : Odrv4
    port map (
            O => \N__27013\,
            I => n13760
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__27010\,
            I => \N__27007\
        );

    \I__3644\ : InMux
    port map (
            O => \N__27007\,
            I => \N__27003\
        );

    \I__3643\ : InMux
    port map (
            O => \N__27006\,
            I => \N__27000\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__26997\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26994\
        );

    \I__3640\ : Span4Mux_s2_h
    port map (
            O => \N__26997\,
            I => \N__26991\
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__26994\,
            I => n1822
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__26991\,
            I => n1822
        );

    \I__3637\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26983\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__26983\,
            I => \N__26980\
        );

    \I__3635\ : Span4Mux_h
    port map (
            O => \N__26980\,
            I => \N__26977\
        );

    \I__3634\ : Odrv4
    port map (
            O => \N__26977\,
            I => n1889
        );

    \I__3633\ : InMux
    port map (
            O => \N__26974\,
            I => \N__26970\
        );

    \I__3632\ : InMux
    port map (
            O => \N__26973\,
            I => \N__26967\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__26970\,
            I => \N__26964\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__26967\,
            I => \N__26961\
        );

    \I__3629\ : Span4Mux_v
    port map (
            O => \N__26964\,
            I => \N__26955\
        );

    \I__3628\ : Span4Mux_v
    port map (
            O => \N__26961\,
            I => \N__26955\
        );

    \I__3627\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26952\
        );

    \I__3626\ : Odrv4
    port map (
            O => \N__26955\,
            I => n1921
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__26952\,
            I => n1921
        );

    \I__3624\ : CascadeMux
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__3623\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26941\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__26941\,
            I => \N__26938\
        );

    \I__3621\ : Odrv12
    port map (
            O => \N__26938\,
            I => n1900
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__26935\,
            I => \N__26932\
        );

    \I__3619\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26928\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__26931\,
            I => \N__26925\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26922\
        );

    \I__3616\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26919\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__26922\,
            I => \N__26916\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__26919\,
            I => n1932
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__26916\,
            I => n1932
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__26911\,
            I => \n1932_cascade_\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__26908\,
            I => \N__26905\
        );

    \I__3610\ : InMux
    port map (
            O => \N__26905\,
            I => \N__26901\
        );

    \I__3609\ : InMux
    port map (
            O => \N__26904\,
            I => \N__26897\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__26901\,
            I => \N__26894\
        );

    \I__3607\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26891\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__26897\,
            I => \N__26888\
        );

    \I__3605\ : Span4Mux_v
    port map (
            O => \N__26894\,
            I => \N__26883\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26883\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__26888\,
            I => n1931
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__26883\,
            I => n1931
        );

    \I__3601\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26875\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__26875\,
            I => n11686
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__26872\,
            I => \N__26868\
        );

    \I__3598\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26865\
        );

    \I__3597\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26862\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__26865\,
            I => \N__26856\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__26862\,
            I => \N__26856\
        );

    \I__3594\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26853\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__26856\,
            I => \N__26850\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__26853\,
            I => n2332
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__26850\,
            I => n2332
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__26845\,
            I => \n2333_cascade_\
        );

    \I__3589\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26838\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__26841\,
            I => \N__26835\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__26838\,
            I => \N__26832\
        );

    \I__3586\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26829\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__26832\,
            I => \N__26826\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__26829\,
            I => n2331
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__26826\,
            I => n2331
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__26821\,
            I => \N__26818\
        );

    \I__3581\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26815\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__26815\,
            I => n11766
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__26812\,
            I => \N__26809\
        );

    \I__3578\ : InMux
    port map (
            O => \N__26809\,
            I => \N__26806\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__26806\,
            I => \N__26803\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__26803\,
            I => \N__26800\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__26800\,
            I => n2190
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__26797\,
            I => \N__26794\
        );

    \I__3573\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26790\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__26793\,
            I => \N__26787\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__26790\,
            I => \N__26784\
        );

    \I__3570\ : InMux
    port map (
            O => \N__26787\,
            I => \N__26781\
        );

    \I__3569\ : Span4Mux_h
    port map (
            O => \N__26784\,
            I => \N__26778\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__26781\,
            I => n2133
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__26778\,
            I => n2133
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__26773\,
            I => \N__26770\
        );

    \I__3565\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26766\
        );

    \I__3564\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26763\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__26766\,
            I => \N__26759\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__26763\,
            I => \N__26756\
        );

    \I__3561\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26753\
        );

    \I__3560\ : Span4Mux_s1_h
    port map (
            O => \N__26759\,
            I => \N__26748\
        );

    \I__3559\ : Span4Mux_h
    port map (
            O => \N__26756\,
            I => \N__26748\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__26753\,
            I => n2129
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__26748\,
            I => n2129
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__26743\,
            I => \N__26740\
        );

    \I__3555\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26736\
        );

    \I__3554\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26733\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26729\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__26733\,
            I => \N__26726\
        );

    \I__3551\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26723\
        );

    \I__3550\ : Span4Mux_s3_h
    port map (
            O => \N__26729\,
            I => \N__26718\
        );

    \I__3549\ : Span4Mux_h
    port map (
            O => \N__26726\,
            I => \N__26718\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__26723\,
            I => n2130
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__26718\,
            I => n2130
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__26713\,
            I => \n11616_cascade_\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__26710\,
            I => \N__26706\
        );

    \I__3544\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26703\
        );

    \I__3543\ : InMux
    port map (
            O => \N__26706\,
            I => \N__26700\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__26703\,
            I => \N__26697\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__26700\,
            I => \N__26694\
        );

    \I__3540\ : Span4Mux_h
    port map (
            O => \N__26697\,
            I => \N__26688\
        );

    \I__3539\ : Span4Mux_s3_h
    port map (
            O => \N__26694\,
            I => \N__26688\
        );

    \I__3538\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26685\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__26688\,
            I => n2131
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__26685\,
            I => n2131
        );

    \I__3535\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26677\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26674\
        );

    \I__3533\ : Odrv12
    port map (
            O => \N__26674\,
            I => n2001
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__26671\,
            I => \N__26668\
        );

    \I__3531\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26665\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__26665\,
            I => \N__26662\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__26662\,
            I => \N__26658\
        );

    \I__3528\ : InMux
    port map (
            O => \N__26661\,
            I => \N__26655\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__26658\,
            I => n2033
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__26655\,
            I => n2033
        );

    \I__3525\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26647\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__26647\,
            I => \N__26644\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__26644\,
            I => \N__26641\
        );

    \I__3522\ : Odrv4
    port map (
            O => \N__26641\,
            I => n2100
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__26638\,
            I => \n2033_cascade_\
        );

    \I__3520\ : CascadeMux
    port map (
            O => \N__26635\,
            I => \N__26632\
        );

    \I__3519\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26629\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__26629\,
            I => \N__26626\
        );

    \I__3517\ : Span4Mux_s1_h
    port map (
            O => \N__26626\,
            I => \N__26623\
        );

    \I__3516\ : Span4Mux_v
    port map (
            O => \N__26623\,
            I => \N__26619\
        );

    \I__3515\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26616\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__26619\,
            I => n2132
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__26616\,
            I => n2132
        );

    \I__3512\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26608\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__26608\,
            I => \N__26605\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__26605\,
            I => \N__26602\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__26602\,
            I => n2199
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__26599\,
            I => \n2132_cascade_\
        );

    \I__3507\ : InMux
    port map (
            O => \N__26596\,
            I => \N__26593\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__26593\,
            I => \N__26589\
        );

    \I__3505\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26586\
        );

    \I__3504\ : Odrv4
    port map (
            O => \N__26589\,
            I => n2314
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__26586\,
            I => n2314
        );

    \I__3502\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__26578\,
            I => \N__26575\
        );

    \I__3500\ : Odrv4
    port map (
            O => \N__26575\,
            I => n2381
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__26572\,
            I => \n2314_cascade_\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__26569\,
            I => \n2326_cascade_\
        );

    \I__3497\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26563\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__26563\,
            I => \N__26560\
        );

    \I__3495\ : Span4Mux_h
    port map (
            O => \N__26560\,
            I => \N__26557\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__26557\,
            I => n2393
        );

    \I__3493\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26551\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__26551\,
            I => \N__26548\
        );

    \I__3491\ : Span4Mux_v
    port map (
            O => \N__26548\,
            I => \N__26545\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__26545\,
            I => n2400
        );

    \I__3489\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__26539\,
            I => n14194
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__26536\,
            I => \n2247_cascade_\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__26533\,
            I => \N__26530\
        );

    \I__3485\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26526\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__26529\,
            I => \N__26523\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__26526\,
            I => \N__26520\
        );

    \I__3482\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26517\
        );

    \I__3481\ : Span4Mux_h
    port map (
            O => \N__26520\,
            I => \N__26514\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__26517\,
            I => n2333
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__26514\,
            I => n2333
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__26509\,
            I => \n2517_cascade_\
        );

    \I__3477\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26503\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__26503\,
            I => n13804
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__26500\,
            I => \N__26497\
        );

    \I__3474\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26494\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__26494\,
            I => \N__26491\
        );

    \I__3472\ : Odrv12
    port map (
            O => \N__26491\,
            I => n2185
        );

    \I__3471\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26485\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__26485\,
            I => \N__26482\
        );

    \I__3469\ : Span4Mux_h
    port map (
            O => \N__26482\,
            I => \N__26479\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__26479\,
            I => n2390
        );

    \I__3467\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26473\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__26473\,
            I => \N__26470\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__3464\ : Odrv4
    port map (
            O => \N__26467\,
            I => n2401
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__26464\,
            I => \n2433_cascade_\
        );

    \I__3462\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26458\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__26458\,
            I => n11670
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__26455\,
            I => \N__26452\
        );

    \I__3459\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26449\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26446\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__26446\,
            I => n2383
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__26443\,
            I => \n2527_cascade_\
        );

    \I__3455\ : InMux
    port map (
            O => \N__26440\,
            I => \N__26437\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__26437\,
            I => n13798
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__26434\,
            I => \n13796_cascade_\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__26431\,
            I => \n14354_cascade_\
        );

    \I__3451\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26425\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__26425\,
            I => n14220
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__26422\,
            I => \n14224_cascade_\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__26419\,
            I => \n2445_cascade_\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__26416\,
            I => \n1158_cascade_\
        );

    \I__3446\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26410\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__26410\,
            I => \N__26407\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__26407\,
            I => n1199
        );

    \I__3443\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26401\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__26401\,
            I => \N__26398\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__26398\,
            I => n1197
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__26395\,
            I => \N__26392\
        );

    \I__3439\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26388\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__26391\,
            I => \N__26385\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26382\
        );

    \I__3436\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26379\
        );

    \I__3435\ : Span4Mux_v
    port map (
            O => \N__26382\,
            I => \N__26376\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__26379\,
            I => n1130
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__26376\,
            I => n1130
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__26371\,
            I => \n1130_cascade_\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__26368\,
            I => \N__26365\
        );

    \I__3430\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26362\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__26362\,
            I => n14068
        );

    \I__3428\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26356\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__26356\,
            I => n11706
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__26353\,
            I => \N__26349\
        );

    \I__3425\ : InMux
    port map (
            O => \N__26352\,
            I => \N__26346\
        );

    \I__3424\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26343\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26340\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__26343\,
            I => \N__26335\
        );

    \I__3421\ : Span4Mux_v
    port map (
            O => \N__26340\,
            I => \N__26335\
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__26335\,
            I => n1224
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__26332\,
            I => \n1257_cascade_\
        );

    \I__3418\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__26326\,
            I => \N__26323\
        );

    \I__3416\ : Span4Mux_v
    port map (
            O => \N__26323\,
            I => \N__26320\
        );

    \I__3415\ : Odrv4
    port map (
            O => \N__26320\,
            I => n1201
        );

    \I__3414\ : InMux
    port map (
            O => \N__26317\,
            I => \N__26314\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__26314\,
            I => n1300
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__26311\,
            I => \n1233_cascade_\
        );

    \I__3411\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26304\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__26307\,
            I => \N__26301\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__26304\,
            I => \N__26297\
        );

    \I__3408\ : InMux
    port map (
            O => \N__26301\,
            I => \N__26294\
        );

    \I__3407\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26291\
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__26297\,
            I => n1332
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__26294\,
            I => n1332
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__26291\,
            I => n1332
        );

    \I__3403\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26281\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__26281\,
            I => n1296
        );

    \I__3401\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26275\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__26275\,
            I => \N__26272\
        );

    \I__3399\ : Odrv12
    port map (
            O => \N__26272\,
            I => n1194
        );

    \I__3398\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__3396\ : Odrv12
    port map (
            O => \N__26263\,
            I => n1200
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__26260\,
            I => \N__26257\
        );

    \I__3394\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26253\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__26256\,
            I => \N__26249\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__26253\,
            I => \N__26246\
        );

    \I__3391\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26243\
        );

    \I__3390\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26240\
        );

    \I__3389\ : Span4Mux_h
    port map (
            O => \N__26246\,
            I => \N__26237\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__26243\,
            I => n1225
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__26240\,
            I => n1225
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__26237\,
            I => n1225
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__26230\,
            I => \N__26227\
        );

    \I__3384\ : InMux
    port map (
            O => \N__26227\,
            I => \N__26224\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__26224\,
            I => n1292
        );

    \I__3382\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26217\
        );

    \I__3381\ : InMux
    port map (
            O => \N__26220\,
            I => \N__26213\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__26217\,
            I => \N__26210\
        );

    \I__3379\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26207\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__26213\,
            I => \N__26204\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__26210\,
            I => n1324
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__26207\,
            I => n1324
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__26204\,
            I => n1324
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__26197\,
            I => \n11640_cascade_\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__26194\,
            I => \N__26191\
        );

    \I__3372\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26188\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__26188\,
            I => \N__26184\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__26187\,
            I => \N__26180\
        );

    \I__3369\ : Span4Mux_s2_h
    port map (
            O => \N__26184\,
            I => \N__26177\
        );

    \I__3368\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26174\
        );

    \I__3367\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26171\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__26177\,
            I => n1331
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__26174\,
            I => n1331
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__26171\,
            I => n1331
        );

    \I__3363\ : CascadeMux
    port map (
            O => \N__26164\,
            I => \N__26161\
        );

    \I__3362\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26157\
        );

    \I__3361\ : InMux
    port map (
            O => \N__26160\,
            I => \N__26154\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26149\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__26154\,
            I => \N__26149\
        );

    \I__3358\ : Odrv4
    port map (
            O => \N__26149\,
            I => n1323
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__26146\,
            I => \n13315_cascade_\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__26143\,
            I => \n1356_cascade_\
        );

    \I__3355\ : InMux
    port map (
            O => \N__26140\,
            I => \N__26137\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__26137\,
            I => n1392
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__26134\,
            I => \N__26130\
        );

    \I__3352\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26125\
        );

    \I__3351\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26125\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__26125\,
            I => \N__26122\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__26122\,
            I => \N__26118\
        );

    \I__3348\ : InMux
    port map (
            O => \N__26121\,
            I => \N__26115\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__26118\,
            I => n1424
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__26115\,
            I => n1424
        );

    \I__3345\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26105\
        );

    \I__3344\ : InMux
    port map (
            O => \N__26109\,
            I => \N__26102\
        );

    \I__3343\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26099\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__26105\,
            I => n299
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__26102\,
            I => n299
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__26099\,
            I => n299
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__26092\,
            I => \N__26087\
        );

    \I__3338\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26082\
        );

    \I__3337\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26082\
        );

    \I__3336\ : InMux
    port map (
            O => \N__26087\,
            I => \N__26079\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__26082\,
            I => n1330
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__26079\,
            I => n1330
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__26074\,
            I => \N__26071\
        );

    \I__3332\ : InMux
    port map (
            O => \N__26071\,
            I => \N__26068\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__26068\,
            I => n1397
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__26065\,
            I => \N__26062\
        );

    \I__3329\ : InMux
    port map (
            O => \N__26062\,
            I => \N__26058\
        );

    \I__3328\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26055\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__26058\,
            I => \N__26051\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__26055\,
            I => \N__26048\
        );

    \I__3325\ : InMux
    port map (
            O => \N__26054\,
            I => \N__26045\
        );

    \I__3324\ : Span4Mux_s3_h
    port map (
            O => \N__26051\,
            I => \N__26042\
        );

    \I__3323\ : Span4Mux_s3_h
    port map (
            O => \N__26048\,
            I => \N__26039\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__26045\,
            I => n1429
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__26042\,
            I => n1429
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__26039\,
            I => n1429
        );

    \I__3319\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__26029\,
            I => n1297
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__26026\,
            I => \N__26023\
        );

    \I__3316\ : InMux
    port map (
            O => \N__26023\,
            I => \N__26020\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__26020\,
            I => \N__26015\
        );

    \I__3314\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26012\
        );

    \I__3313\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26009\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__26015\,
            I => n1329
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__26012\,
            I => n1329
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__26009\,
            I => n1329
        );

    \I__3309\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25999\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__25999\,
            I => n1295
        );

    \I__3307\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25993\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__25993\,
            I => n1294
        );

    \I__3305\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25987\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__25987\,
            I => \N__25984\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__25984\,
            I => n1393
        );

    \I__3302\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25978\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__25978\,
            I => \N__25975\
        );

    \I__3300\ : Odrv4
    port map (
            O => \N__25975\,
            I => n1394
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__25972\,
            I => \N__25969\
        );

    \I__3298\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25965\
        );

    \I__3297\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25961\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__25965\,
            I => \N__25958\
        );

    \I__3295\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25955\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__25961\,
            I => n1426
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__25958\,
            I => n1426
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__25955\,
            I => n1426
        );

    \I__3291\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25945\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__25945\,
            I => n1399
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__25942\,
            I => \N__25939\
        );

    \I__3288\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25935\
        );

    \I__3287\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25931\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__25935\,
            I => \N__25928\
        );

    \I__3285\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25925\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__25931\,
            I => \N__25922\
        );

    \I__3283\ : Span4Mux_s3_h
    port map (
            O => \N__25928\,
            I => \N__25919\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__25925\,
            I => n1431
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__25922\,
            I => n1431
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__25919\,
            I => n1431
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__25912\,
            I => \N__25909\
        );

    \I__3278\ : InMux
    port map (
            O => \N__25909\,
            I => \N__25906\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__25906\,
            I => \N__25903\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__25903\,
            I => n1391
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__25900\,
            I => \N__25897\
        );

    \I__3274\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25893\
        );

    \I__3273\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25890\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__25893\,
            I => \N__25887\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__25890\,
            I => n1423
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__25887\,
            I => n1423
        );

    \I__3269\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25878\
        );

    \I__3268\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25875\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__25878\,
            I => \N__25872\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__25875\,
            I => \N__25869\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__25872\,
            I => n1422
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__25869\,
            I => n1422
        );

    \I__3263\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25861\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__25861\,
            I => \N__25858\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__25858\,
            I => n13334
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__25855\,
            I => \n1423_cascade_\
        );

    \I__3259\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25849\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__25849\,
            I => n14094
        );

    \I__3257\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25841\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__25845\,
            I => \N__25838\
        );

    \I__3255\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25835\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25832\
        );

    \I__3253\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25829\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__25835\,
            I => n1425
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__25832\,
            I => n1425
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__25829\,
            I => n1425
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__25822\,
            I => \n1455_cascade_\
        );

    \I__3248\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__25816\,
            I => \N__25813\
        );

    \I__3246\ : Odrv12
    port map (
            O => \N__25813\,
            I => n1492
        );

    \I__3245\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25806\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__25809\,
            I => \N__25803\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__25806\,
            I => \N__25799\
        );

    \I__3242\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25796\
        );

    \I__3241\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25793\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__25799\,
            I => n1524
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__25796\,
            I => n1524
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__25793\,
            I => n1524
        );

    \I__3237\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25783\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__25783\,
            I => \N__25780\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__25780\,
            I => n1301
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__25777\,
            I => \N__25773\
        );

    \I__3233\ : InMux
    port map (
            O => \N__25776\,
            I => \N__25770\
        );

    \I__3232\ : InMux
    port map (
            O => \N__25773\,
            I => \N__25767\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__25770\,
            I => n1333
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__25767\,
            I => n1333
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__25762\,
            I => \n1333_cascade_\
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__25759\,
            I => \N__25756\
        );

    \I__3227\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25753\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25750\
        );

    \I__3225\ : Span4Mux_s3_h
    port map (
            O => \N__25750\,
            I => \N__25747\
        );

    \I__3224\ : Odrv4
    port map (
            O => \N__25747\,
            I => n1592
        );

    \I__3223\ : InMux
    port map (
            O => \N__25744\,
            I => n12172
        );

    \I__3222\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25738\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__25738\,
            I => n1591
        );

    \I__3220\ : InMux
    port map (
            O => \N__25735\,
            I => n12173
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__25732\,
            I => \N__25729\
        );

    \I__3218\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25726\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__25726\,
            I => \N__25721\
        );

    \I__3216\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25718\
        );

    \I__3215\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25715\
        );

    \I__3214\ : Span4Mux_h
    port map (
            O => \N__25721\,
            I => \N__25712\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__25718\,
            I => \N__25709\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__25715\,
            I => n1523
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__25712\,
            I => n1523
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__25709\,
            I => n1523
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__3208\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__25696\,
            I => n1590
        );

    \I__3206\ : InMux
    port map (
            O => \N__25693\,
            I => n12174
        );

    \I__3205\ : InMux
    port map (
            O => \N__25690\,
            I => \N__25686\
        );

    \I__3204\ : InMux
    port map (
            O => \N__25689\,
            I => \N__25683\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__25686\,
            I => n1522
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__25683\,
            I => n1522
        );

    \I__3201\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25675\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__25675\,
            I => n1589
        );

    \I__3199\ : InMux
    port map (
            O => \N__25672\,
            I => n12175
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__25669\,
            I => \N__25666\
        );

    \I__3197\ : InMux
    port map (
            O => \N__25666\,
            I => \N__25663\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__25663\,
            I => \N__25659\
        );

    \I__3195\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25656\
        );

    \I__3194\ : Span4Mux_h
    port map (
            O => \N__25659\,
            I => \N__25653\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__25656\,
            I => \N__25650\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__25653\,
            I => n1521
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__25650\,
            I => n1521
        );

    \I__3190\ : InMux
    port map (
            O => \N__25645\,
            I => n12176
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__3188\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25635\
        );

    \I__3187\ : InMux
    port map (
            O => \N__25638\,
            I => \N__25632\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__25635\,
            I => \N__25629\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25626\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__25629\,
            I => n1620
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__25626\,
            I => n1620
        );

    \I__3182\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25618\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__25618\,
            I => \N__25615\
        );

    \I__3180\ : Span4Mux_v
    port map (
            O => \N__25615\,
            I => \N__25611\
        );

    \I__3179\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25608\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__25611\,
            I => n1427
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__25608\,
            I => n1427
        );

    \I__3176\ : CascadeMux
    port map (
            O => \N__25603\,
            I => \N__25600\
        );

    \I__3175\ : InMux
    port map (
            O => \N__25600\,
            I => \N__25597\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__25597\,
            I => \N__25594\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__25594\,
            I => n1494
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__25591\,
            I => \N__25587\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__25590\,
            I => \N__25584\
        );

    \I__3170\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25580\
        );

    \I__3169\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25577\
        );

    \I__3168\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25574\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__25580\,
            I => n1526
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__25577\,
            I => n1526
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__25574\,
            I => n1526
        );

    \I__3164\ : CascadeMux
    port map (
            O => \N__25567\,
            I => \N__25564\
        );

    \I__3163\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25561\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__25561\,
            I => \N__25558\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__25558\,
            I => n1493
        );

    \I__3160\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25552\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__25552\,
            I => \N__25548\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__25551\,
            I => \N__25545\
        );

    \I__3157\ : Span4Mux_s3_h
    port map (
            O => \N__25548\,
            I => \N__25541\
        );

    \I__3156\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25538\
        );

    \I__3155\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25535\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__25541\,
            I => n1525
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__25538\,
            I => n1525
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__25535\,
            I => n1525
        );

    \I__3151\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25525\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__25525\,
            I => n1396
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__25522\,
            I => \N__25519\
        );

    \I__3148\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25516\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__25516\,
            I => \N__25511\
        );

    \I__3146\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25508\
        );

    \I__3145\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25505\
        );

    \I__3144\ : Span4Mux_v
    port map (
            O => \N__25511\,
            I => \N__25502\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__25508\,
            I => \N__25499\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__25505\,
            I => n1428
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__25502\,
            I => n1428
        );

    \I__3140\ : Odrv12
    port map (
            O => \N__25499\,
            I => n1428
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__25492\,
            I => \N__25489\
        );

    \I__3138\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25484\
        );

    \I__3137\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25479\
        );

    \I__3136\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25479\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__25484\,
            I => n1533
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__25479\,
            I => n1533
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__25474\,
            I => \N__25471\
        );

    \I__3132\ : InMux
    port map (
            O => \N__25471\,
            I => \N__25468\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__25468\,
            I => n1600
        );

    \I__3130\ : InMux
    port map (
            O => \N__25465\,
            I => n12164
        );

    \I__3129\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25458\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__25461\,
            I => \N__25455\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__25458\,
            I => \N__25451\
        );

    \I__3126\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25448\
        );

    \I__3125\ : InMux
    port map (
            O => \N__25454\,
            I => \N__25445\
        );

    \I__3124\ : Span4Mux_s2_h
    port map (
            O => \N__25451\,
            I => \N__25442\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__25448\,
            I => \N__25437\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__25445\,
            I => \N__25437\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__25442\,
            I => n1532
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__25437\,
            I => n1532
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__25432\,
            I => \N__25429\
        );

    \I__3118\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25426\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__25426\,
            I => \N__25423\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__25423\,
            I => n1599
        );

    \I__3115\ : InMux
    port map (
            O => \N__25420\,
            I => n12165
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__25417\,
            I => \N__25413\
        );

    \I__3113\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25410\
        );

    \I__3112\ : InMux
    port map (
            O => \N__25413\,
            I => \N__25407\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__25410\,
            I => n1531
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__25407\,
            I => n1531
        );

    \I__3109\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25399\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__25399\,
            I => \N__25396\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__25396\,
            I => n1598
        );

    \I__3106\ : InMux
    port map (
            O => \N__25393\,
            I => n12166
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__25390\,
            I => \N__25386\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__25389\,
            I => \N__25382\
        );

    \I__3103\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25379\
        );

    \I__3102\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25374\
        );

    \I__3101\ : InMux
    port map (
            O => \N__25382\,
            I => \N__25374\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__25379\,
            I => n1530
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__25374\,
            I => n1530
        );

    \I__3098\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25366\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__25366\,
            I => \N__25363\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__25363\,
            I => n1597
        );

    \I__3095\ : InMux
    port map (
            O => \N__25360\,
            I => n12167
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__25357\,
            I => \N__25354\
        );

    \I__3093\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25349\
        );

    \I__3092\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25344\
        );

    \I__3091\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25344\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__25349\,
            I => n1529
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__25344\,
            I => n1529
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__25339\,
            I => \N__25336\
        );

    \I__3087\ : InMux
    port map (
            O => \N__25336\,
            I => \N__25333\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__25333\,
            I => \N__25330\
        );

    \I__3085\ : Odrv4
    port map (
            O => \N__25330\,
            I => n1596
        );

    \I__3084\ : InMux
    port map (
            O => \N__25327\,
            I => n12168
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__25324\,
            I => \N__25320\
        );

    \I__3082\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25317\
        );

    \I__3081\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25314\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25309\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25309\
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__25309\,
            I => n1528
        );

    \I__3077\ : InMux
    port map (
            O => \N__25306\,
            I => \N__25303\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__25303\,
            I => n1595
        );

    \I__3075\ : InMux
    port map (
            O => \N__25300\,
            I => n12169
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__25297\,
            I => \N__25293\
        );

    \I__3073\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25290\
        );

    \I__3072\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25287\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__25290\,
            I => \N__25283\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__25287\,
            I => \N__25280\
        );

    \I__3069\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25277\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__25283\,
            I => n1527
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__25280\,
            I => n1527
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__25277\,
            I => n1527
        );

    \I__3065\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25267\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__25267\,
            I => \N__25264\
        );

    \I__3063\ : Span4Mux_s2_h
    port map (
            O => \N__25264\,
            I => \N__25261\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__25261\,
            I => n1594
        );

    \I__3061\ : InMux
    port map (
            O => \N__25258\,
            I => n12170
        );

    \I__3060\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__25252\,
            I => n1593
        );

    \I__3058\ : InMux
    port map (
            O => \N__25249\,
            I => \bfn_4_27_0_\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__25246\,
            I => \N__25242\
        );

    \I__3056\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25238\
        );

    \I__3055\ : InMux
    port map (
            O => \N__25242\,
            I => \N__25235\
        );

    \I__3054\ : InMux
    port map (
            O => \N__25241\,
            I => \N__25232\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__25238\,
            I => n1725
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__25235\,
            I => n1725
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__25232\,
            I => n1725
        );

    \I__3050\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25222\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__25222\,
            I => n1792
        );

    \I__3048\ : InMux
    port map (
            O => \N__25219\,
            I => n12199
        );

    \I__3047\ : InMux
    port map (
            O => \N__25216\,
            I => n12200
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__25213\,
            I => \N__25208\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__25212\,
            I => \N__25205\
        );

    \I__3044\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25202\
        );

    \I__3043\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25199\
        );

    \I__3042\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25196\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__25202\,
            I => n1723
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__25199\,
            I => n1723
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__25196\,
            I => n1723
        );

    \I__3038\ : InMux
    port map (
            O => \N__25189\,
            I => \N__25186\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__25186\,
            I => \N__25183\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__25183\,
            I => \N__25180\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__25180\,
            I => n1790
        );

    \I__3034\ : InMux
    port map (
            O => \N__25177\,
            I => n12201
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__25174\,
            I => \N__25170\
        );

    \I__3032\ : InMux
    port map (
            O => \N__25173\,
            I => \N__25166\
        );

    \I__3031\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25163\
        );

    \I__3030\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25160\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__25166\,
            I => n1722
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__25163\,
            I => n1722
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__25160\,
            I => n1722
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__25153\,
            I => \N__25150\
        );

    \I__3025\ : InMux
    port map (
            O => \N__25150\,
            I => \N__25147\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__25147\,
            I => n1789
        );

    \I__3023\ : InMux
    port map (
            O => \N__25144\,
            I => n12202
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__25141\,
            I => \N__25138\
        );

    \I__3021\ : InMux
    port map (
            O => \N__25138\,
            I => \N__25135\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__25135\,
            I => \N__25130\
        );

    \I__3019\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25125\
        );

    \I__3018\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25125\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__25130\,
            I => n1721
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__25125\,
            I => n1721
        );

    \I__3015\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25117\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__25117\,
            I => n1788
        );

    \I__3013\ : InMux
    port map (
            O => \N__25114\,
            I => n12203
        );

    \I__3012\ : InMux
    port map (
            O => \N__25111\,
            I => \N__25108\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__25108\,
            I => \N__25104\
        );

    \I__3010\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25101\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__25104\,
            I => n1720
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__25101\,
            I => n1720
        );

    \I__3007\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25093\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__25093\,
            I => \N__25090\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__25090\,
            I => n1787
        );

    \I__3004\ : InMux
    port map (
            O => \N__25087\,
            I => n12204
        );

    \I__3003\ : InMux
    port map (
            O => \N__25084\,
            I => \N__25081\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25077\
        );

    \I__3001\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25074\
        );

    \I__3000\ : Span4Mux_v
    port map (
            O => \N__25077\,
            I => \N__25069\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__25074\,
            I => \N__25069\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__25069\,
            I => \N__25066\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__25066\,
            I => n1719
        );

    \I__2996\ : InMux
    port map (
            O => \N__25063\,
            I => n12205
        );

    \I__2995\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25057\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__25057\,
            I => \N__25054\
        );

    \I__2993\ : Odrv12
    port map (
            O => \N__25054\,
            I => n1601
        );

    \I__2992\ : InMux
    port map (
            O => \N__25051\,
            I => \bfn_4_26_0_\
        );

    \I__2991\ : InMux
    port map (
            O => \N__25048\,
            I => \N__25045\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__25045\,
            I => \N__25041\
        );

    \I__2989\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25038\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__25041\,
            I => n1733
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__25038\,
            I => n1733
        );

    \I__2986\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25030\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__25027\
        );

    \I__2984\ : Odrv12
    port map (
            O => \N__25027\,
            I => n1800
        );

    \I__2983\ : InMux
    port map (
            O => \N__25024\,
            I => n12191
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__25021\,
            I => \N__25018\
        );

    \I__2981\ : InMux
    port map (
            O => \N__25018\,
            I => \N__25014\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__25017\,
            I => \N__25011\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__25014\,
            I => \N__25008\
        );

    \I__2978\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25005\
        );

    \I__2977\ : Span4Mux_v
    port map (
            O => \N__25008\,
            I => \N__24999\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__24999\
        );

    \I__2975\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24996\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__24999\,
            I => n1732
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__24996\,
            I => n1732
        );

    \I__2972\ : InMux
    port map (
            O => \N__24991\,
            I => \N__24988\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__24988\,
            I => n1799
        );

    \I__2970\ : InMux
    port map (
            O => \N__24985\,
            I => n12192
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__24982\,
            I => \N__24979\
        );

    \I__2968\ : InMux
    port map (
            O => \N__24979\,
            I => \N__24975\
        );

    \I__2967\ : InMux
    port map (
            O => \N__24978\,
            I => \N__24972\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__24975\,
            I => \N__24969\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__24972\,
            I => n1731
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__24969\,
            I => n1731
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__24964\,
            I => \N__24961\
        );

    \I__2962\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24958\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__24958\,
            I => \N__24955\
        );

    \I__2960\ : Span4Mux_s3_h
    port map (
            O => \N__24955\,
            I => \N__24952\
        );

    \I__2959\ : Odrv4
    port map (
            O => \N__24952\,
            I => n1798
        );

    \I__2958\ : InMux
    port map (
            O => \N__24949\,
            I => n12193
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__24946\,
            I => \N__24942\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__24945\,
            I => \N__24939\
        );

    \I__2955\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24936\
        );

    \I__2954\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24933\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__24936\,
            I => \N__24928\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__24933\,
            I => \N__24928\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__24928\,
            I => \N__24924\
        );

    \I__2950\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24921\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__24924\,
            I => n1730
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__24921\,
            I => n1730
        );

    \I__2947\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24913\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__24913\,
            I => n1797
        );

    \I__2945\ : InMux
    port map (
            O => \N__24910\,
            I => n12194
        );

    \I__2944\ : InMux
    port map (
            O => \N__24907\,
            I => n12195
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__24904\,
            I => \N__24900\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__24903\,
            I => \N__24897\
        );

    \I__2941\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24894\
        );

    \I__2940\ : InMux
    port map (
            O => \N__24897\,
            I => \N__24891\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__24894\,
            I => \N__24888\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__24891\,
            I => \N__24885\
        );

    \I__2937\ : Span4Mux_v
    port map (
            O => \N__24888\,
            I => \N__24882\
        );

    \I__2936\ : Span4Mux_h
    port map (
            O => \N__24885\,
            I => \N__24879\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__24882\,
            I => n1728
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__24879\,
            I => n1728
        );

    \I__2933\ : InMux
    port map (
            O => \N__24874\,
            I => \N__24871\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__24871\,
            I => n1795
        );

    \I__2931\ : InMux
    port map (
            O => \N__24868\,
            I => n12196
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__24865\,
            I => \N__24861\
        );

    \I__2929\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24858\
        );

    \I__2928\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24855\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__24858\,
            I => \N__24852\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__24855\,
            I => \N__24849\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__24852\,
            I => \N__24845\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__24849\,
            I => \N__24842\
        );

    \I__2923\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24839\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__24845\,
            I => n1727
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__24842\,
            I => n1727
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__24839\,
            I => n1727
        );

    \I__2919\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24829\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__24829\,
            I => n1794
        );

    \I__2917\ : InMux
    port map (
            O => \N__24826\,
            I => n12197
        );

    \I__2916\ : InMux
    port map (
            O => \N__24823\,
            I => \bfn_4_25_0_\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__24820\,
            I => \n1851_cascade_\
        );

    \I__2914\ : InMux
    port map (
            O => \N__24817\,
            I => \N__24814\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__24814\,
            I => \N__24811\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__24811\,
            I => \N__24808\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__24808\,
            I => n1895
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__24805\,
            I => \N__24802\
        );

    \I__2909\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24799\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__24799\,
            I => \N__24795\
        );

    \I__2907\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24791\
        );

    \I__2906\ : Span4Mux_s3_h
    port map (
            O => \N__24795\,
            I => \N__24788\
        );

    \I__2905\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24785\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__24791\,
            I => n1927
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__24788\,
            I => n1927
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__24785\,
            I => n1927
        );

    \I__2901\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24775\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__24775\,
            I => \N__24772\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__24772\,
            I => \N__24769\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__24769\,
            I => n1890
        );

    \I__2897\ : InMux
    port map (
            O => \N__24766\,
            I => \N__24762\
        );

    \I__2896\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24759\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24754\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__24759\,
            I => \N__24754\
        );

    \I__2893\ : Span4Mux_v
    port map (
            O => \N__24754\,
            I => \N__24751\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__24751\,
            I => n1922
        );

    \I__2891\ : InMux
    port map (
            O => \N__24748\,
            I => \N__24745\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__24745\,
            I => n13772
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__24742\,
            I => \n1922_cascade_\
        );

    \I__2888\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24736\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__24736\,
            I => n13770
        );

    \I__2886\ : InMux
    port map (
            O => \N__24733\,
            I => \N__24730\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__24730\,
            I => \N__24726\
        );

    \I__2884\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24722\
        );

    \I__2883\ : Span4Mux_v
    port map (
            O => \N__24726\,
            I => \N__24719\
        );

    \I__2882\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24716\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__24722\,
            I => \N__24713\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__24719\,
            I => n1920
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__24716\,
            I => n1920
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__24713\,
            I => n1920
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__24706\,
            I => \n13778_cascade_\
        );

    \I__2876\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24700\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__24700\,
            I => n13782
        );

    \I__2874\ : InMux
    port map (
            O => \N__24697\,
            I => \bfn_4_24_0_\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__24694\,
            I => \N__24690\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__24693\,
            I => \N__24687\
        );

    \I__2871\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24683\
        );

    \I__2870\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24680\
        );

    \I__2869\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24677\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__24683\,
            I => n1928
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__24680\,
            I => n1928
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__24677\,
            I => n1928
        );

    \I__2865\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24667\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__24667\,
            I => \N__24664\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__24664\,
            I => n1995
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__24661\,
            I => \N__24657\
        );

    \I__2861\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24654\
        );

    \I__2860\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24651\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__24654\,
            I => \N__24648\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24645\
        );

    \I__2857\ : Span4Mux_v
    port map (
            O => \N__24648\,
            I => \N__24641\
        );

    \I__2856\ : Span4Mux_s3_h
    port map (
            O => \N__24645\,
            I => \N__24638\
        );

    \I__2855\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24635\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__24641\,
            I => n2027
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__24638\,
            I => n2027
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__24635\,
            I => n2027
        );

    \I__2851\ : InMux
    port map (
            O => \N__24628\,
            I => \N__24625\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__24625\,
            I => \N__24621\
        );

    \I__2849\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24617\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__24621\,
            I => \N__24614\
        );

    \I__2847\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24611\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__24617\,
            I => n2023
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__24614\,
            I => n2023
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__24611\,
            I => n2023
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__24604\,
            I => \N__24601\
        );

    \I__2842\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24598\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__24598\,
            I => \N__24595\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__24595\,
            I => n2090
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__24592\,
            I => \N__24589\
        );

    \I__2838\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24585\
        );

    \I__2837\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24582\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24579\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__24582\,
            I => \N__24576\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__24579\,
            I => \N__24573\
        );

    \I__2833\ : Odrv12
    port map (
            O => \N__24576\,
            I => n2122
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__24573\,
            I => n2122
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__24568\,
            I => \N__24565\
        );

    \I__2830\ : InMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__24562\,
            I => \N__24558\
        );

    \I__2828\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24554\
        );

    \I__2827\ : Span4Mux_s2_h
    port map (
            O => \N__24558\,
            I => \N__24551\
        );

    \I__2826\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24548\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__24554\,
            I => n2128
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__24551\,
            I => n2128
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__24548\,
            I => n2128
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__24541\,
            I => \n2122_cascade_\
        );

    \I__2821\ : InMux
    port map (
            O => \N__24538\,
            I => \N__24534\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__24537\,
            I => \N__24531\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__24534\,
            I => \N__24527\
        );

    \I__2818\ : InMux
    port map (
            O => \N__24531\,
            I => \N__24522\
        );

    \I__2817\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24522\
        );

    \I__2816\ : Span4Mux_h
    port map (
            O => \N__24527\,
            I => \N__24519\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__24522\,
            I => n1918
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__24519\,
            I => n1918
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__24514\,
            I => \N__24510\
        );

    \I__2812\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24507\
        );

    \I__2811\ : InMux
    port map (
            O => \N__24510\,
            I => \N__24504\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__24507\,
            I => n1919
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__24504\,
            I => n1919
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__24499\,
            I => \N__24495\
        );

    \I__2807\ : InMux
    port map (
            O => \N__24498\,
            I => \N__24491\
        );

    \I__2806\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24488\
        );

    \I__2805\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24485\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__24491\,
            I => n1926
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__24488\,
            I => n1926
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__24485\,
            I => n1926
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__24478\,
            I => \n1950_cascade_\
        );

    \I__2800\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24472\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__24472\,
            I => \N__24469\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__24469\,
            I => n1993
        );

    \I__2797\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24463\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__24463\,
            I => \N__24460\
        );

    \I__2795\ : Span4Mux_h
    port map (
            O => \N__24460\,
            I => \N__24457\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__24457\,
            I => n1999
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__24454\,
            I => \N__24450\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__24453\,
            I => \N__24447\
        );

    \I__2791\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24444\
        );

    \I__2790\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24441\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24438\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__24441\,
            I => \N__24435\
        );

    \I__2787\ : Span12Mux_s3_h
    port map (
            O => \N__24438\,
            I => \N__24432\
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__24435\,
            I => n2031
        );

    \I__2785\ : Odrv12
    port map (
            O => \N__24432\,
            I => n2031
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__24427\,
            I => \n2031_cascade_\
        );

    \I__2783\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__24421\,
            I => n11680
        );

    \I__2781\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24415\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__24415\,
            I => \N__24412\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__24412\,
            I => n1992
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__24409\,
            I => \N__24405\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__24408\,
            I => \N__24402\
        );

    \I__2776\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24398\
        );

    \I__2775\ : InMux
    port map (
            O => \N__24402\,
            I => \N__24395\
        );

    \I__2774\ : InMux
    port map (
            O => \N__24401\,
            I => \N__24392\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__24398\,
            I => n1925
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__24395\,
            I => n1925
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__24392\,
            I => n1925
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__2769\ : InMux
    port map (
            O => \N__24382\,
            I => \N__24379\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__24379\,
            I => \N__24374\
        );

    \I__2767\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24371\
        );

    \I__2766\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24368\
        );

    \I__2765\ : Span4Mux_s2_h
    port map (
            O => \N__24374\,
            I => \N__24365\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24362\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__24368\,
            I => n1819
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__24365\,
            I => n1819
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__24362\,
            I => n1819
        );

    \I__2760\ : InMux
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__24352\,
            I => n14134
        );

    \I__2758\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24346\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__24346\,
            I => \N__24343\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__24343\,
            I => \N__24340\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__24340\,
            I => n2187
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__24337\,
            I => \n2219_cascade_\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__24334\,
            I => \N__24330\
        );

    \I__2752\ : InMux
    port map (
            O => \N__24333\,
            I => \N__24326\
        );

    \I__2751\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24321\
        );

    \I__2750\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24321\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__24326\,
            I => n2318
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__24321\,
            I => n2318
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__24316\,
            I => \N__24313\
        );

    \I__2746\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24309\
        );

    \I__2745\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24305\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__24309\,
            I => \N__24302\
        );

    \I__2743\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24299\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24294\
        );

    \I__2741\ : Span4Mux_s3_h
    port map (
            O => \N__24302\,
            I => \N__24294\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__24299\,
            I => n2330
        );

    \I__2739\ : Odrv4
    port map (
            O => \N__24294\,
            I => n2330
        );

    \I__2738\ : InMux
    port map (
            O => \N__24289\,
            I => \N__24286\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__24286\,
            I => \N__24283\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__24283\,
            I => \N__24280\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__24280\,
            I => n2099
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__24277\,
            I => \N__24274\
        );

    \I__2733\ : InMux
    port map (
            O => \N__24274\,
            I => \N__24271\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__24271\,
            I => \N__24268\
        );

    \I__2731\ : Span4Mux_h
    port map (
            O => \N__24268\,
            I => \N__24265\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__24265\,
            I => n1997
        );

    \I__2729\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24258\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__24261\,
            I => \N__24255\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__24258\,
            I => \N__24252\
        );

    \I__2726\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24249\
        );

    \I__2725\ : Span4Mux_v
    port map (
            O => \N__24252\,
            I => \N__24246\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__24249\,
            I => n2029
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__24246\,
            I => n2029
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__24241\,
            I => \N__24237\
        );

    \I__2721\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24234\
        );

    \I__2720\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24231\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__24234\,
            I => \N__24228\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__24231\,
            I => \N__24225\
        );

    \I__2717\ : Span4Mux_v
    port map (
            O => \N__24228\,
            I => \N__24219\
        );

    \I__2716\ : Span4Mux_s2_h
    port map (
            O => \N__24225\,
            I => \N__24219\
        );

    \I__2715\ : InMux
    port map (
            O => \N__24224\,
            I => \N__24216\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__24219\,
            I => n2030
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__24216\,
            I => n2030
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__24211\,
            I => \n2029_cascade_\
        );

    \I__2711\ : InMux
    port map (
            O => \N__24208\,
            I => \N__24205\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__24205\,
            I => n14154
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__24202\,
            I => \N__24199\
        );

    \I__2708\ : InMux
    port map (
            O => \N__24199\,
            I => \N__24196\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__24196\,
            I => \N__24193\
        );

    \I__2706\ : Span4Mux_h
    port map (
            O => \N__24193\,
            I => \N__24190\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__24190\,
            I => n1990
        );

    \I__2704\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24184\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__24184\,
            I => \N__24180\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__24183\,
            I => \N__24177\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__24180\,
            I => \N__24174\
        );

    \I__2700\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24171\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__24174\,
            I => n1923
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__24171\,
            I => n1923
        );

    \I__2697\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24162\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__24165\,
            I => \N__24159\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__24162\,
            I => \N__24156\
        );

    \I__2694\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24153\
        );

    \I__2693\ : Span4Mux_v
    port map (
            O => \N__24156\,
            I => \N__24150\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__24153\,
            I => \N__24147\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__24150\,
            I => n2022
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__24147\,
            I => n2022
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__24142\,
            I => \n2022_cascade_\
        );

    \I__2688\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24136\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__24136\,
            I => n14146
        );

    \I__2686\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24130\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__24130\,
            I => n14152
        );

    \I__2684\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24124\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__24124\,
            I => n2384
        );

    \I__2682\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24118\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__24118\,
            I => n2385
        );

    \I__2680\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24112\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__24112\,
            I => n2389
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__24109\,
            I => \N__24105\
        );

    \I__2677\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24101\
        );

    \I__2676\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24096\
        );

    \I__2675\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24096\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__24101\,
            I => n2317
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__24096\,
            I => n2317
        );

    \I__2672\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24088\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__24088\,
            I => \N__24085\
        );

    \I__2670\ : Odrv12
    port map (
            O => \N__24085\,
            I => n14410
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__24082\,
            I => \n11774_cascade_\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__24079\,
            I => \n14188_cascade_\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__24076\,
            I => \n2429_cascade_\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__24073\,
            I => \n14210_cascade_\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__24070\,
            I => \n14214_cascade_\
        );

    \I__2664\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24064\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__24064\,
            I => n13423
        );

    \I__2662\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24058\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__24058\,
            I => n2396
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__24055\,
            I => \N__24050\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__24054\,
            I => \N__24047\
        );

    \I__2658\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24044\
        );

    \I__2657\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24041\
        );

    \I__2656\ : InMux
    port map (
            O => \N__24047\,
            I => \N__24038\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__24044\,
            I => \N__24035\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__24041\,
            I => n2329
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__24038\,
            I => n2329
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__24035\,
            I => n2329
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__24028\,
            I => \n14016_cascade_\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__24025\,
            I => \n14022_cascade_\
        );

    \I__2649\ : InMux
    port map (
            O => \N__24022\,
            I => \N__24019\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__24019\,
            I => \N__24016\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__24016\,
            I => n2395
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__24013\,
            I => \n2346_cascade_\
        );

    \I__2645\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24007\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__24007\,
            I => \N__24004\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__24004\,
            I => n1193
        );

    \I__2642\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23998\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__23998\,
            I => \N__23995\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__23995\,
            I => n2198
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__23992\,
            I => \n2230_cascade_\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__23989\,
            I => \N__23986\
        );

    \I__2637\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23983\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23980\
        );

    \I__2635\ : Span4Mux_h
    port map (
            O => \N__23980\,
            I => \N__23977\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__23977\,
            I => n2189
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__23974\,
            I => \n2221_cascade_\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__23971\,
            I => \n2320_cascade_\
        );

    \I__2631\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23965\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__23965\,
            I => n2387
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__23962\,
            I => \N__23959\
        );

    \I__2628\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23956\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__23956\,
            I => n2399
        );

    \I__2626\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23950\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__23950\,
            I => n2397
        );

    \I__2624\ : InMux
    port map (
            O => \N__23947\,
            I => n12134
        );

    \I__2623\ : InMux
    port map (
            O => \N__23944\,
            I => n12135
        );

    \I__2622\ : InMux
    port map (
            O => \N__23941\,
            I => n12136
        );

    \I__2621\ : InMux
    port map (
            O => \N__23938\,
            I => n12137
        );

    \I__2620\ : InMux
    port map (
            O => \N__23935\,
            I => \bfn_3_32_0_\
        );

    \I__2619\ : InMux
    port map (
            O => \N__23932\,
            I => n12139
        );

    \I__2618\ : InMux
    port map (
            O => \N__23929\,
            I => n12140
        );

    \I__2617\ : InMux
    port map (
            O => \N__23926\,
            I => \N__23920\
        );

    \I__2616\ : InMux
    port map (
            O => \N__23925\,
            I => \N__23920\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__23920\,
            I => \reg_B_2\
        );

    \I__2614\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23914\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__23914\,
            I => \N__23911\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__23911\,
            I => \debounce.n6\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__23908\,
            I => \N__23904\
        );

    \I__2610\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23901\
        );

    \I__2609\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23898\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__23901\,
            I => \N__23893\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__23898\,
            I => \N__23893\
        );

    \I__2606\ : Span4Mux_s2_v
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__23890\,
            I => \debounce.reg_A_2\
        );

    \I__2604\ : SRMux
    port map (
            O => \N__23887\,
            I => \N__23883\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__23886\,
            I => \N__23880\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__23883\,
            I => \N__23877\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__23880\,
            I => \N__23874\
        );

    \I__2600\ : Span4Mux_v
    port map (
            O => \N__23877\,
            I => \N__23869\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__23874\,
            I => \N__23869\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__23869\,
            I => \debounce.cnt_next_9__N_418\
        );

    \I__2597\ : InMux
    port map (
            O => \N__23866\,
            I => n12150
        );

    \I__2596\ : InMux
    port map (
            O => \N__23863\,
            I => n12151
        );

    \I__2595\ : InMux
    port map (
            O => \N__23860\,
            I => \bfn_3_31_0_\
        );

    \I__2594\ : InMux
    port map (
            O => \N__23857\,
            I => n12131
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__23854\,
            I => \N__23851\
        );

    \I__2592\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23848\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__23848\,
            I => n1299
        );

    \I__2590\ : InMux
    port map (
            O => \N__23845\,
            I => n12132
        );

    \I__2589\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__23839\,
            I => n1298
        );

    \I__2587\ : InMux
    port map (
            O => \N__23836\,
            I => n12133
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__23833\,
            I => \N__23830\
        );

    \I__2585\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__23827\,
            I => n1400
        );

    \I__2583\ : InMux
    port map (
            O => \N__23824\,
            I => n12141
        );

    \I__2582\ : InMux
    port map (
            O => \N__23821\,
            I => n12142
        );

    \I__2581\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23815\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23812\
        );

    \I__2579\ : Span4Mux_s2_h
    port map (
            O => \N__23812\,
            I => \N__23809\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__23809\,
            I => n1398
        );

    \I__2577\ : InMux
    port map (
            O => \N__23806\,
            I => n12143
        );

    \I__2576\ : InMux
    port map (
            O => \N__23803\,
            I => n12144
        );

    \I__2575\ : InMux
    port map (
            O => \N__23800\,
            I => n12145
        );

    \I__2574\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23794\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__23794\,
            I => \N__23791\
        );

    \I__2572\ : Span4Mux_s2_h
    port map (
            O => \N__23791\,
            I => \N__23788\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__23788\,
            I => n1395
        );

    \I__2570\ : InMux
    port map (
            O => \N__23785\,
            I => n12146
        );

    \I__2569\ : InMux
    port map (
            O => \N__23782\,
            I => n12147
        );

    \I__2568\ : InMux
    port map (
            O => \N__23779\,
            I => \bfn_3_30_0_\
        );

    \I__2567\ : InMux
    port map (
            O => \N__23776\,
            I => n12149
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__23773\,
            I => \N__23770\
        );

    \I__2565\ : InMux
    port map (
            O => \N__23770\,
            I => \N__23767\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__23767\,
            I => n1495
        );

    \I__2563\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23761\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__23761\,
            I => n1496
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__23758\,
            I => \n1528_cascade_\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__23755\,
            I => \n13978_cascade_\
        );

    \I__2559\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23749\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__23749\,
            I => \N__23746\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__23746\,
            I => n13984
        );

    \I__2556\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23738\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__23742\,
            I => \N__23735\
        );

    \I__2554\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23732\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__23738\,
            I => \N__23729\
        );

    \I__2552\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23726\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__23732\,
            I => \N__23723\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__23729\,
            I => n1432
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__23726\,
            I => n1432
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__23723\,
            I => n1432
        );

    \I__2547\ : InMux
    port map (
            O => \N__23716\,
            I => \N__23713\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__23713\,
            I => \N__23710\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__23710\,
            I => n14088
        );

    \I__2544\ : CascadeMux
    port map (
            O => \N__23707\,
            I => \N__23703\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__23706\,
            I => \N__23700\
        );

    \I__2542\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23697\
        );

    \I__2541\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23694\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__23697\,
            I => \N__23691\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__23694\,
            I => n1433
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__23691\,
            I => n1433
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__23686\,
            I => \n1433_cascade_\
        );

    \I__2536\ : InMux
    port map (
            O => \N__23683\,
            I => \N__23680\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__23680\,
            I => n1500
        );

    \I__2534\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23674\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__23674\,
            I => n1401
        );

    \I__2532\ : InMux
    port map (
            O => \N__23671\,
            I => \bfn_3_29_0_\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__2530\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23660\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__23664\,
            I => \N__23657\
        );

    \I__2528\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23654\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23651\
        );

    \I__2526\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23648\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__23654\,
            I => n1627
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__23651\,
            I => n1627
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__23648\,
            I => n1627
        );

    \I__2522\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23638\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23635\
        );

    \I__2520\ : Span4Mux_h
    port map (
            O => \N__23635\,
            I => \N__23631\
        );

    \I__2519\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23628\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__23631\,
            I => n1430
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__23628\,
            I => n1430
        );

    \I__2516\ : InMux
    port map (
            O => \N__23623\,
            I => \N__23620\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__23620\,
            I => n1497
        );

    \I__2514\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23614\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__23614\,
            I => n1498
        );

    \I__2512\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23608\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__23608\,
            I => \N__23605\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__23605\,
            I => \N__23600\
        );

    \I__2509\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23597\
        );

    \I__2508\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23594\
        );

    \I__2507\ : Span4Mux_s1_h
    port map (
            O => \N__23600\,
            I => \N__23591\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__23597\,
            I => \N__23588\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__23594\,
            I => \N__23585\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__23591\,
            I => n1622
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__23588\,
            I => n1622
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__23585\,
            I => n1622
        );

    \I__2501\ : InMux
    port map (
            O => \N__23578\,
            I => \N__23574\
        );

    \I__2500\ : InMux
    port map (
            O => \N__23577\,
            I => \N__23571\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__23574\,
            I => \N__23568\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__23571\,
            I => \N__23563\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__23568\,
            I => \N__23563\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__23563\,
            I => n300
        );

    \I__2495\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23557\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__23557\,
            I => n1501
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__23554\,
            I => \n300_cascade_\
        );

    \I__2492\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23548\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__23548\,
            I => \N__23545\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__23545\,
            I => n1490
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__23542\,
            I => \n1522_cascade_\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__23539\,
            I => \N__23536\
        );

    \I__2487\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23533\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__23533\,
            I => \N__23528\
        );

    \I__2485\ : InMux
    port map (
            O => \N__23532\,
            I => \N__23525\
        );

    \I__2484\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23522\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__23528\,
            I => \N__23519\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__23525\,
            I => \N__23516\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__23522\,
            I => \N__23513\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__23519\,
            I => n1621
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__23516\,
            I => n1621
        );

    \I__2478\ : Odrv12
    port map (
            O => \N__23513\,
            I => n1621
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__23506\,
            I => \N__23503\
        );

    \I__2476\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23498\
        );

    \I__2475\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23493\
        );

    \I__2474\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23493\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__23498\,
            I => n1626
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__23493\,
            I => n1626
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__23488\,
            I => \N__23485\
        );

    \I__2470\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23482\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23479\
        );

    \I__2468\ : Span4Mux_h
    port map (
            O => \N__23479\,
            I => \N__23476\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__23476\,
            I => n1693
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__23473\,
            I => \N__23469\
        );

    \I__2465\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23466\
        );

    \I__2464\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23463\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__23466\,
            I => \N__23460\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__23463\,
            I => \N__23457\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__23460\,
            I => n1632
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__23457\,
            I => n1632
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__23452\,
            I => \n1632_cascade_\
        );

    \I__2458\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23445\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__23448\,
            I => \N__23442\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__23445\,
            I => \N__23438\
        );

    \I__2455\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23435\
        );

    \I__2454\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23432\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__23438\,
            I => n1633
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__23435\,
            I => n1633
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__23432\,
            I => n1633
        );

    \I__2450\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23422\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__23422\,
            I => n11634
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__23419\,
            I => \N__23416\
        );

    \I__2447\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23413\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__23413\,
            I => \N__23410\
        );

    \I__2445\ : Span4Mux_s2_h
    port map (
            O => \N__23410\,
            I => \N__23405\
        );

    \I__2444\ : InMux
    port map (
            O => \N__23409\,
            I => \N__23400\
        );

    \I__2443\ : InMux
    port map (
            O => \N__23408\,
            I => \N__23400\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__23405\,
            I => n1625
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__23400\,
            I => n1625
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__23395\,
            I => \N__23392\
        );

    \I__2439\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23389\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__23389\,
            I => \N__23384\
        );

    \I__2437\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23381\
        );

    \I__2436\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23378\
        );

    \I__2435\ : Span4Mux_s2_h
    port map (
            O => \N__23384\,
            I => \N__23373\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23373\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__23378\,
            I => n1623
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__23373\,
            I => n1623
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__23368\,
            I => \N__23365\
        );

    \I__2430\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23362\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__23362\,
            I => n1499
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__23359\,
            I => \n1531_cascade_\
        );

    \I__2427\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23353\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__23353\,
            I => n11698
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__23350\,
            I => \n14110_cascade_\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__23347\,
            I => \n1653_cascade_\
        );

    \I__2423\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23341\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__23341\,
            I => \N__23338\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__23338\,
            I => \N__23335\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__23335\,
            I => n1691
        );

    \I__2419\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23329\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__23329\,
            I => n13962
        );

    \I__2417\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23323\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__23323\,
            I => n11694
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__23320\,
            I => \n13968_cascade_\
        );

    \I__2414\ : InMux
    port map (
            O => \N__23317\,
            I => \N__23314\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__23314\,
            I => n14116
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__23311\,
            I => \N__23308\
        );

    \I__2411\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23305\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__23305\,
            I => n13972
        );

    \I__2409\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23299\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__23299\,
            I => \N__23296\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__23296\,
            I => \N__23293\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__23293\,
            I => n1690
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__23290\,
            I => \N__23286\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__23289\,
            I => \N__23283\
        );

    \I__2403\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23279\
        );

    \I__2402\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23276\
        );

    \I__2401\ : InMux
    port map (
            O => \N__23282\,
            I => \N__23273\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__23279\,
            I => n1628
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__23276\,
            I => n1628
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__23273\,
            I => n1628
        );

    \I__2397\ : InMux
    port map (
            O => \N__23266\,
            I => \N__23263\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__23263\,
            I => n14104
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__23260\,
            I => \N__23257\
        );

    \I__2394\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23254\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__23254\,
            I => \N__23250\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__23253\,
            I => \N__23246\
        );

    \I__2391\ : Span4Mux_s2_h
    port map (
            O => \N__23250\,
            I => \N__23243\
        );

    \I__2390\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23238\
        );

    \I__2389\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23238\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__23243\,
            I => n1624
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__23238\,
            I => n1624
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__23233\,
            I => \N__23230\
        );

    \I__2385\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23227\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__23227\,
            I => \N__23224\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__23224\,
            I => \N__23221\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__23221\,
            I => n1692
        );

    \I__2381\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23215\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__23215\,
            I => \N__23212\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__23212\,
            I => n1894
        );

    \I__2378\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23206\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__23206\,
            I => \N__23203\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__23203\,
            I => \N__23200\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__23200\,
            I => n1688
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__23197\,
            I => \n1720_cascade_\
        );

    \I__2373\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23190\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__23193\,
            I => \N__23187\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__23190\,
            I => \N__23184\
        );

    \I__2370\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23181\
        );

    \I__2369\ : Span4Mux_v
    port map (
            O => \N__23184\,
            I => \N__23177\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__23181\,
            I => \N__23174\
        );

    \I__2367\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23171\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__23177\,
            I => n1820
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__23174\,
            I => n1820
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__23171\,
            I => n1820
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__23164\,
            I => \n1752_cascade_\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__23161\,
            I => \N__23157\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__23160\,
            I => \N__23154\
        );

    \I__2360\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23151\
        );

    \I__2359\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23147\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__23151\,
            I => \N__23144\
        );

    \I__2357\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23141\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__23147\,
            I => n1821
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__23144\,
            I => n1821
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__23141\,
            I => n1821
        );

    \I__2353\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23131\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__23131\,
            I => n13343
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__23128\,
            I => \N__23125\
        );

    \I__2350\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23122\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23119\
        );

    \I__2348\ : Span4Mux_h
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__23116\,
            I => n1892
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__23113\,
            I => \N__23109\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__23112\,
            I => \N__23106\
        );

    \I__2344\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23103\
        );

    \I__2343\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23100\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__23103\,
            I => n1924
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__23100\,
            I => n1924
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \n1924_cascade_\
        );

    \I__2339\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23089\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__23089\,
            I => \N__23086\
        );

    \I__2337\ : Span4Mux_h
    port map (
            O => \N__23086\,
            I => \N__23083\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__23083\,
            I => n1893
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__23080\,
            I => \N__23077\
        );

    \I__2334\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__23071\,
            I => \N__23068\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__23068\,
            I => n1891
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__23065\,
            I => \n1923_cascade_\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__23062\,
            I => \N__23059\
        );

    \I__2328\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23056\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__23056\,
            I => \N__23053\
        );

    \I__2326\ : Span4Mux_h
    port map (
            O => \N__23053\,
            I => \N__23050\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__23050\,
            I => n1896
        );

    \I__2324\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23044\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__23041\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__23041\,
            I => n1899
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__23038\,
            I => \n1822_cascade_\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__23035\,
            I => \N__23031\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__23034\,
            I => \N__23028\
        );

    \I__2318\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23025\
        );

    \I__2317\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23022\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23018\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__23022\,
            I => \N__23015\
        );

    \I__2314\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23012\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__23018\,
            I => n2028
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__23015\,
            I => n2028
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__23012\,
            I => n2028
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__23005\,
            I => \N__23002\
        );

    \I__2309\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22999\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__22999\,
            I => n1989
        );

    \I__2307\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22993\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__22993\,
            I => n1998
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__2304\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22984\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__22984\,
            I => n1994
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__22981\,
            I => \N__22977\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__22980\,
            I => \N__22973\
        );

    \I__2300\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22970\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__22976\,
            I => \N__22967\
        );

    \I__2298\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22964\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__22970\,
            I => \N__22961\
        );

    \I__2296\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22958\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__22964\,
            I => n2026
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__22961\,
            I => n2026
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__22958\,
            I => n2026
        );

    \I__2292\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__22948\,
            I => \N__22945\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__22945\,
            I => \N__22942\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__22942\,
            I => n1887
        );

    \I__2288\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22936\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__22936\,
            I => n1986
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__22933\,
            I => \n1919_cascade_\
        );

    \I__2285\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22926\
        );

    \I__2284\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22923\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__22926\,
            I => \N__22919\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__22923\,
            I => \N__22916\
        );

    \I__2281\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22913\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__22919\,
            I => \N__22910\
        );

    \I__2279\ : Span4Mux_s3_h
    port map (
            O => \N__22916\,
            I => \N__22907\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__22913\,
            I => n2018
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__22910\,
            I => n2018
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__22907\,
            I => n2018
        );

    \I__2275\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__22897\,
            I => n1988
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__22894\,
            I => \N__22891\
        );

    \I__2272\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22886\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__22890\,
            I => \N__22883\
        );

    \I__2270\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22880\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__22886\,
            I => \N__22877\
        );

    \I__2268\ : InMux
    port map (
            O => \N__22883\,
            I => \N__22874\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__22880\,
            I => n2020
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__22877\,
            I => n2020
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__22874\,
            I => n2020
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__22867\,
            I => \N__22864\
        );

    \I__2263\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22861\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__22861\,
            I => n1987
        );

    \I__2261\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22855\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__22855\,
            I => n1991
        );

    \I__2259\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22849\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__22849\,
            I => \N__22846\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__22846\,
            I => \N__22843\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__22843\,
            I => n2098
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__22840\,
            I => \N__22837\
        );

    \I__2254\ : InMux
    port map (
            O => \N__22837\,
            I => \N__22834\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__22834\,
            I => n2392
        );

    \I__2252\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22828\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__22828\,
            I => \N__22825\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__22825\,
            I => n2096
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__22822\,
            I => \N__22819\
        );

    \I__2248\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22816\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__22816\,
            I => \N__22813\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__22813\,
            I => \N__22810\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__22810\,
            I => n2197
        );

    \I__2244\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22804\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__22804\,
            I => n1996
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22798\
        );

    \I__2241\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22792\
        );

    \I__2239\ : Span4Mux_h
    port map (
            O => \N__22792\,
            I => \N__22789\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__22789\,
            I => n2196
        );

    \I__2237\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22783\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__22780\,
            I => \N__22777\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__22777\,
            I => n2201
        );

    \I__2233\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22771\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__22771\,
            I => n14160
        );

    \I__2231\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22765\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__22765\,
            I => \N__22762\
        );

    \I__2229\ : Span4Mux_h
    port map (
            O => \N__22762\,
            I => \N__22759\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__22759\,
            I => n2186
        );

    \I__2227\ : InMux
    port map (
            O => \N__22756\,
            I => n12308
        );

    \I__2226\ : InMux
    port map (
            O => \N__22753\,
            I => n12309
        );

    \I__2225\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__22747\,
            I => n2386
        );

    \I__2223\ : InMux
    port map (
            O => \N__22744\,
            I => n12310
        );

    \I__2222\ : InMux
    port map (
            O => \N__22741\,
            I => \bfn_3_19_0_\
        );

    \I__2221\ : InMux
    port map (
            O => \N__22738\,
            I => n12312
        );

    \I__2220\ : InMux
    port map (
            O => \N__22735\,
            I => n12313
        );

    \I__2219\ : InMux
    port map (
            O => \N__22732\,
            I => n12314
        );

    \I__2218\ : InMux
    port map (
            O => \N__22729\,
            I => n12315
        );

    \I__2217\ : InMux
    port map (
            O => \N__22726\,
            I => n12316
        );

    \I__2216\ : InMux
    port map (
            O => \N__22723\,
            I => n12299
        );

    \I__2215\ : InMux
    port map (
            O => \N__22720\,
            I => n12300
        );

    \I__2214\ : InMux
    port map (
            O => \N__22717\,
            I => n12301
        );

    \I__2213\ : InMux
    port map (
            O => \N__22714\,
            I => n12302
        );

    \I__2212\ : InMux
    port map (
            O => \N__22711\,
            I => \bfn_3_18_0_\
        );

    \I__2211\ : InMux
    port map (
            O => \N__22708\,
            I => n12304
        );

    \I__2210\ : InMux
    port map (
            O => \N__22705\,
            I => n12305
        );

    \I__2209\ : InMux
    port map (
            O => \N__22702\,
            I => n12306
        );

    \I__2208\ : InMux
    port map (
            O => \N__22699\,
            I => n12307
        );

    \I__2207\ : InMux
    port map (
            O => \N__22696\,
            I => n12739
        );

    \I__2206\ : InMux
    port map (
            O => \N__22693\,
            I => \bfn_2_32_0_\
        );

    \I__2205\ : InMux
    port map (
            O => \N__22690\,
            I => n12741
        );

    \I__2204\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22683\
        );

    \I__2203\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22680\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22677\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__22680\,
            I => \debounce.cnt_reg_4\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__22677\,
            I => \debounce.cnt_reg_4\
        );

    \I__2199\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22668\
        );

    \I__2198\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22665\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__22668\,
            I => \N__22662\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__22665\,
            I => \debounce.cnt_reg_6\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__22662\,
            I => \debounce.cnt_reg_6\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__2193\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22651\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__22651\,
            I => \N__22647\
        );

    \I__2191\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22644\
        );

    \I__2190\ : Span4Mux_s1_v
    port map (
            O => \N__22647\,
            I => \N__22641\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__22644\,
            I => \debounce.cnt_reg_0\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__22641\,
            I => \debounce.cnt_reg_0\
        );

    \I__2187\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22632\
        );

    \I__2186\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22629\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__22632\,
            I => \N__22626\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__22629\,
            I => \debounce.cnt_reg_7\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__22626\,
            I => \debounce.cnt_reg_7\
        );

    \I__2182\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22618\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__22618\,
            I => \debounce.n13\
        );

    \I__2180\ : InMux
    port map (
            O => \N__22615\,
            I => \bfn_3_17_0_\
        );

    \I__2179\ : InMux
    port map (
            O => \N__22612\,
            I => n12296
        );

    \I__2178\ : InMux
    port map (
            O => \N__22609\,
            I => n12297
        );

    \I__2177\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22603\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__22603\,
            I => n2398
        );

    \I__2175\ : InMux
    port map (
            O => \N__22600\,
            I => n12298
        );

    \I__2174\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__22594\,
            I => n11_adj_663
        );

    \I__2172\ : InMux
    port map (
            O => \N__22591\,
            I => n12731
        );

    \I__2171\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22585\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__22585\,
            I => n10_adj_662
        );

    \I__2169\ : InMux
    port map (
            O => \N__22582\,
            I => \bfn_2_31_0_\
        );

    \I__2168\ : InMux
    port map (
            O => \N__22579\,
            I => \N__22576\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__22576\,
            I => n9_adj_661
        );

    \I__2166\ : InMux
    port map (
            O => \N__22573\,
            I => n12733
        );

    \I__2165\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22567\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__22567\,
            I => n8_adj_660
        );

    \I__2163\ : InMux
    port map (
            O => \N__22564\,
            I => n12734
        );

    \I__2162\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22558\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__22558\,
            I => n7_adj_659
        );

    \I__2160\ : InMux
    port map (
            O => \N__22555\,
            I => n12735
        );

    \I__2159\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22549\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__22549\,
            I => n6_adj_658
        );

    \I__2157\ : InMux
    port map (
            O => \N__22546\,
            I => n12736
        );

    \I__2156\ : InMux
    port map (
            O => \N__22543\,
            I => n12737
        );

    \I__2155\ : InMux
    port map (
            O => \N__22540\,
            I => n12738
        );

    \I__2154\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__22534\,
            I => n20_adj_672
        );

    \I__2152\ : InMux
    port map (
            O => \N__22531\,
            I => n12722
        );

    \I__2151\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22525\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__22525\,
            I => n19_adj_671
        );

    \I__2149\ : InMux
    port map (
            O => \N__22522\,
            I => n12723
        );

    \I__2148\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22516\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__22516\,
            I => n18_adj_670
        );

    \I__2146\ : InMux
    port map (
            O => \N__22513\,
            I => \bfn_2_30_0_\
        );

    \I__2145\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22507\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__22507\,
            I => n17_adj_669
        );

    \I__2143\ : InMux
    port map (
            O => \N__22504\,
            I => n12725
        );

    \I__2142\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22498\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__22498\,
            I => n16_adj_668
        );

    \I__2140\ : InMux
    port map (
            O => \N__22495\,
            I => n12726
        );

    \I__2139\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22489\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__22489\,
            I => n15_adj_667
        );

    \I__2137\ : InMux
    port map (
            O => \N__22486\,
            I => n12727
        );

    \I__2136\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22480\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__22480\,
            I => n14_adj_666
        );

    \I__2134\ : InMux
    port map (
            O => \N__22477\,
            I => n12728
        );

    \I__2133\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22471\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__22471\,
            I => n13_adj_665
        );

    \I__2131\ : InMux
    port map (
            O => \N__22468\,
            I => n12729
        );

    \I__2130\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22462\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__22462\,
            I => n12_adj_664
        );

    \I__2128\ : InMux
    port map (
            O => \N__22459\,
            I => n12730
        );

    \I__2127\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22453\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__22453\,
            I => n1491
        );

    \I__2125\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22447\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__22447\,
            I => n26_adj_678
        );

    \I__2123\ : InMux
    port map (
            O => \N__22444\,
            I => \bfn_2_29_0_\
        );

    \I__2122\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__22438\,
            I => n25_adj_677
        );

    \I__2120\ : InMux
    port map (
            O => \N__22435\,
            I => n12717
        );

    \I__2119\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__22429\,
            I => n24_adj_676
        );

    \I__2117\ : InMux
    port map (
            O => \N__22426\,
            I => n12718
        );

    \I__2116\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22420\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__22420\,
            I => n23_adj_675
        );

    \I__2114\ : InMux
    port map (
            O => \N__22417\,
            I => n12719
        );

    \I__2113\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__22411\,
            I => n22_adj_674
        );

    \I__2111\ : InMux
    port map (
            O => \N__22408\,
            I => n12720
        );

    \I__2110\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22402\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__22402\,
            I => n21_adj_673
        );

    \I__2108\ : InMux
    port map (
            O => \N__22399\,
            I => n12721
        );

    \I__2107\ : InMux
    port map (
            O => \N__22396\,
            I => n12154
        );

    \I__2106\ : InMux
    port map (
            O => \N__22393\,
            I => n12155
        );

    \I__2105\ : InMux
    port map (
            O => \N__22390\,
            I => n12156
        );

    \I__2104\ : InMux
    port map (
            O => \N__22387\,
            I => n12157
        );

    \I__2103\ : InMux
    port map (
            O => \N__22384\,
            I => n12158
        );

    \I__2102\ : InMux
    port map (
            O => \N__22381\,
            I => \bfn_2_28_0_\
        );

    \I__2101\ : InMux
    port map (
            O => \N__22378\,
            I => n12160
        );

    \I__2100\ : InMux
    port map (
            O => \N__22375\,
            I => n12161
        );

    \I__2099\ : InMux
    port map (
            O => \N__22372\,
            I => n12162
        );

    \I__2098\ : InMux
    port map (
            O => \N__22369\,
            I => n12163
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__22366\,
            I => \n13986_cascade_\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__22363\,
            I => \n1554_cascade_\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__22360\,
            I => \N__22356\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__22359\,
            I => \N__22352\
        );

    \I__2093\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22349\
        );

    \I__2092\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22344\
        );

    \I__2091\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22344\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__22349\,
            I => n1629
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__22344\,
            I => n1629
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__2087\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22331\
        );

    \I__2086\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22326\
        );

    \I__2085\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22326\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__22331\,
            I => n1631
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__22326\,
            I => n1631
        );

    \I__2082\ : InMux
    port map (
            O => \N__22321\,
            I => \bfn_2_27_0_\
        );

    \I__2081\ : InMux
    port map (
            O => \N__22318\,
            I => n12152
        );

    \I__2080\ : InMux
    port map (
            O => \N__22315\,
            I => n12153
        );

    \I__2079\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22309\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__22309\,
            I => n1698
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__22306\,
            I => \N__22303\
        );

    \I__2076\ : InMux
    port map (
            O => \N__22303\,
            I => \N__22300\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__22300\,
            I => n1696
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__22297\,
            I => \n1728_cascade_\
        );

    \I__2073\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22291\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__22291\,
            I => n1695
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__22288\,
            I => \N__22285\
        );

    \I__2070\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22282\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__22282\,
            I => n1694
        );

    \I__2068\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22276\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__22276\,
            I => \N__22273\
        );

    \I__2066\ : Span4Mux_h
    port map (
            O => \N__22273\,
            I => \N__22270\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__22270\,
            I => n1689
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__22267\,
            I => \N__22264\
        );

    \I__2063\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22260\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__22263\,
            I => \N__22257\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__22260\,
            I => \N__22253\
        );

    \I__2060\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22250\
        );

    \I__2059\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22247\
        );

    \I__2058\ : Odrv12
    port map (
            O => \N__22253\,
            I => n1630
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__22250\,
            I => n1630
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__22247\,
            I => n1630
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__2054\ : InMux
    port map (
            O => \N__22237\,
            I => \N__22234\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__22234\,
            I => \N__22231\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__22231\,
            I => n1700
        );

    \I__2051\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22225\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__22225\,
            I => \N__22222\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__22222\,
            I => n1699
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__22219\,
            I => \n1731_cascade_\
        );

    \I__2047\ : InMux
    port map (
            O => \N__22216\,
            I => \N__22213\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__22213\,
            I => \N__22210\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__22210\,
            I => n1697
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__22207\,
            I => \n1729_cascade_\
        );

    \I__2043\ : InMux
    port map (
            O => \N__22204\,
            I => \N__22201\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__22201\,
            I => \N__22198\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__22198\,
            I => n1701
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__22195\,
            I => \n1733_cascade_\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__22192\,
            I => \N__22189\
        );

    \I__2038\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22186\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__22186\,
            I => n1886
        );

    \I__2036\ : InMux
    port map (
            O => \N__22183\,
            I => n12233
        );

    \I__2035\ : InMux
    port map (
            O => \N__22180\,
            I => n12234
        );

    \I__2034\ : InMux
    port map (
            O => \N__22177\,
            I => n12235
        );

    \I__2033\ : InMux
    port map (
            O => \N__22174\,
            I => n12236
        );

    \I__2032\ : InMux
    port map (
            O => \N__22171\,
            I => \bfn_2_23_0_\
        );

    \I__2031\ : InMux
    port map (
            O => \N__22168\,
            I => n12238
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__22165\,
            I => \N__22162\
        );

    \I__2029\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22159\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__22159\,
            I => \N__22155\
        );

    \I__2027\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22152\
        );

    \I__2026\ : Span4Mux_s2_h
    port map (
            O => \N__22155\,
            I => \N__22149\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__22152\,
            I => n2016
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__22149\,
            I => n2016
        );

    \I__2023\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__22141\,
            I => n1888
        );

    \I__2021\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__22135\,
            I => n1985
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__2018\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22126\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__22126\,
            I => \N__22122\
        );

    \I__2016\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22118\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__22122\,
            I => \N__22115\
        );

    \I__2014\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22112\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__22118\,
            I => \N__22109\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__22115\,
            I => n2017
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__22112\,
            I => n2017
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__22109\,
            I => n2017
        );

    \I__2009\ : InMux
    port map (
            O => \N__22102\,
            I => n12223
        );

    \I__2008\ : InMux
    port map (
            O => \N__22099\,
            I => n12224
        );

    \I__2007\ : InMux
    port map (
            O => \N__22096\,
            I => n12225
        );

    \I__2006\ : InMux
    port map (
            O => \N__22093\,
            I => n12226
        );

    \I__2005\ : InMux
    port map (
            O => \N__22090\,
            I => n12227
        );

    \I__2004\ : InMux
    port map (
            O => \N__22087\,
            I => n12228
        );

    \I__2003\ : InMux
    port map (
            O => \N__22084\,
            I => \bfn_2_22_0_\
        );

    \I__2002\ : InMux
    port map (
            O => \N__22081\,
            I => n12230
        );

    \I__2001\ : InMux
    port map (
            O => \N__22078\,
            I => n12231
        );

    \I__2000\ : InMux
    port map (
            O => \N__22075\,
            I => n12232
        );

    \I__1999\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22069\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__22069\,
            I => \N__22066\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__22066\,
            I => n2084
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__1995\ : InMux
    port map (
            O => \N__22060\,
            I => \N__22056\
        );

    \I__1994\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22053\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__22056\,
            I => n2116
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__22053\,
            I => n2116
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__22048\,
            I => \N__22045\
        );

    \I__1990\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22041\
        );

    \I__1989\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22038\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__22041\,
            I => \N__22033\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__22033\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__22033\,
            I => n2115
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \n2116_cascade_\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__22027\,
            I => \n2148_cascade_\
        );

    \I__1983\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__22018\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__22018\,
            I => n2195
        );

    \I__1980\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22012\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__22012\,
            I => n2087
        );

    \I__1978\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__22006\,
            I => n2093
        );

    \I__1976\ : InMux
    port map (
            O => \N__22003\,
            I => \N__22000\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__21997\,
            I => \N__21994\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__21994\,
            I => n2085
        );

    \I__1972\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21986\
        );

    \I__1971\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21981\
        );

    \I__1970\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21981\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__21986\,
            I => n2117
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__21981\,
            I => n2117
        );

    \I__1967\ : InMux
    port map (
            O => \N__21976\,
            I => \bfn_2_21_0_\
        );

    \I__1966\ : InMux
    port map (
            O => \N__21973\,
            I => n12222
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__21970\,
            I => \n2331_cascade_\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__21967\,
            I => \N__21964\
        );

    \I__1963\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21961\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__21961\,
            I => \N__21958\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__21958\,
            I => n2089
        );

    \I__1960\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21952\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__21952\,
            I => n2188
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__21949\,
            I => \n2121_cascade_\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__21946\,
            I => \n2220_cascade_\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__21943\,
            I => \n2319_cascade_\
        );

    \I__1955\ : InMux
    port map (
            O => \N__21940\,
            I => \N__21937\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__21937\,
            I => n2097
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__21934\,
            I => \n2049_cascade_\
        );

    \I__1952\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21928\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__21928\,
            I => n2183
        );

    \I__1950\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21922\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__21922\,
            I => n2184
        );

    \I__1948\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21915\
        );

    \I__1947\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21912\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__21915\,
            I => \N__21909\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__21912\,
            I => \debounce.cnt_reg_3\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__21909\,
            I => \debounce.cnt_reg_3\
        );

    \I__1943\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21900\
        );

    \I__1942\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21897\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__21900\,
            I => \N__21894\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__21897\,
            I => \debounce.cnt_reg_9\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__21894\,
            I => \debounce.cnt_reg_9\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__1937\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21882\
        );

    \I__1936\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21879\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__21882\,
            I => \N__21876\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__21879\,
            I => \debounce.cnt_reg_5\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__21876\,
            I => \debounce.cnt_reg_5\
        );

    \I__1932\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21867\
        );

    \I__1931\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21864\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__21867\,
            I => \N__21861\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__21864\,
            I => \debounce.cnt_reg_8\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__21861\,
            I => \debounce.cnt_reg_8\
        );

    \I__1927\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21852\
        );

    \I__1926\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21849\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__21852\,
            I => \N__21846\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__21849\,
            I => \debounce.cnt_reg_1\
        );

    \I__1923\ : Odrv12
    port map (
            O => \N__21846\,
            I => \debounce.cnt_reg_1\
        );

    \I__1922\ : InMux
    port map (
            O => \N__21841\,
            I => \N__21837\
        );

    \I__1921\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21834\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__21837\,
            I => \N__21831\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__21834\,
            I => \debounce.cnt_reg_2\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__21831\,
            I => \debounce.cnt_reg_2\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__21826\,
            I => \debounce.n14472_cascade_\
        );

    \I__1916\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__21817\,
            I => n2095
        );

    \I__1913\ : InMux
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21808\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__21808\,
            I => \N__21805\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__21805\,
            I => n2094
        );

    \I__1909\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__21796\,
            I => n2101
        );

    \I__1906\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21790\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__21790\,
            I => n2200
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__21787\,
            I => \n2133_cascade_\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__21784\,
            I => \n2232_cascade_\
        );

    \I__1902\ : InMux
    port map (
            O => \N__21781\,
            I => n12122
        );

    \I__1901\ : InMux
    port map (
            O => \N__21778\,
            I => n12123
        );

    \I__1900\ : InMux
    port map (
            O => \N__21775\,
            I => n12124
        );

    \I__1899\ : InMux
    port map (
            O => \N__21772\,
            I => n12125
        );

    \I__1898\ : InMux
    port map (
            O => \N__21769\,
            I => n12126
        );

    \I__1897\ : InMux
    port map (
            O => \N__21766\,
            I => n12127
        );

    \I__1896\ : InMux
    port map (
            O => \N__21763\,
            I => n12128
        );

    \I__1895\ : InMux
    port map (
            O => \N__21760\,
            I => \bfn_1_32_0_\
        );

    \I__1894\ : InMux
    port map (
            O => \N__21757\,
            I => n12130
        );

    \I__1893\ : InMux
    port map (
            O => \N__21754\,
            I => \debounce.n12655\
        );

    \I__1892\ : InMux
    port map (
            O => \N__21751\,
            I => \debounce.n12656\
        );

    \I__1891\ : InMux
    port map (
            O => \N__21748\,
            I => \debounce.n12657\
        );

    \I__1890\ : InMux
    port map (
            O => \N__21745\,
            I => \debounce.n12658\
        );

    \I__1889\ : InMux
    port map (
            O => \N__21742\,
            I => \debounce.n12659\
        );

    \I__1888\ : InMux
    port map (
            O => \N__21739\,
            I => \debounce.n12660\
        );

    \I__1887\ : InMux
    port map (
            O => \N__21736\,
            I => \bfn_1_30_0_\
        );

    \I__1886\ : InMux
    port map (
            O => \N__21733\,
            I => \debounce.n12662\
        );

    \I__1885\ : InMux
    port map (
            O => \N__21730\,
            I => \bfn_1_31_0_\
        );

    \I__1884\ : InMux
    port map (
            O => \N__21727\,
            I => n12188
        );

    \I__1883\ : InMux
    port map (
            O => \N__21724\,
            I => n12189
        );

    \I__1882\ : InMux
    port map (
            O => \N__21721\,
            I => n12190
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__21718\,
            I => \n1427_cascade_\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__21715\,
            I => \n1430_cascade_\
        );

    \I__1879\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__21709\,
            I => n11638
        );

    \I__1877\ : InMux
    port map (
            O => \N__21706\,
            I => \bfn_1_29_0_\
        );

    \I__1876\ : InMux
    port map (
            O => \N__21703\,
            I => \debounce.n12654\
        );

    \I__1875\ : InMux
    port map (
            O => \N__21700\,
            I => n12179
        );

    \I__1874\ : InMux
    port map (
            O => \N__21697\,
            I => n12180
        );

    \I__1873\ : InMux
    port map (
            O => \N__21694\,
            I => n12181
        );

    \I__1872\ : InMux
    port map (
            O => \N__21691\,
            I => n12182
        );

    \I__1871\ : InMux
    port map (
            O => \N__21688\,
            I => n12183
        );

    \I__1870\ : InMux
    port map (
            O => \N__21685\,
            I => \bfn_1_27_0_\
        );

    \I__1869\ : InMux
    port map (
            O => \N__21682\,
            I => n12185
        );

    \I__1868\ : InMux
    port map (
            O => \N__21679\,
            I => n12186
        );

    \I__1867\ : InMux
    port map (
            O => \N__21676\,
            I => n12187
        );

    \I__1866\ : InMux
    port map (
            O => \N__21673\,
            I => n12216
        );

    \I__1865\ : InMux
    port map (
            O => \N__21670\,
            I => n12217
        );

    \I__1864\ : InMux
    port map (
            O => \N__21667\,
            I => n12218
        );

    \I__1863\ : InMux
    port map (
            O => \N__21664\,
            I => n12219
        );

    \I__1862\ : InMux
    port map (
            O => \N__21661\,
            I => n12220
        );

    \I__1861\ : InMux
    port map (
            O => \N__21658\,
            I => \bfn_1_25_0_\
        );

    \I__1860\ : InMux
    port map (
            O => \N__21655\,
            I => \bfn_1_26_0_\
        );

    \I__1859\ : InMux
    port map (
            O => \N__21652\,
            I => n12177
        );

    \I__1858\ : InMux
    port map (
            O => \N__21649\,
            I => n12178
        );

    \I__1857\ : InMux
    port map (
            O => \N__21646\,
            I => n12207
        );

    \I__1856\ : InMux
    port map (
            O => \N__21643\,
            I => n12208
        );

    \I__1855\ : InMux
    port map (
            O => \N__21640\,
            I => n12209
        );

    \I__1854\ : InMux
    port map (
            O => \N__21637\,
            I => n12210
        );

    \I__1853\ : InMux
    port map (
            O => \N__21634\,
            I => n12211
        );

    \I__1852\ : InMux
    port map (
            O => \N__21631\,
            I => n12212
        );

    \I__1851\ : InMux
    port map (
            O => \N__21628\,
            I => \bfn_1_24_0_\
        );

    \I__1850\ : InMux
    port map (
            O => \N__21625\,
            I => n12214
        );

    \I__1849\ : InMux
    port map (
            O => \N__21622\,
            I => n12215
        );

    \I__1848\ : InMux
    port map (
            O => \N__21619\,
            I => n12250
        );

    \I__1847\ : InMux
    port map (
            O => \N__21616\,
            I => n12251
        );

    \I__1846\ : InMux
    port map (
            O => \N__21613\,
            I => n12252
        );

    \I__1845\ : InMux
    port map (
            O => \N__21610\,
            I => n12253
        );

    \I__1844\ : InMux
    port map (
            O => \N__21607\,
            I => \bfn_1_22_0_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__21604\,
            I => n12255
        );

    \I__1842\ : InMux
    port map (
            O => \N__21601\,
            I => n12256
        );

    \I__1841\ : InMux
    port map (
            O => \N__21598\,
            I => \bfn_1_23_0_\
        );

    \I__1840\ : InMux
    port map (
            O => \N__21595\,
            I => n12206
        );

    \I__1839\ : InMux
    port map (
            O => \N__21592\,
            I => n12241
        );

    \I__1838\ : InMux
    port map (
            O => \N__21589\,
            I => n12242
        );

    \I__1837\ : InMux
    port map (
            O => \N__21586\,
            I => n12243
        );

    \I__1836\ : InMux
    port map (
            O => \N__21583\,
            I => n12244
        );

    \I__1835\ : InMux
    port map (
            O => \N__21580\,
            I => n12245
        );

    \I__1834\ : InMux
    port map (
            O => \N__21577\,
            I => \bfn_1_21_0_\
        );

    \I__1833\ : InMux
    port map (
            O => \N__21574\,
            I => n12247
        );

    \I__1832\ : InMux
    port map (
            O => \N__21571\,
            I => n12248
        );

    \I__1831\ : InMux
    port map (
            O => \N__21568\,
            I => n12249
        );

    \I__1830\ : InMux
    port map (
            O => \N__21565\,
            I => n12271
        );

    \I__1829\ : InMux
    port map (
            O => \N__21562\,
            I => \bfn_1_19_0_\
        );

    \I__1828\ : InMux
    port map (
            O => \N__21559\,
            I => n12273
        );

    \I__1827\ : InMux
    port map (
            O => \N__21556\,
            I => n12274
        );

    \I__1826\ : InMux
    port map (
            O => \N__21553\,
            I => n12275
        );

    \I__1825\ : InMux
    port map (
            O => \N__21550\,
            I => \bfn_1_20_0_\
        );

    \I__1824\ : InMux
    port map (
            O => \N__21547\,
            I => n12239
        );

    \I__1823\ : InMux
    port map (
            O => \N__21544\,
            I => n12240
        );

    \I__1822\ : InMux
    port map (
            O => \N__21541\,
            I => n12262
        );

    \I__1821\ : InMux
    port map (
            O => \N__21538\,
            I => n12263
        );

    \I__1820\ : InMux
    port map (
            O => \N__21535\,
            I => \bfn_1_18_0_\
        );

    \I__1819\ : InMux
    port map (
            O => \N__21532\,
            I => n12265
        );

    \I__1818\ : InMux
    port map (
            O => \N__21529\,
            I => n12266
        );

    \I__1817\ : InMux
    port map (
            O => \N__21526\,
            I => n12267
        );

    \I__1816\ : InMux
    port map (
            O => \N__21523\,
            I => n12268
        );

    \I__1815\ : InMux
    port map (
            O => \N__21520\,
            I => n12269
        );

    \I__1814\ : InMux
    port map (
            O => \N__21517\,
            I => n12270
        );

    \I__1813\ : InMux
    port map (
            O => \N__21514\,
            I => \bfn_1_17_0_\
        );

    \I__1812\ : InMux
    port map (
            O => \N__21511\,
            I => n12257
        );

    \I__1811\ : InMux
    port map (
            O => \N__21508\,
            I => n12258
        );

    \I__1810\ : InMux
    port map (
            O => \N__21505\,
            I => n12259
        );

    \I__1809\ : InMux
    port map (
            O => \N__21502\,
            I => n12260
        );

    \I__1808\ : InMux
    port map (
            O => \N__21499\,
            I => n12261
        );

    \I__1807\ : IoInMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__21493\,
            I => \N__21490\
        );

    \I__1805\ : IoSpan4Mux
    port map (
            O => \N__21490\,
            I => \N__21487\
        );

    \I__1804\ : IoSpan4Mux
    port map (
            O => \N__21487\,
            I => \N__21484\
        );

    \I__1803\ : IoSpan4Mux
    port map (
            O => \N__21484\,
            I => \N__21481\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__21481\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12528,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12536,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12544,
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_13_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_28_0_\
        );

    \IN_MUX_bfv_13_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12057,
            carryinitout => \bfn_13_29_0_\
        );

    \IN_MUX_bfv_13_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12065,
            carryinitout => \bfn_13_30_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12613,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12621,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_6_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_23_0_\
        );

    \IN_MUX_bfv_6_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n12630\,
            carryinitout => \bfn_6_24_0_\
        );

    \IN_MUX_bfv_6_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n12638\,
            carryinitout => \bfn_6_25_0_\
        );

    \IN_MUX_bfv_6_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n12646\,
            carryinitout => \bfn_6_26_0_\
        );

    \IN_MUX_bfv_16_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_26_0_\
        );

    \IN_MUX_bfv_16_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12670,
            carryinitout => \bfn_16_27_0_\
        );

    \IN_MUX_bfv_16_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12678,
            carryinitout => \bfn_16_28_0_\
        );

    \IN_MUX_bfv_14_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_26_0_\
        );

    \IN_MUX_bfv_14_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12080,
            carryinitout => \bfn_14_27_0_\
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12088,
            carryinitout => \bfn_14_28_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12582,
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_7_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12590,
            carryinitout => \bfn_7_27_0_\
        );

    \IN_MUX_bfv_7_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12598,
            carryinitout => \bfn_7_28_0_\
        );

    \IN_MUX_bfv_2_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_27_0_\
        );

    \IN_MUX_bfv_2_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12159,
            carryinitout => \bfn_2_28_0_\
        );

    \IN_MUX_bfv_3_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_29_0_\
        );

    \IN_MUX_bfv_3_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12148,
            carryinitout => \bfn_3_30_0_\
        );

    \IN_MUX_bfv_3_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_31_0_\
        );

    \IN_MUX_bfv_3_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12138,
            carryinitout => \bfn_3_32_0_\
        );

    \IN_MUX_bfv_1_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_31_0_\
        );

    \IN_MUX_bfv_1_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12129,
            carryinitout => \bfn_1_32_0_\
        );

    \IN_MUX_bfv_6_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_31_0_\
        );

    \IN_MUX_bfv_6_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12121,
            carryinitout => \bfn_6_32_0_\
        );

    \IN_MUX_bfv_7_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_30_0_\
        );

    \IN_MUX_bfv_7_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_29_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12499,
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12507,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12515,
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12471,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12479,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12487,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12444,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12452,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12460,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12418,
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12426,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12434,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12393,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12401,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12409,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12369,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12377,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12385,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12346,
            carryinitout => \bfn_6_15_0_\
        );

    \IN_MUX_bfv_6_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12354,
            carryinitout => \bfn_6_16_0_\
        );

    \IN_MUX_bfv_6_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_17_0_\
        );

    \IN_MUX_bfv_6_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12324,
            carryinitout => \bfn_6_18_0_\
        );

    \IN_MUX_bfv_6_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12332,
            carryinitout => \bfn_6_19_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12303,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12311,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12283,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12291,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_1_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_17_0_\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12264,
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12272,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12246,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12254,
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_2_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_21_0_\
        );

    \IN_MUX_bfv_2_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12229,
            carryinitout => \bfn_2_22_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12237,
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12213,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12221,
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_4_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_24_0_\
        );

    \IN_MUX_bfv_4_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12198,
            carryinitout => \bfn_4_25_0_\
        );

    \IN_MUX_bfv_1_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_26_0_\
        );

    \IN_MUX_bfv_1_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12184,
            carryinitout => \bfn_1_27_0_\
        );

    \IN_MUX_bfv_4_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_26_0_\
        );

    \IN_MUX_bfv_4_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12171,
            carryinitout => \bfn_4_27_0_\
        );

    \IN_MUX_bfv_12_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_27_0_\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_1_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \debounce.n12661\,
            carryinitout => \bfn_1_30_0_\
        );

    \IN_MUX_bfv_2_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_29_0_\
        );

    \IN_MUX_bfv_2_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12724,
            carryinitout => \bfn_2_30_0_\
        );

    \IN_MUX_bfv_2_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12732,
            carryinitout => \bfn_2_31_0_\
        );

    \IN_MUX_bfv_2_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12740,
            carryinitout => \bfn_2_32_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12559,
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12567,
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_5_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_28_0_\
        );

    \IN_MUX_bfv_11_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_29_0_\
        );

    \IN_MUX_bfv_11_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n12693\,
            carryinitout => \bfn_11_30_0_\
        );

    \IN_MUX_bfv_11_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n12701\,
            carryinitout => \bfn_11_31_0_\
        );

    \IN_MUX_bfv_11_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n12709\,
            carryinitout => \bfn_11_32_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21496\,
            GLOBALBUFFEROUTPUT => \CLK_N\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_2_lut_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27994\,
            in2 => \_gnd_net_\,
            in3 => \N__21514\,
            lcout => n2201,
            ltout => OPEN,
            carryin => \bfn_1_17_0_\,
            carryout => n12257,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_3_lut_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53827\,
            in2 => \N__26793\,
            in3 => \N__21511\,
            lcout => n2200,
            ltout => OPEN,
            carryin => n12257,
            carryout => n12258,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_4_lut_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26635\,
            in3 => \N__21508\,
            lcout => n2199,
            ltout => OPEN,
            carryin => n12258,
            carryout => n12259,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_5_lut_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53828\,
            in2 => \N__26710\,
            in3 => \N__21505\,
            lcout => n2198,
            ltout => OPEN,
            carryin => n12259,
            carryout => n12260,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_6_lut_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26743\,
            in3 => \N__21502\,
            lcout => n2197,
            ltout => OPEN,
            carryin => n12260,
            carryout => n12261,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_7_lut_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26773\,
            in3 => \N__21499\,
            lcout => n2196,
            ltout => OPEN,
            carryin => n12261,
            carryout => n12262,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_8_lut_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53830\,
            in2 => \N__24568\,
            in3 => \N__21541\,
            lcout => n2195,
            ltout => OPEN,
            carryin => n12262,
            carryout => n12263,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_9_lut_LC_1_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53829\,
            in2 => \N__29366\,
            in3 => \N__21538\,
            lcout => n2194,
            ltout => OPEN,
            carryin => n12263,
            carryout => n12264,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_10_lut_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53611\,
            in2 => \N__29177\,
            in3 => \N__21535\,
            lcout => n2193,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => n12265,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_11_lut_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29501\,
            in2 => \N__53990\,
            in3 => \N__21532\,
            lcout => n2192,
            ltout => OPEN,
            carryin => n12265,
            carryout => n12266,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_12_lut_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53615\,
            in2 => \N__29581\,
            in3 => \N__21529\,
            lcout => n2191,
            ltout => OPEN,
            carryin => n12266,
            carryout => n12267,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_13_lut_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53620\,
            in2 => \N__27112\,
            in3 => \N__21526\,
            lcout => n2190,
            ltout => OPEN,
            carryin => n12267,
            carryout => n12268,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_14_lut_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53616\,
            in2 => \N__24592\,
            in3 => \N__21523\,
            lcout => n2189,
            ltout => OPEN,
            carryin => n12268,
            carryout => n12269,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_15_lut_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53621\,
            in2 => \N__27087\,
            in3 => \N__21520\,
            lcout => n2188,
            ltout => OPEN,
            carryin => n12269,
            carryout => n12270,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_16_lut_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27607\,
            in2 => \N__53992\,
            in3 => \N__21517\,
            lcout => n2187,
            ltout => OPEN,
            carryin => n12270,
            carryout => n12271,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_17_lut_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27057\,
            in2 => \N__53991\,
            in3 => \N__21565\,
            lcout => n2186,
            ltout => OPEN,
            carryin => n12271,
            carryout => n12272,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_18_lut_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29692\,
            in2 => \N__54920\,
            in3 => \N__21562\,
            lcout => n2185,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => n12273,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_19_lut_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21991\,
            in2 => \N__54925\,
            in3 => \N__21559\,
            lcout => n2184,
            ltout => OPEN,
            carryin => n12273,
            carryout => n12274,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_20_lut_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22059\,
            in2 => \N__54921\,
            in3 => \N__21556\,
            lcout => n2183,
            ltout => OPEN,
            carryin => n12274,
            carryout => n12275,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_21_lut_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54517\,
            in1 => \N__36222\,
            in2 => \N__22048\,
            in3 => \N__21553\,
            lcout => n2214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12563_1_lut_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35994\,
            lcout => n15035,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_2_lut_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27922\,
            in2 => \_gnd_net_\,
            in3 => \N__21550\,
            lcout => n2101,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => n12239,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_3_lut_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54518\,
            in2 => \N__26671\,
            in3 => \N__21547\,
            lcout => n2100,
            ltout => OPEN,
            carryin => n12239,
            carryout => n12240,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_4_lut_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27181\,
            in3 => \N__21544\,
            lcout => n2099,
            ltout => OPEN,
            carryin => n12240,
            carryout => n12241,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_5_lut_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54519\,
            in2 => \N__24454\,
            in3 => \N__21592\,
            lcout => n2098,
            ltout => OPEN,
            carryin => n12241,
            carryout => n12242,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_6_lut_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24241\,
            in3 => \N__21589\,
            lcout => n2097,
            ltout => OPEN,
            carryin => n12242,
            carryout => n12243,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_7_lut_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24262\,
            in2 => \_gnd_net_\,
            in3 => \N__21586\,
            lcout => n2096,
            ltout => OPEN,
            carryin => n12243,
            carryout => n12244,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_8_lut_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54521\,
            in2 => \N__23034\,
            in3 => \N__21583\,
            lcout => n2095,
            ltout => OPEN,
            carryin => n12244,
            carryout => n12245,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_9_lut_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54520\,
            in2 => \N__24661\,
            in3 => \N__21580\,
            lcout => n2094,
            ltout => OPEN,
            carryin => n12245,
            carryout => n12246,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_10_lut_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54501\,
            in2 => \N__22981\,
            in3 => \N__21577\,
            lcout => n2093,
            ltout => OPEN,
            carryin => \bfn_1_21_0_\,
            carryout => n12247,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_11_lut_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29626\,
            in2 => \N__54922\,
            in3 => \N__21574\,
            lcout => n2092,
            ltout => OPEN,
            carryin => n12247,
            carryout => n12248,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_12_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54505\,
            in2 => \N__27139\,
            in3 => \N__21571\,
            lcout => n2091,
            ltout => OPEN,
            carryin => n12248,
            carryout => n12249,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_13_lut_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24628\,
            in2 => \N__54923\,
            in3 => \N__21568\,
            lcout => n2090,
            ltout => OPEN,
            carryin => n12249,
            carryout => n12250,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_14_lut_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54509\,
            in2 => \N__24165\,
            in3 => \N__21619\,
            lcout => n2089,
            ltout => OPEN,
            carryin => n12250,
            carryout => n12251,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_15_lut_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54531\,
            in2 => \N__27652\,
            in3 => \N__21616\,
            lcout => n2088,
            ltout => OPEN,
            carryin => n12251,
            carryout => n12252,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_16_lut_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54510\,
            in2 => \N__22894\,
            in3 => \N__21613\,
            lcout => n2087,
            ltout => OPEN,
            carryin => n12252,
            carryout => n12253,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_17_lut_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29712\,
            in2 => \N__54924\,
            in3 => \N__21610\,
            lcout => n2086,
            ltout => OPEN,
            carryin => n12253,
            carryout => n12254,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_18_lut_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22930\,
            in2 => \N__54934\,
            in3 => \N__21607\,
            lcout => n2085,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => n12255,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_19_lut_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22121\,
            in2 => \N__54935\,
            in3 => \N__21604\,
            lcout => n2084,
            ltout => OPEN,
            carryin => n12255,
            carryout => n12256,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_20_lut_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54535\,
            in1 => \N__22158\,
            in2 => \N__36072\,
            in3 => \N__21601\,
            lcout => n2115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_2_lut_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32694\,
            in2 => \_gnd_net_\,
            in3 => \N__21598\,
            lcout => n1901,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => n12206,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_3_lut_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54936\,
            in2 => \N__28024\,
            in3 => \N__21595\,
            lcout => n1900,
            ltout => OPEN,
            carryin => n12206,
            carryout => n12207,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_4_lut_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27711\,
            in3 => \N__21646\,
            lcout => n1899,
            ltout => OPEN,
            carryin => n12207,
            carryout => n12208,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_5_lut_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54937\,
            in2 => \N__27685\,
            in3 => \N__21643\,
            lcout => n1898,
            ltout => OPEN,
            carryin => n12208,
            carryout => n12209,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_6_lut_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27272\,
            in3 => \N__21640\,
            lcout => n1897,
            ltout => OPEN,
            carryin => n12209,
            carryout => n12210,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_7_lut_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27244\,
            in3 => \N__21637\,
            lcout => n1896,
            ltout => OPEN,
            carryin => n12210,
            carryout => n12211,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_8_lut_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54939\,
            in2 => \N__27742\,
            in3 => \N__21634\,
            lcout => n1895,
            ltout => OPEN,
            carryin => n12211,
            carryout => n12212,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_9_lut_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54938\,
            in2 => \N__27834\,
            in3 => \N__21631\,
            lcout => n1894,
            ltout => OPEN,
            carryin => n12212,
            carryout => n12213,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_10_lut_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54940\,
            in2 => \N__27808\,
            in3 => \N__21628\,
            lcout => n1893,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => n12214,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_11_lut_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54947\,
            in2 => \N__27858\,
            in3 => \N__21625\,
            lcout => n1892,
            ltout => OPEN,
            carryin => n12214,
            carryout => n12215,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_12_lut_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54941\,
            in2 => \N__27310\,
            in3 => \N__21622\,
            lcout => n1891,
            ltout => OPEN,
            carryin => n12215,
            carryout => n12216,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_13_lut_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27325\,
            in2 => \N__55134\,
            in3 => \N__21673\,
            lcout => n1890,
            ltout => OPEN,
            carryin => n12216,
            carryout => n12217,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_14_lut_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54945\,
            in2 => \N__27010\,
            in3 => \N__21670\,
            lcout => n1889,
            ltout => OPEN,
            carryin => n12217,
            carryout => n12218,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_15_lut_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54948\,
            in2 => \N__23161\,
            in3 => \N__21667\,
            lcout => n1888,
            ltout => OPEN,
            carryin => n12218,
            carryout => n12219,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_16_lut_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54946\,
            in2 => \N__23193\,
            in3 => \N__21664\,
            lcout => n1887,
            ltout => OPEN,
            carryin => n12219,
            carryout => n12220,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_17_lut_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54949\,
            in2 => \N__24385\,
            in3 => \N__21661\,
            lcout => n1886,
            ltout => OPEN,
            carryin => n12220,
            carryout => n12221,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_18_lut_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__54950\,
            in1 => \_gnd_net_\,
            in2 => \N__27414\,
            in3 => \N__21658\,
            lcout => n1885,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_2_lut_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28098\,
            in2 => \_gnd_net_\,
            in3 => \N__21655\,
            lcout => n1701,
            ltout => OPEN,
            carryin => \bfn_1_26_0_\,
            carryout => n12177,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_3_lut_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54581\,
            in2 => \N__23448\,
            in3 => \N__21652\,
            lcout => n1700,
            ltout => OPEN,
            carryin => n12177,
            carryout => n12178,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_4_lut_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23473\,
            in3 => \N__21649\,
            lcout => n1699,
            ltout => OPEN,
            carryin => n12178,
            carryout => n12179,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_5_lut_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54582\,
            in2 => \N__22339\,
            in3 => \N__21700\,
            lcout => n1698,
            ltout => OPEN,
            carryin => n12179,
            carryout => n12180,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_6_lut_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22263\,
            in3 => \N__21697\,
            lcout => n1697,
            ltout => OPEN,
            carryin => n12180,
            carryout => n12181,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_7_lut_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22360\,
            in3 => \N__21694\,
            lcout => n1696,
            ltout => OPEN,
            carryin => n12181,
            carryout => n12182,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_8_lut_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54951\,
            in2 => \N__23289\,
            in3 => \N__21691\,
            lcout => n1695,
            ltout => OPEN,
            carryin => n12182,
            carryout => n12183,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_9_lut_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54583\,
            in2 => \N__23668\,
            in3 => \N__21688\,
            lcout => n1694,
            ltout => OPEN,
            carryin => n12183,
            carryout => n12184,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_10_lut_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55135\,
            in2 => \N__23506\,
            in3 => \N__21685\,
            lcout => n1693,
            ltout => OPEN,
            carryin => \bfn_1_27_0_\,
            carryout => n12185,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_11_lut_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55140\,
            in2 => \N__23419\,
            in3 => \N__21682\,
            lcout => n1692,
            ltout => OPEN,
            carryin => n12185,
            carryout => n12186,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_12_lut_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55136\,
            in2 => \N__23260\,
            in3 => \N__21679\,
            lcout => n1691,
            ltout => OPEN,
            carryin => n12186,
            carryout => n12187,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_13_lut_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55141\,
            in2 => \N__23395\,
            in3 => \N__21676\,
            lcout => n1690,
            ltout => OPEN,
            carryin => n12187,
            carryout => n12188,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_14_lut_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23604\,
            in2 => \N__55219\,
            in3 => \N__21727\,
            lcout => n1689,
            ltout => OPEN,
            carryin => n12188,
            carryout => n12189,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_15_lut_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23532\,
            in2 => \N__55218\,
            in3 => \N__21724\,
            lcout => n1688,
            ltout => OPEN,
            carryin => n12189,
            carryout => n12190,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_16_lut_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__55145\,
            in1 => \N__35520\,
            in2 => \N__25642\,
            in3 => \N__21721\,
            lcout => n1719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i907_3_lut_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23797\,
            in2 => \N__28336\,
            in3 => \N__36743\,
            lcout => n1427,
            ltout => \n1427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_73_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21718\,
            in3 => \N__25515\,
            lcout => n14088,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i910_3_lut_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23818\,
            in2 => \N__26194\,
            in3 => \N__36744\,
            lcout => n1430,
            ltout => \n1430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_74_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__25938\,
            in1 => \N__26061\,
            in2 => \N__21715\,
            in3 => \N__21712\,
            lcout => n13334,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9924_3_lut_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23578\,
            in2 => \N__23707\,
            in3 => \N__23741\,
            lcout => n11638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.cnt_reg_636__i0_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22650\,
            in2 => \_gnd_net_\,
            in3 => \N__21706\,
            lcout => \debounce.cnt_reg_0\,
            ltout => OPEN,
            carryin => \bfn_1_29_0_\,
            carryout => \debounce.n12654\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i1_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21855\,
            in2 => \_gnd_net_\,
            in3 => \N__21703\,
            lcout => \debounce.cnt_reg_1\,
            ltout => OPEN,
            carryin => \debounce.n12654\,
            carryout => \debounce.n12655\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i2_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21840\,
            in2 => \_gnd_net_\,
            in3 => \N__21754\,
            lcout => \debounce.cnt_reg_2\,
            ltout => OPEN,
            carryin => \debounce.n12655\,
            carryout => \debounce.n12656\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i3_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21918\,
            in2 => \_gnd_net_\,
            in3 => \N__21751\,
            lcout => \debounce.cnt_reg_3\,
            ltout => OPEN,
            carryin => \debounce.n12656\,
            carryout => \debounce.n12657\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i4_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22686\,
            in2 => \_gnd_net_\,
            in3 => \N__21748\,
            lcout => \debounce.cnt_reg_4\,
            ltout => OPEN,
            carryin => \debounce.n12657\,
            carryout => \debounce.n12658\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i5_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21885\,
            in2 => \_gnd_net_\,
            in3 => \N__21745\,
            lcout => \debounce.cnt_reg_5\,
            ltout => OPEN,
            carryin => \debounce.n12658\,
            carryout => \debounce.n12659\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i6_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22671\,
            in2 => \_gnd_net_\,
            in3 => \N__21742\,
            lcout => \debounce.cnt_reg_6\,
            ltout => OPEN,
            carryin => \debounce.n12659\,
            carryout => \debounce.n12660\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i7_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22635\,
            in2 => \_gnd_net_\,
            in3 => \N__21739\,
            lcout => \debounce.cnt_reg_7\,
            ltout => OPEN,
            carryin => \debounce.n12660\,
            carryout => \debounce.n12661\,
            clk => \N__56042\,
            ce => 'H',
            sr => \N__23887\
        );

    \debounce.cnt_reg_636__i8_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21870\,
            in2 => \_gnd_net_\,
            in3 => \N__21736\,
            lcout => \debounce.cnt_reg_8\,
            ltout => OPEN,
            carryin => \bfn_1_30_0_\,
            carryout => \debounce.n12662\,
            clk => \N__56044\,
            ce => 'H',
            sr => \N__23886\
        );

    \debounce.cnt_reg_636__i9_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21903\,
            in2 => \_gnd_net_\,
            in3 => \N__21733\,
            lcout => \debounce.cnt_reg_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56044\,
            ce => 'H',
            sr => \N__23886\
        );

    \encoder0_position_31__I_0_add_766_2_lut_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28176\,
            in2 => \_gnd_net_\,
            in3 => \N__21730\,
            lcout => n1201,
            ltout => OPEN,
            carryin => \bfn_1_31_0_\,
            carryout => n12122,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_3_lut_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55220\,
            in2 => \N__28633\,
            in3 => \N__21781\,
            lcout => n1200,
            ltout => OPEN,
            carryin => n12122,
            carryout => n12123,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_4_lut_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28687\,
            in3 => \N__21778\,
            lcout => n1199,
            ltout => OPEN,
            carryin => n12123,
            carryout => n12124,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_5_lut_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55221\,
            in2 => \N__30457\,
            in3 => \N__21775\,
            lcout => n1198,
            ltout => OPEN,
            carryin => n12124,
            carryout => n12125,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_6_lut_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26395\,
            in3 => \N__21772\,
            lcout => n1197,
            ltout => OPEN,
            carryin => n12125,
            carryout => n12126,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_7_lut_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28663\,
            in3 => \N__21769\,
            lcout => n1196,
            ltout => OPEN,
            carryin => n12126,
            carryout => n12127,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_8_lut_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55223\,
            in2 => \N__30550\,
            in3 => \N__21766\,
            lcout => n1195,
            ltout => OPEN,
            carryin => n12127,
            carryout => n12128,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_9_lut_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55222\,
            in2 => \N__28765\,
            in3 => \N__21763\,
            lcout => n1194,
            ltout => OPEN,
            carryin => n12128,
            carryout => n12129,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_10_lut_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55224\,
            in2 => \N__28788\,
            in3 => \N__21760\,
            lcout => n1193,
            ltout => OPEN,
            carryin => \bfn_1_32_0_\,
            carryout => n12130,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_11_lut_LC_1_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__55225\,
            in1 => \N__36570\,
            in2 => \N__28807\,
            in3 => \N__21757\,
            lcout => n1224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i12061_4_lut_LC_1_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21919\,
            in1 => \N__21904\,
            in2 => \N__21889\,
            in3 => \N__21871\,
            lcout => OPEN,
            ltout => \debounce.n14472_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i2_4_lut_LC_1_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__21856\,
            in1 => \N__21841\,
            in2 => \N__21826\,
            in3 => \N__22621\,
            lcout => n13490,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1383_3_lut_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21823\,
            in2 => \N__23035\,
            in3 => \N__35987\,
            lcout => n2127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1382_3_lut_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21814\,
            in2 => \N__36017\,
            in3 => \N__24660\,
            lcout => n2126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37554\,
            lcout => n23_adj_647,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1389_3_lut_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21802\,
            in1 => \N__27921\,
            in2 => \_gnd_net_\,
            in3 => \N__35986\,
            lcout => n2133,
            ltout => \n2133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1456_3_lut_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__21793\,
            in1 => \_gnd_net_\,
            in2 => \N__21787\,
            in3 => \N__36168\,
            lcout => n2232,
            ltout => \n2232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1523_3_lut_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31456\,
            in1 => \_gnd_net_\,
            in2 => \N__21784\,
            in3 => \N__39145\,
            lcout => n2331,
            ltout => \n2331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1590_3_lut_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22606\,
            in2 => \N__21970\,
            in3 => \N__34929\,
            lcout => n2430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12587_1_lut_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36158\,
            lcout => n15059,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1377_3_lut_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24166\,
            in2 => \N__21967\,
            in3 => \N__35993\,
            lcout => n2121,
            ltout => \n2121_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1444_3_lut_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21955\,
            in2 => \N__21949\,
            in3 => \N__36157\,
            lcout => n2220,
            ltout => \n2220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1511_3_lut_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31642\,
            in2 => \N__21946\,
            in3 => \N__39134\,
            lcout => n2319,
            ltout => \n2319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1578_3_lut_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22750\,
            in2 => \N__21943\,
            in3 => \N__34935\,
            lcout => n2418,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12566_4_lut_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22125\,
            in1 => \N__22929\,
            in2 => \N__22165\,
            in3 => \N__22774\,
            lcout => n2049,
            ltout => \n2049_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1385_3_lut_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21940\,
            in1 => \_gnd_net_\,
            in2 => \N__21934\,
            in3 => \N__24240\,
            lcout => n2129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1439_3_lut_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21931\,
            in2 => \N__22063\,
            in3 => \N__36159\,
            lcout => n2215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1440_3_lut_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__21990\,
            in1 => \N__21925\,
            in2 => \N__36193\,
            in3 => \_gnd_net_\,
            lcout => n2216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1372_3_lut_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22072\,
            in2 => \N__22132\,
            in3 => \N__35985\,
            lcout => n2116,
            ltout => \n2116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12590_4_lut_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21989\,
            in1 => \N__22044\,
            in2 => \N__22030\,
            in3 => \N__27022\,
            lcout => n2148,
            ltout => \n2148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1451_3_lut_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24561\,
            in2 => \N__22027\,
            in3 => \N__22024\,
            lcout => n2227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1375_3_lut_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22015\,
            in1 => \_gnd_net_\,
            in2 => \N__36015\,
            in3 => \N__22889\,
            lcout => n2119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1381_3_lut_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22009\,
            in2 => \N__22980\,
            in3 => \N__35978\,
            lcout => n2125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1373_3_lut_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__22922\,
            in1 => \_gnd_net_\,
            in2 => \N__36016\,
            in3 => \N__22003\,
            lcout => n2117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_2_lut_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37603\,
            in2 => \_gnd_net_\,
            in3 => \N__21976\,
            lcout => n2001,
            ltout => OPEN,
            carryin => \bfn_2_21_0_\,
            carryout => n12222,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_3_lut_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53790\,
            in2 => \N__27493\,
            in3 => \N__21973\,
            lcout => n2000,
            ltout => OPEN,
            carryin => n12222,
            carryout => n12223,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_4_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26935\,
            in3 => \N__22102\,
            lcout => n1999,
            ltout => OPEN,
            carryin => n12223,
            carryout => n12224,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_5_lut_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53791\,
            in2 => \N__26908\,
            in3 => \N__22099\,
            lcout => n1998,
            ltout => OPEN,
            carryin => n12224,
            carryout => n12225,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_6_lut_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27454\,
            in3 => \N__22096\,
            lcout => n1997,
            ltout => OPEN,
            carryin => n12225,
            carryout => n12226,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_7_lut_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27538\,
            in3 => \N__22093\,
            lcout => n1996,
            ltout => OPEN,
            carryin => n12226,
            carryout => n12227,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_8_lut_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54254\,
            in2 => \N__24693\,
            in3 => \N__22090\,
            lcout => n1995,
            ltout => OPEN,
            carryin => n12227,
            carryout => n12228,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_9_lut_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53792\,
            in2 => \N__24805\,
            in3 => \N__22087\,
            lcout => n1994,
            ltout => OPEN,
            carryin => n12228,
            carryout => n12229,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_10_lut_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54255\,
            in2 => \N__24499\,
            in3 => \N__22084\,
            lcout => n1993,
            ltout => OPEN,
            carryin => \bfn_2_22_0_\,
            carryout => n12230,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_11_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54926\,
            in2 => \N__24408\,
            in3 => \N__22081\,
            lcout => n1992,
            ltout => OPEN,
            carryin => n12230,
            carryout => n12231,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_12_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54256\,
            in2 => \N__23112\,
            in3 => \N__22078\,
            lcout => n1991,
            ltout => OPEN,
            carryin => n12231,
            carryout => n12232,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_13_lut_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54927\,
            in2 => \N__24183\,
            in3 => \N__22075\,
            lcout => n1990,
            ltout => OPEN,
            carryin => n12232,
            carryout => n12233,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_14_lut_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24765\,
            in2 => \N__55132\,
            in3 => \N__22183\,
            lcout => n1989,
            ltout => OPEN,
            carryin => n12233,
            carryout => n12234,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_15_lut_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26973\,
            in2 => \N__54729\,
            in3 => \N__22180\,
            lcout => n1988,
            ltout => OPEN,
            carryin => n12234,
            carryout => n12235,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_16_lut_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24725\,
            in2 => \N__55133\,
            in3 => \N__22177\,
            lcout => n1987,
            ltout => OPEN,
            carryin => n12235,
            carryout => n12236,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_17_lut_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24513\,
            in2 => \N__54730\,
            in3 => \N__22174\,
            lcout => n1986,
            ltout => OPEN,
            carryin => n12236,
            carryout => n12237,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_18_lut_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24530\,
            in2 => \N__54731\,
            in3 => \N__22171\,
            lcout => n1985,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => n12238,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_19_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54266\,
            in1 => \N__35910\,
            in2 => \N__27379\,
            in3 => \N__22168\,
            lcout => n2016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1240_3_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22144\,
            in2 => \N__23160\,
            in3 => \N__35765\,
            lcout => n1920,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1182_3_lut_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24978\,
            in2 => \N__24964\,
            in3 => \N__35594\,
            lcout => n1830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1305_3_lut_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__35895\,
            in1 => \N__22138\,
            in2 => \N__24537\,
            in3 => \_gnd_net_\,
            lcout => n2017,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1116_3_lut_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__35481\,
            in1 => \N__23449\,
            in2 => \N__22240\,
            in3 => \_gnd_net_\,
            lcout => n1732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1115_3_lut_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23472\,
            in1 => \N__35482\,
            in2 => \_gnd_net_\,
            in3 => \N__22228\,
            lcout => n1731,
            ltout => \n1731_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9979_4_lut_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__28048\,
            in1 => \N__25044\,
            in2 => \N__22219\,
            in3 => \N__25004\,
            lcout => n11694,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1113_3_lut_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35483\,
            in2 => \N__22267\,
            in3 => \N__22216\,
            lcout => n1729,
            ltout => \n1729_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_81_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24927\,
            in2 => \N__22207\,
            in3 => \_gnd_net_\,
            lcout => n14116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1117_3_lut_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22204\,
            in1 => \N__28099\,
            in2 => \_gnd_net_\,
            in3 => \N__35480\,
            lcout => n1733,
            ltout => \n1733_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1184_3_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25033\,
            in2 => \N__22195\,
            in3 => \N__35584\,
            lcout => n1832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1238_3_lut_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24377\,
            in2 => \N__22192\,
            in3 => \N__35766\,
            lcout => n1918,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_148_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__22334\,
            in1 => \N__22256\,
            in2 => \N__22359\,
            in3 => \N__23425\,
            lcout => n13343,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1114_3_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22312\,
            in2 => \N__35492\,
            in3 => \N__22335\,
            lcout => n1730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1112_3_lut_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__22355\,
            in1 => \_gnd_net_\,
            in2 => \N__22306\,
            in3 => \N__35476\,
            lcout => n1728,
            ltout => \n1728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_79_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24848\,
            in2 => \N__22297\,
            in3 => \N__27872\,
            lcout => n13962,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12374_3_lut_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22294\,
            in2 => \N__23290\,
            in3 => \N__35469\,
            lcout => n1727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12477_1_lut_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35491\,
            in3 => \_gnd_net_\,
            lcout => n14949,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1110_3_lut_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23663\,
            in2 => \N__22288\,
            in3 => \N__35468\,
            lcout => n1726,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1105_3_lut_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23611\,
            in2 => \N__35493\,
            in3 => \N__22279\,
            lcout => n1721,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1046_3_lut_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__25402\,
            in1 => \N__25416\,
            in2 => \N__35388\,
            in3 => \_gnd_net_\,
            lcout => n1630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1049_3_lut_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25060\,
            in2 => \N__27574\,
            in3 => \N__35364\,
            lcout => n1633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_127_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__25352\,
            in1 => \N__23356\,
            in2 => \N__25389\,
            in3 => \N__23752\,
            lcout => OPEN,
            ltout => \n13986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12825_4_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25725\,
            in1 => \N__25689\,
            in2 => \N__22366\,
            in3 => \N__25662\,
            lcout => n1554,
            ltout => \n1554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1042_3_lut_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25296\,
            in1 => \_gnd_net_\,
            in2 => \N__22363\,
            in3 => \N__25270\,
            lcout => n1626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1044_rep_37_3_lut_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25353\,
            in2 => \N__25339\,
            in3 => \N__35365\,
            lcout => n1628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1045_3_lut_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25385\,
            in1 => \_gnd_net_\,
            in2 => \N__35389\,
            in3 => \N__25369\,
            lcout => n1629,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1047_3_lut_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25462\,
            in2 => \N__25432\,
            in3 => \N__35372\,
            lcout => n1631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_2_lut_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23577\,
            in2 => \_gnd_net_\,
            in3 => \N__22321\,
            lcout => n1501,
            ltout => OPEN,
            carryin => \bfn_2_27_0_\,
            carryout => n12152,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_3_lut_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54732\,
            in2 => \N__23706\,
            in3 => \N__22318\,
            lcout => n1500,
            ltout => OPEN,
            carryin => n12152,
            carryout => n12153,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_4_lut_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23742\,
            in3 => \N__22315\,
            lcout => n1499,
            ltout => OPEN,
            carryin => n12153,
            carryout => n12154,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_5_lut_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54733\,
            in2 => \N__25942\,
            in3 => \N__22396\,
            lcout => n1498,
            ltout => OPEN,
            carryin => n12154,
            carryout => n12155,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_6_lut_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23634\,
            in2 => \_gnd_net_\,
            in3 => \N__22393\,
            lcout => n1497,
            ltout => OPEN,
            carryin => n12155,
            carryout => n12156,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_7_lut_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26065\,
            in3 => \N__22390\,
            lcout => n1496,
            ltout => OPEN,
            carryin => n12156,
            carryout => n12157,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_8_lut_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54734\,
            in2 => \N__25522\,
            in3 => \N__22387\,
            lcout => n1495,
            ltout => OPEN,
            carryin => n12157,
            carryout => n12158,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_9_lut_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25614\,
            in2 => \N__55061\,
            in3 => \N__22384\,
            lcout => n1494,
            ltout => OPEN,
            carryin => n12158,
            carryout => n12159,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_10_lut_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54744\,
            in2 => \N__25972\,
            in3 => \N__22381\,
            lcout => n1493,
            ltout => OPEN,
            carryin => \bfn_2_28_0_\,
            carryout => n12160,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_11_lut_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25846\,
            in2 => \N__55062\,
            in3 => \N__22378\,
            lcout => n1492,
            ltout => OPEN,
            carryin => n12160,
            carryout => n12161,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_12_lut_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54748\,
            in2 => \N__26134\,
            in3 => \N__22375\,
            lcout => n1491,
            ltout => OPEN,
            carryin => n12161,
            carryout => n12162,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_13_lut_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54742\,
            in2 => \N__25900\,
            in3 => \N__22372\,
            lcout => n1490,
            ltout => OPEN,
            carryin => n12162,
            carryout => n12163,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_14_lut_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54743\,
            in1 => \N__25882\,
            in2 => \N__35310\,
            in3 => \N__22369\,
            lcout => n1521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12804_1_lut_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35275\,
            lcout => n15276,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i971_3_lut_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26133\,
            in2 => \N__35286\,
            in3 => \N__22456\,
            lcout => n1523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i0_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22450\,
            in2 => \_gnd_net_\,
            in3 => \N__22444\,
            lcout => n26_adj_678,
            ltout => OPEN,
            carryin => \bfn_2_29_0_\,
            carryout => n12717,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i1_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22441\,
            in2 => \_gnd_net_\,
            in3 => \N__22435\,
            lcout => n25_adj_677,
            ltout => OPEN,
            carryin => n12717,
            carryout => n12718,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i2_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22432\,
            in2 => \_gnd_net_\,
            in3 => \N__22426\,
            lcout => n24_adj_676,
            ltout => OPEN,
            carryin => n12718,
            carryout => n12719,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i3_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22423\,
            in2 => \_gnd_net_\,
            in3 => \N__22417\,
            lcout => n23_adj_675,
            ltout => OPEN,
            carryin => n12719,
            carryout => n12720,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i4_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22414\,
            in2 => \_gnd_net_\,
            in3 => \N__22408\,
            lcout => n22_adj_674,
            ltout => OPEN,
            carryin => n12720,
            carryout => n12721,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i5_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22405\,
            in2 => \_gnd_net_\,
            in3 => \N__22399\,
            lcout => n21_adj_673,
            ltout => OPEN,
            carryin => n12721,
            carryout => n12722,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i6_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22537\,
            in2 => \_gnd_net_\,
            in3 => \N__22531\,
            lcout => n20_adj_672,
            ltout => OPEN,
            carryin => n12722,
            carryout => n12723,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i7_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22528\,
            in2 => \_gnd_net_\,
            in3 => \N__22522\,
            lcout => n19_adj_671,
            ltout => OPEN,
            carryin => n12723,
            carryout => n12724,
            clk => \N__56045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i8_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22519\,
            in2 => \_gnd_net_\,
            in3 => \N__22513\,
            lcout => n18_adj_670,
            ltout => OPEN,
            carryin => \bfn_2_30_0_\,
            carryout => n12725,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i9_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22510\,
            in2 => \_gnd_net_\,
            in3 => \N__22504\,
            lcout => n17_adj_669,
            ltout => OPEN,
            carryin => n12725,
            carryout => n12726,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i10_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22501\,
            in2 => \_gnd_net_\,
            in3 => \N__22495\,
            lcout => n16_adj_668,
            ltout => OPEN,
            carryin => n12726,
            carryout => n12727,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i11_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22492\,
            in2 => \_gnd_net_\,
            in3 => \N__22486\,
            lcout => n15_adj_667,
            ltout => OPEN,
            carryin => n12727,
            carryout => n12728,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i12_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22483\,
            in2 => \_gnd_net_\,
            in3 => \N__22477\,
            lcout => n14_adj_666,
            ltout => OPEN,
            carryin => n12728,
            carryout => n12729,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i13_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22474\,
            in2 => \_gnd_net_\,
            in3 => \N__22468\,
            lcout => n13_adj_665,
            ltout => OPEN,
            carryin => n12729,
            carryout => n12730,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i14_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22465\,
            in2 => \_gnd_net_\,
            in3 => \N__22459\,
            lcout => n12_adj_664,
            ltout => OPEN,
            carryin => n12730,
            carryout => n12731,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i15_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22597\,
            in2 => \_gnd_net_\,
            in3 => \N__22591\,
            lcout => n11_adj_663,
            ltout => OPEN,
            carryin => n12731,
            carryout => n12732,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i16_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22588\,
            in2 => \_gnd_net_\,
            in3 => \N__22582\,
            lcout => n10_adj_662,
            ltout => OPEN,
            carryin => \bfn_2_31_0_\,
            carryout => n12733,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i17_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22579\,
            in2 => \_gnd_net_\,
            in3 => \N__22573\,
            lcout => n9_adj_661,
            ltout => OPEN,
            carryin => n12733,
            carryout => n12734,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i18_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22570\,
            in2 => \_gnd_net_\,
            in3 => \N__22564\,
            lcout => n8_adj_660,
            ltout => OPEN,
            carryin => n12734,
            carryout => n12735,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i19_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22561\,
            in2 => \_gnd_net_\,
            in3 => \N__22555\,
            lcout => n7_adj_659,
            ltout => OPEN,
            carryin => n12735,
            carryout => n12736,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i20_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22552\,
            in2 => \_gnd_net_\,
            in3 => \N__22546\,
            lcout => n6_adj_658,
            ltout => OPEN,
            carryin => n12736,
            carryout => n12737,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i21_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36825\,
            in2 => \_gnd_net_\,
            in3 => \N__22543\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n12737,
            carryout => n12738,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i22_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36804\,
            in2 => \_gnd_net_\,
            in3 => \N__22540\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n12738,
            carryout => n12739,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i23_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36783\,
            in2 => \_gnd_net_\,
            in3 => \N__22696\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n12739,
            carryout => n12740,
            clk => \N__56051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i24_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36843\,
            in2 => \_gnd_net_\,
            in3 => \N__22693\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_2_32_0_\,
            carryout => n12741,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_634__i25_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36882\,
            in2 => \_gnd_net_\,
            in3 => \N__22690\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i5_4_lut_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__22687\,
            in1 => \N__22672\,
            in2 => \N__22657\,
            in3 => \N__22636\,
            lcout => \debounce.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i2_LC_2_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23907\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \reg_B_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_2_lut_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37516\,
            in2 => \_gnd_net_\,
            in3 => \N__22615\,
            lcout => n2401,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => n12296,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_3_lut_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53415\,
            in2 => \N__26533\,
            in3 => \N__22612\,
            lcout => n2400,
            ltout => OPEN,
            carryin => n12296,
            carryout => n12297,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_4_lut_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26872\,
            in3 => \N__22609\,
            lcout => n2399,
            ltout => OPEN,
            carryin => n12297,
            carryout => n12298,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_5_lut_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53416\,
            in2 => \N__26841\,
            in3 => \N__22600\,
            lcout => n2398,
            ltout => OPEN,
            carryin => n12298,
            carryout => n12299,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_6_lut_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24316\,
            in3 => \N__22723\,
            lcout => n2397,
            ltout => OPEN,
            carryin => n12299,
            carryout => n12300,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_7_lut_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24054\,
            in3 => \N__22720\,
            lcout => n2396,
            ltout => OPEN,
            carryin => n12300,
            carryout => n12301,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_8_lut_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53418\,
            in2 => \N__32394\,
            in3 => \N__22717\,
            lcout => n2395,
            ltout => OPEN,
            carryin => n12301,
            carryout => n12302,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_9_lut_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53417\,
            in2 => \N__32362\,
            in3 => \N__22714\,
            lcout => n2394,
            ltout => OPEN,
            carryin => n12302,
            carryout => n12303,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_10_lut_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53764\,
            in2 => \N__32302\,
            in3 => \N__22711\,
            lcout => n2393,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => n12304,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_11_lut_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53767\,
            in2 => \N__32278\,
            in3 => \N__22708\,
            lcout => n2392,
            ltout => OPEN,
            carryin => n12304,
            carryout => n12305,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_12_lut_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53765\,
            in2 => \N__32425\,
            in3 => \N__22705\,
            lcout => n2391,
            ltout => OPEN,
            carryin => n12305,
            carryout => n12306,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_13_lut_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53768\,
            in2 => \N__32245\,
            in3 => \N__22702\,
            lcout => n2390,
            ltout => OPEN,
            carryin => n12306,
            carryout => n12307,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_14_lut_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53766\,
            in2 => \N__32335\,
            in3 => \N__22699\,
            lcout => n2389,
            ltout => OPEN,
            carryin => n12307,
            carryout => n12308,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_15_lut_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53769\,
            in2 => \N__32455\,
            in3 => \N__22756\,
            lcout => n2388,
            ltout => OPEN,
            carryin => n12308,
            carryout => n12309,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_16_lut_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32655\,
            in2 => \N__54248\,
            in3 => \N__22753\,
            lcout => n2387,
            ltout => OPEN,
            carryin => n12309,
            carryout => n12310,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_17_lut_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53773\,
            in2 => \N__32640\,
            in3 => \N__22744\,
            lcout => n2386,
            ltout => OPEN,
            carryin => n12310,
            carryout => n12311,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_18_lut_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24333\,
            in2 => \N__54249\,
            in3 => \N__22741\,
            lcout => n2385,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => n12312,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_19_lut_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24108\,
            in2 => \N__54252\,
            in3 => \N__22738\,
            lcout => n2384,
            ltout => OPEN,
            carryin => n12312,
            carryout => n12313,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_20_lut_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39012\,
            in2 => \N__54250\,
            in3 => \N__22735\,
            lcout => n2383,
            ltout => OPEN,
            carryin => n12313,
            carryout => n12314,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_21_lut_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29539\,
            in2 => \N__54253\,
            in3 => \N__22732\,
            lcout => n2382,
            ltout => OPEN,
            carryin => n12314,
            carryout => n12315,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_22_lut_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26596\,
            in2 => \N__54251\,
            in3 => \N__22729\,
            lcout => n2381,
            ltout => OPEN,
            carryin => n12315,
            carryout => n12316,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_23_lut_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53789\,
            in1 => \N__34950\,
            in2 => \N__31921\,
            in3 => \N__22726\,
            lcout => n2412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1386_3_lut_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22852\,
            in2 => \N__24453\,
            in3 => \N__35991\,
            lcout => n2130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1584_3_lut_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32276\,
            in2 => \N__22840\,
            in3 => \N__34906\,
            lcout => n2424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1384_3_lut_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22831\,
            in2 => \N__24261\,
            in3 => \N__35992\,
            lcout => n2128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1453_3_lut_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26732\,
            in2 => \N__22822\,
            in3 => \N__36150\,
            lcout => n2229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1316_3_lut_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27537\,
            in1 => \_gnd_net_\,
            in2 => \N__35894\,
            in3 => \N__22807\,
            lcout => n2028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1452_3_lut_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26762\,
            in2 => \N__22801\,
            in3 => \N__36149\,
            lcout => n2228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1457_3_lut_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27993\,
            in2 => \N__36191\,
            in3 => \N__22786\,
            lcout => n2233,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_95_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29705\,
            in1 => \N__27635\,
            in2 => \N__22890\,
            in3 => \N__24208\,
            lcout => n14160,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1442_3_lut_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22768\,
            in2 => \N__36192\,
            in3 => \N__27053\,
            lcout => n2218,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_92_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24644\,
            in1 => \N__29615\,
            in2 => \N__22976\,
            in3 => \N__23021\,
            lcout => n14146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1309_3_lut_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24766\,
            in2 => \N__23005\,
            in3 => \N__35863\,
            lcout => n2021,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1318_3_lut_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22996\,
            in1 => \_gnd_net_\,
            in2 => \N__35888\,
            in3 => \N__26904\,
            lcout => n2030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1314_3_lut_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__24798\,
            in1 => \_gnd_net_\,
            in2 => \N__22990\,
            in3 => \N__35858\,
            lcout => n2026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1239_3_lut_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35747\,
            in1 => \N__22951\,
            in2 => \_gnd_net_\,
            in3 => \N__23194\,
            lcout => n1919,
            ltout => \n1919_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1306_3_lut_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22939\,
            in2 => \N__22933\,
            in3 => \N__35867\,
            lcout => n2018,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1308_3_lut_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26974\,
            in1 => \_gnd_net_\,
            in2 => \N__35889\,
            in3 => \N__22900\,
            lcout => n2020,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1307_3_lut_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24733\,
            in2 => \N__22867\,
            in3 => \N__35862\,
            lcout => n2019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1311_3_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22858\,
            in2 => \N__23113\,
            in3 => \N__35875\,
            lcout => n2023,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1244_3_lut_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__35727\,
            in1 => \N__27859\,
            in2 => \N__23128\,
            in3 => \_gnd_net_\,
            lcout => n1924,
            ltout => \n1924_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_87_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24794\,
            in2 => \N__23095\,
            in3 => \N__24401\,
            lcout => n13770,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1245_3_lut_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27801\,
            in2 => \N__35752\,
            in3 => \N__23092\,
            lcout => n1925,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1243_3_lut_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__27306\,
            in1 => \_gnd_net_\,
            in2 => \N__23080\,
            in3 => \N__35726\,
            lcout => n1923,
            ltout => \n1923_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_88_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24494\,
            in2 => \N__23065\,
            in3 => \N__24686\,
            lcout => n13772,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1248_3_lut_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__35725\,
            in1 => \_gnd_net_\,
            in2 => \N__23062\,
            in3 => \N__27236\,
            lcout => n1928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1251_3_lut_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23047\,
            in2 => \N__27712\,
            in3 => \N__35721\,
            lcout => n1931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1174_3_lut_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__25189\,
            in1 => \N__25211\,
            in2 => \N__35622\,
            in3 => \_gnd_net_\,
            lcout => n1822,
            ltout => \n1822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_86_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23150\,
            in2 => \N__23038\,
            in3 => \N__23180\,
            lcout => n14134,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1246_3_lut_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23218\,
            in2 => \N__27835\,
            in3 => \N__35720\,
            lcout => n1926,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12540_1_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35890\,
            in3 => \_gnd_net_\,
            lcout => n15012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1104_3_lut_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35487\,
            in1 => \_gnd_net_\,
            in2 => \N__23539\,
            in3 => \N__23209\,
            lcout => n1720,
            ltout => \n1720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1171_3_lut_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35600\,
            in2 => \N__23197\,
            in3 => \N__25096\,
            lcout => n1819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12497_1_lut_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35595\,
            lcout => n14969,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1172_3_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25134\,
            in1 => \_gnd_net_\,
            in2 => \N__35621\,
            in3 => \N__25120\,
            lcout => n1820,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12500_4_lut_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25107\,
            in1 => \N__25133\,
            in2 => \N__23311\,
            in3 => \N__25080\,
            lcout => n1752,
            ltout => \n1752_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1176_3_lut_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25245\,
            in1 => \_gnd_net_\,
            in2 => \N__23164\,
            in3 => \N__25225\,
            lcout => n1824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1173_3_lut_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35599\,
            in2 => \N__25153\,
            in3 => \N__25173\,
            lcout => n1821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_149_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23266\,
            in1 => \N__23388\,
            in2 => \N__23253\,
            in3 => \N__23134\,
            lcout => OPEN,
            ltout => \n14110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12480_4_lut_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25638\,
            in1 => \N__23603\,
            in2 => \N__23350\,
            in3 => \N__23531\,
            lcout => n1653,
            ltout => \n1653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1107_3_lut_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23249\,
            in1 => \_gnd_net_\,
            in2 => \N__23347\,
            in3 => \N__23344\,
            lcout => n1723,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_80_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25241\,
            in1 => \N__27341\,
            in2 => \N__25212\,
            in3 => \N__23332\,
            lcout => OPEN,
            ltout => \n13968_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_82_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__25169\,
            in1 => \N__23326\,
            in2 => \N__23320\,
            in3 => \N__23317\,
            lcout => n13972,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1106_3_lut_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23387\,
            in1 => \N__35486\,
            in2 => \_gnd_net_\,
            in3 => \N__23302\,
            lcout => n1722,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_147_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23501\,
            in1 => \N__23282\,
            in2 => \N__23664\,
            in3 => \N__23408\,
            lcout => n14104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1040_3_lut_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__25555\,
            in1 => \_gnd_net_\,
            in2 => \N__25759\,
            in3 => \N__35382\,
            lcout => n1624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1108_3_lut_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__35484\,
            in1 => \_gnd_net_\,
            in2 => \N__23233\,
            in3 => \N__23409\,
            lcout => n1724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1109_3_lut_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23502\,
            in2 => \N__23488\,
            in3 => \N__35485\,
            lcout => n1725,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29897\,
            lcout => n13_adj_637,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1048_3_lut_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__25488\,
            in1 => \_gnd_net_\,
            in2 => \N__25474\,
            in3 => \N__35373\,
            lcout => n1632,
            ltout => \n1632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9920_3_lut_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__28097\,
            in1 => \_gnd_net_\,
            in2 => \N__23452\,
            in3 => \N__23441\,
            lcout => n11634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1041_3_lut_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25255\,
            in2 => \N__25591\,
            in3 => \N__35378\,
            lcout => n1625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1039_3_lut_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25810\,
            in2 => \N__35391\,
            in3 => \N__25741\,
            lcout => n1623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12820_1_lut_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35374\,
            lcout => n15292,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i979_3_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23743\,
            in2 => \N__23368\,
            in3 => \N__35282\,
            lcout => n1531,
            ltout => \n1531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9983_4_lut_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__25487\,
            in1 => \N__27570\,
            in2 => \N__23359\,
            in3 => \N__25454\,
            lcout => n11698,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1043_3_lut_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__25306\,
            in1 => \N__25323\,
            in2 => \N__35390\,
            in3 => \_gnd_net_\,
            lcout => n1627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i977_3_lut_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__23641\,
            in1 => \N__23623\,
            in2 => \N__35279\,
            in3 => \_gnd_net_\,
            lcout => n1529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29928\,
            lcout => n14_adj_638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i978_3_lut_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23617\,
            in2 => \N__35280\,
            in3 => \N__25934\,
            lcout => n1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1038_3_lut_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25724\,
            in2 => \N__25702\,
            in3 => \N__35384\,
            lcout => n1622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i20_3_lut_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29929\,
            in1 => \N__33271\,
            in2 => \_gnd_net_\,
            in3 => \N__39546\,
            lcout => n300,
            ltout => \n300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i981_3_lut_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23560\,
            in2 => \N__23554\,
            in3 => \N__35258\,
            lcout => n1533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i970_3_lut_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25896\,
            in2 => \N__35281\,
            in3 => \N__23551\,
            lcout => n1522,
            ltout => \n1522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1037_3_lut_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25678\,
            in2 => \N__23542\,
            in3 => \N__35383\,
            lcout => n1621,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i975_3_lut_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25514\,
            in2 => \N__23773\,
            in3 => \N__35246\,
            lcout => n1527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i976_3_lut_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__26054\,
            in1 => \N__23764\,
            in2 => \N__35274\,
            in3 => \_gnd_net_\,
            lcout => n1528,
            ltout => \n1528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_78_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23758\,
            in3 => \N__25286\,
            lcout => OPEN,
            ltout => \n13978_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_126_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25544\,
            in1 => \N__25802\,
            in2 => \N__23755\,
            in3 => \N__25583\,
            lcout => n13984,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i912_3_lut_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__25776\,
            in1 => \_gnd_net_\,
            in2 => \N__23833\,
            in3 => \N__36720\,
            lcout => n1432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_75_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26121\,
            in1 => \N__25964\,
            in2 => \N__25845\,
            in3 => \N__23716\,
            lcout => n14094,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i913_3_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23677\,
            in1 => \N__26110\,
            in2 => \_gnd_net_\,
            in3 => \N__36721\,
            lcout => n1433,
            ltout => \n1433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i980_3_lut_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35247\,
            in1 => \_gnd_net_\,
            in2 => \N__23686\,
            in3 => \N__23683\,
            lcout => n1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_2_lut_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26109\,
            in2 => \_gnd_net_\,
            in3 => \N__23671\,
            lcout => n1401,
            ltout => OPEN,
            carryin => \bfn_3_29_0_\,
            carryout => n12141,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_3_lut_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54738\,
            in2 => \N__25777\,
            in3 => \N__23824\,
            lcout => n1400,
            ltout => OPEN,
            carryin => n12141,
            carryout => n12142,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_4_lut_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26307\,
            in3 => \N__23821\,
            lcout => n1399,
            ltout => OPEN,
            carryin => n12142,
            carryout => n12143,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_5_lut_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54739\,
            in2 => \N__26187\,
            in3 => \N__23806\,
            lcout => n1398,
            ltout => OPEN,
            carryin => n12143,
            carryout => n12144,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_6_lut_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26092\,
            in3 => \N__23803\,
            lcout => n1397,
            ltout => OPEN,
            carryin => n12144,
            carryout => n12145,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_7_lut_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26019\,
            in2 => \_gnd_net_\,
            in3 => \N__23800\,
            lcout => n1396,
            ltout => OPEN,
            carryin => n12145,
            carryout => n12146,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_8_lut_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54741\,
            in2 => \N__28329\,
            in3 => \N__23785\,
            lcout => n1395,
            ltout => OPEN,
            carryin => n12146,
            carryout => n12147,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_9_lut_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54740\,
            in2 => \N__28362\,
            in3 => \N__23782\,
            lcout => n1394,
            ltout => OPEN,
            carryin => n12147,
            carryout => n12148,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_10_lut_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55070\,
            in2 => \N__28389\,
            in3 => \N__23779\,
            lcout => n1393,
            ltout => OPEN,
            carryin => \bfn_3_30_0_\,
            carryout => n12149,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_11_lut_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55072\,
            in2 => \N__28408\,
            in3 => \N__23776\,
            lcout => n1392,
            ltout => OPEN,
            carryin => n12149,
            carryout => n12150,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_12_lut_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26216\,
            in2 => \N__55209\,
            in3 => \N__23866\,
            lcout => n1391,
            ltout => OPEN,
            carryin => n12150,
            carryout => n12151,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_13_lut_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__55071\,
            in1 => \N__36756\,
            in2 => \N__26164\,
            in3 => \N__23863\,
            lcout => n1422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i842_3_lut_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23842\,
            in2 => \N__28516\,
            in3 => \N__36629\,
            lcout => n1330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i2_4_lut_adj_26_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__28143\,
            in1 => \N__28119\,
            in2 => \N__28450\,
            in3 => \N__28473\,
            lcout => \debounce.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i843_3_lut_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28263\,
            in2 => \N__23854\,
            in3 => \N__36628\,
            lcout => n1331,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_2_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28300\,
            in2 => \_gnd_net_\,
            in3 => \N__23860\,
            lcout => n1301,
            ltout => OPEN,
            carryin => \bfn_3_31_0_\,
            carryout => n12131,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_3_lut_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55063\,
            in2 => \N__28282\,
            in3 => \N__23857\,
            lcout => n1300,
            ltout => OPEN,
            carryin => n12131,
            carryout => n12132,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_4_lut_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28264\,
            in3 => \N__23845\,
            lcout => n1299,
            ltout => OPEN,
            carryin => n12132,
            carryout => n12133,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_5_lut_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55064\,
            in2 => \N__28515\,
            in3 => \N__23836\,
            lcout => n1298,
            ltout => OPEN,
            carryin => n12133,
            carryout => n12134,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_6_lut_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28558\,
            in3 => \N__23947\,
            lcout => n1297,
            ltout => OPEN,
            carryin => n12134,
            carryout => n12135,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_7_lut_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28537\,
            in3 => \N__23944\,
            lcout => n1296,
            ltout => OPEN,
            carryin => n12135,
            carryout => n12136,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_8_lut_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55066\,
            in2 => \N__28231\,
            in3 => \N__23941\,
            lcout => n1295,
            ltout => OPEN,
            carryin => n12136,
            carryout => n12137,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_9_lut_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55065\,
            in2 => \N__28594\,
            in3 => \N__23938\,
            lcout => n1294,
            ltout => OPEN,
            carryin => n12137,
            carryout => n12138,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_10_lut_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55067\,
            in2 => \N__28714\,
            in3 => \N__23935\,
            lcout => n1293,
            ltout => OPEN,
            carryin => \bfn_3_32_0_\,
            carryout => n12139,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_11_lut_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55068\,
            in2 => \N__26256\,
            in3 => \N__23932\,
            lcout => n1292,
            ltout => OPEN,
            carryin => n12139,
            carryout => n12140,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_12_lut_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__55069\,
            in1 => \N__36663\,
            in2 => \N__26353\,
            in3 => \N__23929\,
            lcout => n1323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i2_LC_3_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__27944\,
            in1 => \N__23926\,
            in2 => \_gnd_net_\,
            in3 => \N__38070\,
            lcout => h1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56057\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i3_4_lut_LC_3_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011111111"
        )
    port map (
            in0 => \N__23925\,
            in1 => \N__23917\,
            in2 => \N__23908\,
            in3 => \N__27943\,
            lcout => \debounce.cnt_next_9__N_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i769_3_lut_LC_3_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36541\,
            in2 => \N__28789\,
            in3 => \N__24010\,
            lcout => n1225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_104_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31395\,
            in3 => \N__31358\,
            lcout => n14410,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1454_3_lut_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24001\,
            in2 => \N__36207\,
            in3 => \N__26709\,
            lcout => n2230,
            ltout => \n2230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1521_3_lut_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__39133\,
            in1 => \_gnd_net_\,
            in2 => \N__23992\,
            in3 => \N__31378\,
            lcout => n2329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1656_3_lut_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28960\,
            in2 => \N__28980\,
            in3 => \N__35046\,
            lcout => n2528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1445_3_lut_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24588\,
            in2 => \N__23989\,
            in3 => \N__36194\,
            lcout => n2221,
            ltout => \n2221_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1512_3_lut_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31678\,
            in2 => \N__23974\,
            in3 => \N__39132\,
            lcout => n2320,
            ltout => \n2320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1579_3_lut_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34925\,
            in1 => \_gnd_net_\,
            in2 => \N__23971\,
            in3 => \N__23968\,
            lcout => n2419,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1591_3_lut_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26871\,
            in2 => \N__23962\,
            in3 => \N__34924\,
            lcout => n2431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1589_3_lut_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23953\,
            in2 => \N__34927\,
            in3 => \N__24312\,
            lcout => n2429,
            ltout => \n2429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_114_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__29411\,
            in1 => \N__29018\,
            in2 => \N__24076\,
            in3 => \N__26461\,
            lcout => n13423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_112_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28937\,
            in1 => \N__30884\,
            in2 => \N__31239\,
            in3 => \N__31292\,
            lcout => OPEN,
            ltout => \n14210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_113_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30681\,
            in1 => \N__28895\,
            in2 => \N__24073\,
            in3 => \N__29207\,
            lcout => OPEN,
            ltout => \n14214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_115_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31138\,
            in1 => \N__31019\,
            in2 => \N__24070\,
            in3 => \N__24067\,
            lcout => n14220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1588_3_lut_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24061\,
            in2 => \N__24055\,
            in3 => \N__34896\,
            lcout => n2428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_110_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__24308\,
            in1 => \N__24053\,
            in2 => \N__26821\,
            in3 => \N__32605\,
            lcout => OPEN,
            ltout => \n14016_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_111_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24329\,
            in1 => \N__24104\,
            in2 => \N__24028\,
            in3 => \N__39011\,
            lcout => OPEN,
            ltout => \n14022_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12879_4_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26592\,
            in1 => \N__29538\,
            in2 => \N__24025\,
            in3 => \N__31917\,
            lcout => n2346,
            ltout => \n2346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1587_3_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24022\,
            in2 => \N__24013\,
            in3 => \N__32384\,
            lcout => n2427,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1576_3_lut_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34905\,
            in1 => \N__24127\,
            in2 => \N__24109\,
            in3 => \_gnd_net_\,
            lcout => n2416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1577_3_lut_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24121\,
            in1 => \_gnd_net_\,
            in2 => \N__24334\,
            in3 => \N__34904\,
            lcout => n2417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1581_3_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24115\,
            in2 => \N__34928\,
            in3 => \N__32334\,
            lcout => n2421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12876_1_lut_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34900\,
            lcout => n15348,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1509_3_lut_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32088\,
            in2 => \N__32074\,
            in3 => \N__39072\,
            lcout => n2317,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10059_4_lut_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__31517\,
            in1 => \N__32160\,
            in2 => \N__31437\,
            in3 => \N__31476\,
            lcout => OPEN,
            ltout => \n11774_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_105_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__31659\,
            in1 => \N__24091\,
            in2 => \N__24082\,
            in3 => \N__29464\,
            lcout => OPEN,
            ltout => \n14188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_106_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__32121\,
            in2 => \N__24079\,
            in3 => \N__39179\,
            lcout => n14194,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1520_3_lut_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31333\,
            in1 => \_gnd_net_\,
            in2 => \N__31362\,
            in3 => \N__39067\,
            lcout => n2328,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1443_3_lut_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24349\,
            in2 => \N__36206\,
            in3 => \N__27606\,
            lcout => n2219,
            ltout => \n2219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1510_3_lut_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32110\,
            in1 => \_gnd_net_\,
            in2 => \N__24337\,
            in3 => \N__39071\,
            lcout => n2318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1522_3_lut_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__31433\,
            in1 => \_gnd_net_\,
            in2 => \N__39105\,
            in3 => \N__31414\,
            lcout => n2330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1387_3_lut_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24289\,
            in1 => \_gnd_net_\,
            in2 => \N__27180\,
            in3 => \N__36031\,
            lcout => n2131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1317_3_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35870\,
            in2 => \N__24277\,
            in3 => \N__27453\,
            lcout => n2029,
            ltout => \n2029_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_94_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__24224\,
            in1 => \N__24424\,
            in2 => \N__24211\,
            in3 => \N__24133\,
            lcout => n14154,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1310_3_lut_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35869\,
            in2 => \N__24202\,
            in3 => \N__24187\,
            lcout => n2022,
            ltout => \n2022_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_93_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27128\,
            in1 => \N__24620\,
            in2 => \N__24142\,
            in3 => \N__24139\,
            lcout => n14152,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1315_3_lut_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35868\,
            in2 => \N__24694\,
            in3 => \N__24670\,
            lcout => n2027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1378_3_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__24624\,
            in1 => \_gnd_net_\,
            in2 => \N__24604\,
            in3 => \N__36032\,
            lcout => n2122,
            ltout => \n2122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_97_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__24557\,
            in1 => \_gnd_net_\,
            in2 => \N__24541\,
            in3 => \N__29505\,
            lcout => n13748,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12543_4_lut_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24538\,
            in1 => \N__27372\,
            in2 => \N__24514\,
            in3 => \N__24703\,
            lcout => n1950,
            ltout => \n1950_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1313_3_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24498\,
            in1 => \_gnd_net_\,
            in2 => \N__24478\,
            in3 => \N__24475\,
            lcout => n2025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1319_3_lut_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24466\,
            in2 => \N__26931\,
            in3 => \N__35874\,
            lcout => n2031,
            ltout => \n2031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9965_4_lut_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__27164\,
            in1 => \N__26661\,
            in2 => \N__24427\,
            in3 => \N__27914\,
            lcout => n11680,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1312_3_lut_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24418\,
            in2 => \N__24409\,
            in3 => \N__35873\,
            lcout => n2024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12521_4_lut_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24378\,
            in1 => \N__24355\,
            in2 => \N__27211\,
            in3 => \N__27413\,
            lcout => n1851,
            ltout => \n1851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1247_3_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27741\,
            in1 => \_gnd_net_\,
            in2 => \N__24820\,
            in3 => \N__24817\,
            lcout => n1927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1181_3_lut_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24916\,
            in2 => \N__24946\,
            in3 => \N__35620\,
            lcout => n1829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1242_3_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27324\,
            in1 => \_gnd_net_\,
            in2 => \N__35761\,
            in3 => \N__24778\,
            lcout => n1922,
            ltout => \n1922_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_89_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26960\,
            in1 => \N__24748\,
            in2 => \N__24742\,
            in3 => \N__24739\,
            lcout => OPEN,
            ltout => \n13778_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_91_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__27508\,
            in1 => \N__24729\,
            in2 => \N__24706\,
            in3 => \N__26878\,
            lcout => n13782,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1183_3_lut_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__35619\,
            in1 => \N__24991\,
            in2 => \N__25021\,
            in3 => \_gnd_net_\,
            lcout => n1831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1179_3_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24874\,
            in2 => \N__24904\,
            in3 => \N__35615\,
            lcout => n1827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12375_3_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24832\,
            in2 => \N__35628\,
            in3 => \N__24864\,
            lcout => n1826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_2_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28043\,
            in2 => \_gnd_net_\,
            in3 => \N__24697\,
            lcout => n1801,
            ltout => OPEN,
            carryin => \bfn_4_24_0_\,
            carryout => n12191,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_3_lut_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25048\,
            in2 => \N__54589\,
            in3 => \N__25024\,
            lcout => n1800,
            ltout => OPEN,
            carryin => n12191,
            carryout => n12192,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_4_lut_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25017\,
            in3 => \N__24985\,
            lcout => n1799,
            ltout => OPEN,
            carryin => n12192,
            carryout => n12193,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_5_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54083\,
            in2 => \N__24982\,
            in3 => \N__24949\,
            lcout => n1798,
            ltout => OPEN,
            carryin => n12193,
            carryout => n12194,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_6_lut_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24945\,
            in3 => \N__24910\,
            lcout => n1797,
            ltout => OPEN,
            carryin => n12194,
            carryout => n12195,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_7_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27771\,
            in3 => \N__24907\,
            lcout => n1796,
            ltout => OPEN,
            carryin => n12195,
            carryout => n12196,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_8_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54082\,
            in2 => \N__24903\,
            in3 => \N__24868\,
            lcout => n1795,
            ltout => OPEN,
            carryin => n12196,
            carryout => n12197,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_9_lut_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54084\,
            in2 => \N__24865\,
            in3 => \N__24826\,
            lcout => n1794,
            ltout => OPEN,
            carryin => n12197,
            carryout => n12198,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_10_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55162\,
            in2 => \N__27885\,
            in3 => \N__24823\,
            lcout => n1793,
            ltout => OPEN,
            carryin => \bfn_4_25_0_\,
            carryout => n12199,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_11_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55166\,
            in2 => \N__25246\,
            in3 => \N__25219\,
            lcout => n1792,
            ltout => OPEN,
            carryin => n12199,
            carryout => n12200,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_12_lut_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55163\,
            in2 => \N__27348\,
            in3 => \N__25216\,
            lcout => n1791,
            ltout => OPEN,
            carryin => n12200,
            carryout => n12201,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_13_lut_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55167\,
            in2 => \N__25213\,
            in3 => \N__25177\,
            lcout => n1790,
            ltout => OPEN,
            carryin => n12201,
            carryout => n12202,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_14_lut_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55164\,
            in2 => \N__25174\,
            in3 => \N__25144\,
            lcout => n1789,
            ltout => OPEN,
            carryin => n12202,
            carryout => n12203,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_15_lut_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55168\,
            in2 => \N__25141\,
            in3 => \N__25114\,
            lcout => n1788,
            ltout => OPEN,
            carryin => n12203,
            carryout => n12204,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_16_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25111\,
            in2 => \N__55226\,
            in3 => \N__25087\,
            lcout => n1787,
            ltout => OPEN,
            carryin => n12204,
            carryout => n12205,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_17_lut_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__55165\,
            in1 => \N__25084\,
            in2 => \N__35646\,
            in3 => \N__25063\,
            lcout => n1818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_2_lut_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27563\,
            in2 => \_gnd_net_\,
            in3 => \N__25051\,
            lcout => n1601,
            ltout => OPEN,
            carryin => \bfn_4_26_0_\,
            carryout => n12164,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_3_lut_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54057\,
            in2 => \N__25492\,
            in3 => \N__25465\,
            lcout => n1600,
            ltout => OPEN,
            carryin => n12164,
            carryout => n12165,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_4_lut_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25461\,
            in3 => \N__25420\,
            lcout => n1599,
            ltout => OPEN,
            carryin => n12165,
            carryout => n12166,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_5_lut_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54058\,
            in2 => \N__25417\,
            in3 => \N__25393\,
            lcout => n1598,
            ltout => OPEN,
            carryin => n12166,
            carryout => n12167,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_6_lut_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25390\,
            in3 => \N__25360\,
            lcout => n1597,
            ltout => OPEN,
            carryin => n12167,
            carryout => n12168,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_7_lut_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25357\,
            in3 => \N__25327\,
            lcout => n1596,
            ltout => OPEN,
            carryin => n12168,
            carryout => n12169,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_8_lut_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54580\,
            in2 => \N__25324\,
            in3 => \N__25300\,
            lcout => n1595,
            ltout => OPEN,
            carryin => n12169,
            carryout => n12170,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_9_lut_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54059\,
            in2 => \N__25297\,
            in3 => \N__25258\,
            lcout => n1594,
            ltout => OPEN,
            carryin => n12170,
            carryout => n12171,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_10_lut_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54771\,
            in2 => \N__25590\,
            in3 => \N__25249\,
            lcout => n1593,
            ltout => OPEN,
            carryin => \bfn_4_27_0_\,
            carryout => n12172,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_11_lut_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54584\,
            in2 => \N__25551\,
            in3 => \N__25744\,
            lcout => n1592,
            ltout => OPEN,
            carryin => n12172,
            carryout => n12173,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_12_lut_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54772\,
            in2 => \N__25809\,
            in3 => \N__25735\,
            lcout => n1591,
            ltout => OPEN,
            carryin => n12173,
            carryout => n12174,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_13_lut_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54585\,
            in2 => \N__25732\,
            in3 => \N__25693\,
            lcout => n1590,
            ltout => OPEN,
            carryin => n12174,
            carryout => n12175,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_14_lut_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25690\,
            in2 => \N__54975\,
            in3 => \N__25672\,
            lcout => n1589,
            ltout => OPEN,
            carryin => n12175,
            carryout => n12176,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_15_lut_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54773\,
            in1 => \N__35409\,
            in2 => \N__25669\,
            in3 => \N__25645\,
            lcout => n1620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i974_3_lut_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25621\,
            in2 => \N__25603\,
            in3 => \N__35257\,
            lcout => n1526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i973_3_lut_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25968\,
            in2 => \N__25567\,
            in3 => \N__35256\,
            lcout => n1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i908_3_lut_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25528\,
            in2 => \N__26026\,
            in3 => \N__36711\,
            lcout => n1428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i905_3_lut_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25990\,
            in2 => \N__36733\,
            in3 => \N__28390\,
            lcout => n1425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i906_3_lut_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36715\,
            in2 => \N__28366\,
            in3 => \N__25981\,
            lcout => n1426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i911_3_lut_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__26308\,
            in1 => \N__25948\,
            in2 => \N__36732\,
            in3 => \_gnd_net_\,
            lcout => n1431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i903_3_lut_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26221\,
            in2 => \N__25912\,
            in3 => \N__36719\,
            lcout => n1423,
            ltout => \n1423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12807_4_lut_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25881\,
            in1 => \N__25864\,
            in2 => \N__25855\,
            in3 => \N__25852\,
            lcout => n1455,
            ltout => \n1455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i972_3_lut_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25844\,
            in2 => \N__25822\,
            in3 => \N__25819\,
            lcout => n1524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i845_3_lut_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25786\,
            in1 => \N__28296\,
            in2 => \_gnd_net_\,
            in3 => \N__36627\,
            lcout => n1333,
            ltout => \n1333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9926_3_lut_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26108\,
            in2 => \N__25762\,
            in3 => \N__26300\,
            lcout => OPEN,
            ltout => \n11640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_72_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__26090\,
            in1 => \N__26018\,
            in2 => \N__26197\,
            in3 => \N__26183\,
            lcout => OPEN,
            ltout => \n13315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12790_4_lut_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26220\,
            in1 => \N__26160\,
            in2 => \N__26146\,
            in3 => \N__28306\,
            lcout => n1356,
            ltout => \n1356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i904_3_lut_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28404\,
            in2 => \N__26143\,
            in3 => \N__26140\,
            lcout => n1424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i21_3_lut_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39535\,
            in1 => \N__33244\,
            in2 => \_gnd_net_\,
            in3 => \N__29905\,
            lcout => n299,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12787_1_lut_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36739\,
            in3 => \_gnd_net_\,
            lcout => n15259,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i909_3_lut_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26091\,
            in2 => \N__26074\,
            in3 => \N__36725\,
            lcout => n1429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i841_3_lut_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26032\,
            in2 => \N__28557\,
            in3 => \N__36626\,
            lcout => n1329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i839_3_lut_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28227\,
            in2 => \N__36635\,
            in3 => \N__26002\,
            lcout => n1327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i838_3_lut_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25996\,
            in2 => \N__28593\,
            in3 => \N__36618\,
            lcout => n1326,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12774_4_lut_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28483\,
            in1 => \N__26352\,
            in2 => \N__26260\,
            in3 => \N__28693\,
            lcout => n1257,
            ltout => \n1257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12771_1_lut_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26332\,
            in3 => \_gnd_net_\,
            lcout => n15243,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i777_3_lut_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28169\,
            in1 => \N__26329\,
            in2 => \_gnd_net_\,
            in3 => \N__36537\,
            lcout => n1233,
            ltout => \n1233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i844_3_lut_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26317\,
            in2 => \N__26311\,
            in3 => \N__36625\,
            lcout => n1332,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i840_3_lut_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26284\,
            in1 => \_gnd_net_\,
            in2 => \N__36636\,
            in3 => \N__28536\,
            lcout => n1328,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i770_3_lut_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28758\,
            in2 => \N__36546\,
            in3 => \N__26278\,
            lcout => n1226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i776_3_lut_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26269\,
            in2 => \N__28629\,
            in3 => \N__36529\,
            lcout => n1232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i836_3_lut_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26252\,
            in2 => \N__26230\,
            in3 => \N__36630\,
            lcout => n1324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12755_4_lut_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__28800\,
            in1 => \N__26359\,
            in2 => \N__26368\,
            in3 => \N__28738\,
            lcout => n1158,
            ltout => \n1158_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12752_1_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26416\,
            in3 => \_gnd_net_\,
            lcout => n15224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i775_3_lut_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28683\,
            in2 => \N__36545\,
            in3 => \N__26413\,
            lcout => n1231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i773_3_lut_LC_4_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26404\,
            in2 => \N__26391\,
            in3 => \N__36536\,
            lcout => n1229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i706_3_lut_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30343\,
            in2 => \N__33904\,
            in3 => \N__36957\,
            lcout => n1130,
            ltout => \n1130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_68_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26371\,
            in3 => \N__28649\,
            lcout => n14068,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9991_4_lut_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__28177\,
            in1 => \N__28682\,
            in2 => \N__30453\,
            in3 => \N__28622\,
            lcout => n11706,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i1_LC_4_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38171\,
            in1 => \N__28120\,
            in2 => \_gnd_net_\,
            in3 => \N__27945\,
            lcout => h2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_118_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37391\,
            in1 => \N__30728\,
            in2 => \N__34511\,
            in3 => \N__30800\,
            lcout => n13798,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1709_3_lut_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30972\,
            in2 => \N__38943\,
            in3 => \N__28849\,
            lcout => n2613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1653_3_lut_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29134\,
            in2 => \N__31240\,
            in3 => \N__35048\,
            lcout => n2525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1655_3_lut_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28921\,
            in1 => \_gnd_net_\,
            in2 => \N__35092\,
            in3 => \N__28941\,
            lcout => n2527,
            ltout => \n2527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_119_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34346\,
            in1 => \N__30665\,
            in2 => \N__26443\,
            in3 => \N__30852\,
            lcout => OPEN,
            ltout => \n13796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_120_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26440\,
            in1 => \N__34598\,
            in2 => \N__26434\,
            in3 => \N__31107\,
            lcout => n13804,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1654_3_lut_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28876\,
            in1 => \_gnd_net_\,
            in2 => \N__28912\,
            in3 => \N__35047\,
            lcout => n2526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_116_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29105\,
            in2 => \N__29073\,
            in3 => \N__29322\,
            lcout => OPEN,
            ltout => \n14354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_117_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31571\,
            in1 => \N__29279\,
            in2 => \N__26431\,
            in3 => \N__26428\,
            lcout => OPEN,
            ltout => \n14224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12906_4_lut_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31193\,
            in1 => \N__29782\,
            in2 => \N__26422\,
            in3 => \N__29248\,
            lcout => n2445,
            ltout => \n2445_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1649_3_lut_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29106\,
            in1 => \_gnd_net_\,
            in2 => \N__26419\,
            in3 => \N__29092\,
            lcout => n2521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1650_3_lut_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29119\,
            in2 => \N__31297\,
            in3 => \N__35085\,
            lcout => n2522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1645_3_lut_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29323\,
            in1 => \_gnd_net_\,
            in2 => \N__35108\,
            in3 => \N__29299\,
            lcout => n2517,
            ltout => \n2517_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_122_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29734\,
            in1 => \N__31049\,
            in2 => \N__26509\,
            in3 => \N__26506\,
            lcout => n13810,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1646_3_lut_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29069\,
            in2 => \N__35107\,
            in3 => \N__29053\,
            lcout => n2518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1642_3_lut_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29263\,
            in2 => \N__29284\,
            in3 => \N__35053\,
            lcout => n2514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29691\,
            in1 => \_gnd_net_\,
            in2 => \N__26500\,
            in3 => \N__36205\,
            lcout => n2217,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1582_3_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__26488\,
            in1 => \_gnd_net_\,
            in2 => \N__34926\,
            in3 => \N__32241\,
            lcout => n2422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1593_3_lut_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37505\,
            in1 => \N__26476\,
            in2 => \_gnd_net_\,
            in3 => \N__34890\,
            lcout => n2433,
            ltout => \n2433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9955_3_lut_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37679\,
            in2 => \N__26464\,
            in3 => \N__29657\,
            lcout => n11670,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1575_3_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39013\,
            in2 => \N__26455\,
            in3 => \N__34894\,
            lcout => n2415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1506_3_lut_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31969\,
            in2 => \N__32008\,
            in3 => \N__39104\,
            lcout => n2314,
            ltout => \n2314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1573_3_lut_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26581\,
            in2 => \N__26572\,
            in3 => \N__34895\,
            lcout => n2413,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1518_3_lut_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__31839\,
            in1 => \_gnd_net_\,
            in2 => \N__31816\,
            in3 => \N__39095\,
            lcout => n2326,
            ltout => \n2326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1585_3_lut_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34865\,
            in1 => \_gnd_net_\,
            in2 => \N__26569\,
            in3 => \N__26566\,
            lcout => n2425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1524_3_lut_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31521\,
            in2 => \N__31498\,
            in3 => \N__39096\,
            lcout => n2332,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1657_3_lut_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28996\,
            in2 => \N__35103\,
            in3 => \N__29025\,
            lcout => n2529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1592_3_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26554\,
            in2 => \N__26529\,
            in3 => \N__34864\,
            lcout => n2432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12853_4_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32039\,
            in1 => \N__31991\,
            in2 => \N__31953\,
            in3 => \N__26542\,
            lcout => n2247,
            ltout => \n2247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1525_3_lut_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__32161\,
            in1 => \N__31534\,
            in2 => \N__26536\,
            in3 => \_gnd_net_\,
            lcout => n2333,
            ltout => \n2333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10051_4_lut_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__26861\,
            in1 => \N__37512\,
            in2 => \N__26845\,
            in3 => \N__26842\,
            lcout => n11766,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1446_3_lut_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__36201\,
            in1 => \N__27105\,
            in2 => \N__26812\,
            in3 => \_gnd_net_\,
            lcout => n2222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9902_3_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27977\,
            in2 => \N__26797\,
            in3 => \N__26622\,
            lcout => OPEN,
            ltout => \n11616_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_99_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__26769\,
            in1 => \N__26739\,
            in2 => \N__26713\,
            in3 => \N__26693\,
            lcout => n13382,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12518_1_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35751\,
            lcout => n14990,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1321_3_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37599\,
            in1 => \N__26680\,
            in2 => \_gnd_net_\,
            in3 => \N__35871\,
            lcout => n2033,
            ltout => \n2033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1388_3_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26650\,
            in2 => \N__26638\,
            in3 => \N__36018\,
            lcout => n2132,
            ltout => \n2132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1455_3_lut_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26611\,
            in2 => \N__26599\,
            in3 => \N__36200\,
            lcout => n2231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1320_3_lut_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27193\,
            in2 => \N__27489\,
            in3 => \N__35872\,
            lcout => n2032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1379_3_lut_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27151\,
            in2 => \N__36045\,
            in3 => \N__27132\,
            lcout => n2123,
            ltout => \n2123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_96_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29370\,
            in1 => \N__29181\,
            in2 => \N__27091\,
            in3 => \N__29571\,
            lcout => OPEN,
            ltout => \n13746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_98_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27088\,
            in1 => \N__27596\,
            in2 => \N__27067\,
            in3 => \N__27064\,
            lcout => OPEN,
            ltout => \n13754_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_100_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27058\,
            in1 => \N__29676\,
            in2 => \N__27031\,
            in3 => \N__27028\,
            lcout => n13760,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1241_3_lut_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27006\,
            in1 => \_gnd_net_\,
            in2 => \N__35754\,
            in3 => \N__26986\,
            lcout => n1921,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1252_3_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28020\,
            in2 => \N__26947\,
            in3 => \N__35729\,
            lcout => n1932,
            ltout => \n1932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9971_4_lut_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__27482\,
            in1 => \N__37598\,
            in2 => \N__26911\,
            in3 => \N__26900\,
            lcout => n11686,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1249_3_lut_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27547\,
            in2 => \N__27277\,
            in3 => \N__35733\,
            lcout => n1929,
            ltout => \n1929_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_90_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27511\,
            in3 => \N__27438\,
            lcout => n14136,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1253_3_lut_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27502\,
            in1 => \N__32695\,
            in2 => \_gnd_net_\,
            in3 => \N__35728\,
            lcout => n1933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1250_3_lut_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27680\,
            in2 => \N__35753\,
            in3 => \N__27463\,
            lcout => n1930,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1237_3_lut_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27427\,
            in2 => \N__27415\,
            in3 => \N__35737\,
            lcout => n1917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1175_3_lut_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27361\,
            in2 => \N__27355\,
            in3 => \N__35611\,
            lcout => n1823,
            ltout => \n1823_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_84_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__27302\,
            in1 => \_gnd_net_\,
            in2 => \N__27280\,
            in3 => \N__27778\,
            lcout => OPEN,
            ltout => \n14126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_85_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__27276\,
            in1 => \N__27240\,
            in2 => \N__27214\,
            in3 => \N__27658\,
            lcout => n14128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1177_3_lut_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27199\,
            in1 => \_gnd_net_\,
            in2 => \N__35624\,
            in3 => \N__27886\,
            lcout => n1825,
            ltout => \n1825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_83_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27821\,
            in1 => \N__27797\,
            in2 => \N__27781\,
            in3 => \N__27725\,
            lcout => n14122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1180_3_lut_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27772\,
            in2 => \N__27751\,
            in3 => \N__35607\,
            lcout => n1828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9973_4_lut_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__32690\,
            in1 => \N__27710\,
            in2 => \N__27681\,
            in3 => \N__28019\,
            lcout => n11688,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1376_3_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27651\,
            in2 => \N__27622\,
            in3 => \N__36036\,
            lcout => n2120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i19_3_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33301\,
            in1 => \N__39465\,
            in2 => \_gnd_net_\,
            in3 => \N__29951\,
            lcout => n301,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29819\,
            lcout => n21_adj_645,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39309\,
            in3 => \_gnd_net_\,
            lcout => n29_adj_653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30064\,
            lcout => n4_adj_628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i17_3_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32971\,
            in1 => \N__39466\,
            in2 => \_gnd_net_\,
            in3 => \N__30140\,
            lcout => n303,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1185_3_lut_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28060\,
            in1 => \N__28044\,
            in2 => \_gnd_net_\,
            in3 => \N__35623\,
            lcout => n1833,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36287\,
            lcout => n8_adj_632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i13_3_lut_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33034\,
            in1 => \N__39396\,
            in2 => \_gnd_net_\,
            in3 => \N__29826\,
            lcout => n307,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i0_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38132\,
            in1 => \N__28446\,
            in2 => \_gnd_net_\,
            in3 => \N__27952\,
            lcout => h3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39394\,
            lcout => n2_adj_626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i14_3_lut_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39395\,
            in1 => \N__33022\,
            in2 => \_gnd_net_\,
            in3 => \N__38305\,
            lcout => n306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30106\,
            lcout => n6_adj_630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32182\,
            lcout => n22_adj_646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29976\,
            lcout => n16_adj_640,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10846_3_lut_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33427\,
            in2 => \N__30318\,
            in3 => \N__28210\,
            lcout => OPEN,
            ltout => \n13257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10847_3_lut_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__39444\,
            in1 => \_gnd_net_\,
            in2 => \N__28102\,
            in3 => \N__30068\,
            lcout => n830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2139_2_lut_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39443\,
            in2 => \_gnd_net_\,
            in3 => \N__33367\,
            lcout => n402,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30390\,
            in3 => \_gnd_net_\,
            lcout => n9_adj_633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i18_3_lut_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29977\,
            in1 => \N__33325\,
            in2 => \_gnd_net_\,
            in3 => \N__39445\,
            lcout => n302,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29955\,
            lcout => n15_adj_639,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_709_2_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30199\,
            in3 => \N__28069\,
            lcout => n2290,
            ltout => OPEN,
            carryin => \bfn_5_28_0_\,
            carryout => n12096,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_709_3_lut_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54599\,
            in2 => \N__30085\,
            in3 => \N__28066\,
            lcout => n2289,
            ltout => OPEN,
            carryin => n12096,
            carryout => n12097,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_709_4_lut_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30157\,
            in3 => \N__28063\,
            lcout => n2288,
            ltout => OPEN,
            carryin => n12097,
            carryout => n12098,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_709_5_lut_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30043\,
            in2 => \N__54977\,
            in3 => \N__28204\,
            lcout => n2287,
            ltout => OPEN,
            carryin => n12098,
            carryout => n12099,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_709_6_lut_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30223\,
            in3 => \N__28201\,
            lcout => n2286,
            ltout => OPEN,
            carryin => n12099,
            carryout => n12100,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_709_7_lut_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28198\,
            in3 => \N__28189\,
            lcout => n2285,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10850_3_lut_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33496\,
            in2 => \N__30317\,
            in3 => \N__28186\,
            lcout => OPEN,
            ltout => \n13261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10851_3_lut_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__39486\,
            in1 => \_gnd_net_\,
            in2 => \N__28180\,
            in3 => \N__30121\,
            lcout => n832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i3_3_lut_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32929\,
            in1 => \N__39497\,
            in2 => \_gnd_net_\,
            in3 => \N__32479\,
            lcout => n317,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i23_3_lut_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39496\,
            in1 => \N__33184\,
            in2 => \_gnd_net_\,
            in3 => \N__30037\,
            lcout => n297,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i1_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28147\,
            lcout => \reg_B_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32209\,
            lcout => n30_adj_654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i0_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28477\,
            lcout => \reg_B_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30036\,
            lcout => n11_adj_635,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10848_3_lut_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30307\,
            in2 => \N__33472\,
            in3 => \N__28426\,
            lcout => n13259,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29871\,
            lcout => n12_adj_636,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i837_3_lut_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36631\,
            in2 => \N__28713\,
            in3 => \N__28420\,
            lcout => n1325,
            ltout => \n1325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_71_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28382\,
            in1 => \N__28355\,
            in2 => \N__28339\,
            in3 => \N__28322\,
            lcout => n13734,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i22_3_lut_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33214\,
            in1 => \N__39534\,
            in2 => \_gnd_net_\,
            in3 => \N__29872\,
            lcout => n298,
            ltout => \n298_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9928_3_lut_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28278\,
            in2 => \N__28267\,
            in3 => \N__28259\,
            lcout => n11642,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i772_3_lut_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36540\,
            in2 => \N__28659\,
            in3 => \N__28243\,
            lcout => n1228,
            ltout => \n1228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_69_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28583\,
            in2 => \N__28717\,
            in3 => \N__28706\,
            lcout => n14078,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i708_3_lut_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__33928\,
            in1 => \N__30355\,
            in2 => \N__36958\,
            in3 => \_gnd_net_\,
            lcout => n1132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i705_3_lut_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30328\,
            in2 => \N__36959\,
            in3 => \N__33850\,
            lcout => n1129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i709_3_lut_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33948\,
            in2 => \N__30367\,
            in3 => \N__36941\,
            lcout => n1133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i771_3_lut_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__36539\,
            in1 => \_gnd_net_\,
            in2 => \N__30543\,
            in3 => \N__28603\,
            lcout => n1227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i774_3_lut_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36538\,
            in2 => \N__30449\,
            in3 => \N__28567\,
            lcout => n1230,
            ltout => \n1230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_70_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__28532\,
            in1 => \N__28511\,
            in2 => \N__28492\,
            in3 => \N__28489\,
            lcout => n13318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30418\,
            in3 => \_gnd_net_\,
            lcout => n10_adj_634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i703_3_lut_LC_5_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30586\,
            in2 => \N__30517\,
            in3 => \N__36948\,
            lcout => n1127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i701_3_lut_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30565\,
            in2 => \N__33778\,
            in3 => \N__36950\,
            lcout => n1125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i702_3_lut_LC_5_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30577\,
            in2 => \N__30493\,
            in3 => \N__36949\,
            lcout => n1126,
            ltout => \n1126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_63_LC_5_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30536\,
            in2 => \N__28768\,
            in3 => \N__28754\,
            lcout => n13994,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_2_lut_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32776\,
            in2 => \_gnd_net_\,
            in3 => \N__28732\,
            lcout => n2601,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => n12339,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_3_lut_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38985\,
            in2 => \N__53063\,
            in3 => \N__28729\,
            lcout => n2600,
            ltout => OPEN,
            carryin => n12339,
            carryout => n12340,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_4_lut_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31627\,
            in3 => \N__28726\,
            lcout => n2599,
            ltout => OPEN,
            carryin => n12340,
            carryout => n12341,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_5_lut_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53064\,
            in2 => \N__34461\,
            in3 => \N__28723\,
            lcout => n2598,
            ltout => OPEN,
            carryin => n12341,
            carryout => n12342,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_6_lut_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34297\,
            in3 => \N__28720\,
            lcout => n2597,
            ltout => OPEN,
            carryin => n12342,
            carryout => n12343,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_7_lut_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30619\,
            in3 => \N__28834\,
            lcout => n2596,
            ltout => OPEN,
            carryin => n12343,
            carryout => n12344,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_8_lut_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52985\,
            in2 => \N__30745\,
            in3 => \N__28831\,
            lcout => n2595,
            ltout => OPEN,
            carryin => n12344,
            carryout => n12345,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_9_lut_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53065\,
            in2 => \N__34414\,
            in3 => \N__28828\,
            lcout => n2594,
            ltout => OPEN,
            carryin => n12345,
            carryout => n12346,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_10_lut_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53007\,
            in2 => \N__34518\,
            in3 => \N__28825\,
            lcout => n2593,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => n12347,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_11_lut_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53014\,
            in2 => \N__30813\,
            in3 => \N__28822\,
            lcout => n2592,
            ltout => OPEN,
            carryin => n12347,
            carryout => n12348,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_12_lut_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53008\,
            in2 => \N__30853\,
            in3 => \N__28819\,
            lcout => n2591,
            ltout => OPEN,
            carryin => n12348,
            carryout => n12349,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_13_lut_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53015\,
            in2 => \N__30670\,
            in3 => \N__28816\,
            lcout => n2590,
            ltout => OPEN,
            carryin => n12349,
            carryout => n12350,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_14_lut_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53009\,
            in2 => \N__34353\,
            in3 => \N__28813\,
            lcout => n2589,
            ltout => OPEN,
            carryin => n12350,
            carryout => n12351,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_15_lut_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53016\,
            in2 => \N__37404\,
            in3 => \N__28810\,
            lcout => n2588,
            ltout => OPEN,
            carryin => n12351,
            carryout => n12352,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_16_lut_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53010\,
            in2 => \N__34609\,
            in3 => \N__28867\,
            lcout => n2587,
            ltout => OPEN,
            carryin => n12352,
            carryout => n12353,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_17_lut_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31108\,
            in2 => \N__53108\,
            in3 => \N__28864\,
            lcout => n2586,
            ltout => OPEN,
            carryin => n12353,
            carryout => n12354,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_18_lut_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31056\,
            in2 => \N__53662\,
            in3 => \N__28861\,
            lcout => n2585,
            ltout => OPEN,
            carryin => \bfn_6_16_0_\,
            carryout => n12355,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_19_lut_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53340\,
            in2 => \N__30783\,
            in3 => \N__28858\,
            lcout => n2584,
            ltout => OPEN,
            carryin => n12355,
            carryout => n12356,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_20_lut_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30993\,
            in2 => \N__53663\,
            in3 => \N__28855\,
            lcout => n2583,
            ltout => OPEN,
            carryin => n12356,
            carryout => n12357,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_21_lut_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31555\,
            in2 => \N__53347\,
            in3 => \N__28852\,
            lcout => n2582,
            ltout => OPEN,
            carryin => n12357,
            carryout => n12358,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_22_lut_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30971\,
            in2 => \N__53664\,
            in3 => \N__28843\,
            lcout => n2581,
            ltout => OPEN,
            carryin => n12358,
            carryout => n12359,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_23_lut_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34547\,
            in2 => \N__53348\,
            in3 => \N__28840\,
            lcout => n2580,
            ltout => OPEN,
            carryin => n12359,
            carryout => n12360,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_24_lut_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53124\,
            in2 => \N__31177\,
            in3 => \N__28837\,
            lcout => n2579,
            ltout => OPEN,
            carryin => n12360,
            carryout => n12361,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_25_lut_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__53125\,
            in1 => \N__30931\,
            in2 => \N__35157\,
            in3 => \N__29044\,
            lcout => n2610,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_2_lut_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37686\,
            in2 => \_gnd_net_\,
            in3 => \N__29041\,
            lcout => n2501,
            ltout => OPEN,
            carryin => \bfn_6_17_0_\,
            carryout => n12317,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_3_lut_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53177\,
            in2 => \N__29446\,
            in3 => \N__29038\,
            lcout => n2500,
            ltout => OPEN,
            carryin => n12317,
            carryout => n12318,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_4_lut_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29665\,
            in3 => \N__29035\,
            lcout => n2499,
            ltout => OPEN,
            carryin => n12318,
            carryout => n12319,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_5_lut_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53178\,
            in2 => \N__29424\,
            in3 => \N__29032\,
            lcout => n2498,
            ltout => OPEN,
            carryin => n12319,
            carryout => n12320,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_6_lut_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29029\,
            in3 => \N__28987\,
            lcout => n2497,
            ltout => OPEN,
            carryin => n12320,
            carryout => n12321,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_7_lut_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28984\,
            in3 => \N__28951\,
            lcout => n2496,
            ltout => OPEN,
            carryin => n12321,
            carryout => n12322,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_8_lut_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53736\,
            in2 => \N__28948\,
            in3 => \N__28915\,
            lcout => n2495,
            ltout => OPEN,
            carryin => n12322,
            carryout => n12323,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_9_lut_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53179\,
            in2 => \N__28911\,
            in3 => \N__28870\,
            lcout => n2494,
            ltout => OPEN,
            carryin => n12323,
            carryout => n12324,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_10_lut_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53349\,
            in2 => \N__31232\,
            in3 => \N__29128\,
            lcout => n2493,
            ltout => OPEN,
            carryin => \bfn_6_18_0_\,
            carryout => n12325,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_11_lut_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53356\,
            in2 => \N__30891\,
            in3 => \N__29125\,
            lcout => n2492,
            ltout => OPEN,
            carryin => n12325,
            carryout => n12326,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_12_lut_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53350\,
            in2 => \N__30699\,
            in3 => \N__29122\,
            lcout => n2491,
            ltout => OPEN,
            carryin => n12326,
            carryout => n12327,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_13_lut_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53357\,
            in2 => \N__31296\,
            in3 => \N__29113\,
            lcout => n2490,
            ltout => OPEN,
            carryin => n12327,
            carryout => n12328,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_14_lut_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53351\,
            in2 => \N__29110\,
            in3 => \N__29086\,
            lcout => n2489,
            ltout => OPEN,
            carryin => n12328,
            carryout => n12329,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_15_lut_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53358\,
            in2 => \N__29224\,
            in3 => \N__29083\,
            lcout => n2488,
            ltout => OPEN,
            carryin => n12329,
            carryout => n12330,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_16_lut_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53352\,
            in2 => \N__31137\,
            in3 => \N__29080\,
            lcout => n2487,
            ltout => OPEN,
            carryin => n12330,
            carryout => n12331,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_17_lut_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29077\,
            in2 => \N__53665\,
            in3 => \N__29047\,
            lcout => n2486,
            ltout => OPEN,
            carryin => n12331,
            carryout => n12332,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_18_lut_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29321\,
            in2 => \N__53666\,
            in3 => \N__29293\,
            lcout => n2485,
            ltout => OPEN,
            carryin => \bfn_6_19_0_\,
            carryout => n12333,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_19_lut_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53366\,
            in2 => \N__31032\,
            in3 => \N__29290\,
            lcout => n2484,
            ltout => OPEN,
            carryin => n12333,
            carryout => n12334,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_20_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31578\,
            in2 => \N__53667\,
            in3 => \N__29287\,
            lcout => n2483,
            ltout => OPEN,
            carryin => n12334,
            carryout => n12335,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_21_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29280\,
            in2 => \N__54676\,
            in3 => \N__29257\,
            lcout => n2482,
            ltout => OPEN,
            carryin => n12335,
            carryout => n12336,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_22_lut_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29781\,
            in2 => \N__53668\,
            in3 => \N__29254\,
            lcout => n2481,
            ltout => OPEN,
            carryin => n12336,
            carryout => n12337,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_23_lut_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31194\,
            in2 => \N__54677\,
            in3 => \N__29251\,
            lcout => n2480,
            ltout => OPEN,
            carryin => n12337,
            carryout => n12338,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_24_lut_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__53373\,
            in1 => \N__29247\,
            in2 => \N__35133\,
            in3 => \N__29227\,
            lcout => n2511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1648_3_lut_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29223\,
            in2 => \N__29191\,
            in3 => \N__35052\,
            lcout => n2520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1449_rep_27_3_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29182\,
            in2 => \N__36198\,
            in3 => \N__29149\,
            lcout => n2225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1448_3_lut_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29521\,
            in2 => \N__29506\,
            in3 => \N__36173\,
            lcout => n2224,
            ltout => \n2224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_101_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29473\,
            in3 => \N__31835\,
            lcout => OPEN,
            ltout => \n14174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_102_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31892\,
            in1 => \N__31793\,
            in2 => \N__29470\,
            in3 => \N__32498\,
            lcout => OPEN,
            ltout => \n14178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_103_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31730\,
            in1 => \N__31761\,
            in2 => \N__29467\,
            in3 => \N__31701\,
            lcout => n14184,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1660_3_lut_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__29455\,
            in1 => \_gnd_net_\,
            in2 => \N__29445\,
            in3 => \N__35067\,
            lcout => n2532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1658_3_lut_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29425\,
            in1 => \_gnd_net_\,
            in2 => \N__35102\,
            in3 => \N__29398\,
            lcout => n2530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1450_3_lut_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29389\,
            in2 => \N__29374\,
            in3 => \N__36169\,
            lcout => n2226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1661_3_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29338\,
            in1 => \N__37690\,
            in2 => \_gnd_net_\,
            in3 => \N__35075\,
            lcout => n2533,
            ltout => \n2533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9967_3_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32771\,
            in2 => \N__29326\,
            in3 => \N__31619\,
            lcout => OPEN,
            ltout => \n11682_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_121_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__30602\,
            in1 => \N__34280\,
            in2 => \N__29737\,
            in3 => \N__34443\,
            lcout => n13397,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1517_3_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31777\,
            in2 => \N__31801\,
            in3 => \N__39098\,
            lcout => n2325,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1374_3_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29725\,
            in2 => \N__29716\,
            in3 => \N__36044\,
            lcout => n2118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1659_3_lut_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29661\,
            in1 => \_gnd_net_\,
            in2 => \N__29641\,
            in3 => \N__35074\,
            lcout => n2531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1513_3_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31734\,
            in2 => \N__31714\,
            in3 => \N__39097\,
            lcout => n2321,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1380_3_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29625\,
            in2 => \N__29599\,
            in3 => \N__36037\,
            lcout => n2124,
            ltout => \n2124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1447_3_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29560\,
            in2 => \N__29545\,
            in3 => \N__36199\,
            lcout => n2223,
            ltout => \n2223_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1514_3_lut_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31744\,
            in1 => \_gnd_net_\,
            in2 => \N__29542\,
            in3 => \N__39119\,
            lcout => n2322,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1507_3_lut_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32046\,
            in2 => \N__39144\,
            in3 => \N__32017\,
            lcout => n2315,
            ltout => \n2315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1574_3_lut_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29797\,
            in2 => \N__29785\,
            in3 => \N__34931\,
            lcout => n2414,
            ltout => \n2414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1641_3_lut_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35105\,
            in1 => \_gnd_net_\,
            in2 => \N__29764\,
            in3 => \N__29761\,
            lcout => n2513,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12903_1_lut_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35104\,
            lcout => n15375,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12850_1_lut_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39143\,
            in3 => \_gnd_net_\,
            lcout => n15322,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i0_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32568\,
            in2 => \_gnd_net_\,
            in3 => \N__29752\,
            lcout => encoder0_position_0,
            ltout => OPEN,
            carryin => \bfn_6_23_0_\,
            carryout => \quad_counter0.n12623\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i1_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49765\,
            in2 => \N__32590\,
            in3 => \N__29749\,
            lcout => encoder0_position_1,
            ltout => OPEN,
            carryin => \quad_counter0.n12623\,
            carryout => \quad_counter0.n12624\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i2_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32475\,
            in2 => \N__49829\,
            in3 => \N__29746\,
            lcout => encoder0_position_2,
            ltout => OPEN,
            carryin => \quad_counter0.n12624\,
            carryout => \quad_counter0.n12625\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i3_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49769\,
            in2 => \N__32208\,
            in3 => \N__29743\,
            lcout => encoder0_position_3,
            ltout => OPEN,
            carryin => \quad_counter0.n12625\,
            carryout => \quad_counter0.n12626\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i4_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39302\,
            in2 => \N__49830\,
            in3 => \N__29740\,
            lcout => encoder0_position_4,
            ltout => OPEN,
            carryin => \quad_counter0.n12626\,
            carryout => \quad_counter0.n12627\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i5_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49773\,
            in2 => \N__32737\,
            in3 => \N__29848\,
            lcout => encoder0_position_5,
            ltout => OPEN,
            carryin => \quad_counter0.n12627\,
            carryout => \quad_counter0.n12628\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i6_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37772\,
            in2 => \N__49831\,
            in3 => \N__29845\,
            lcout => encoder0_position_6,
            ltout => OPEN,
            carryin => \quad_counter0.n12628\,
            carryout => \quad_counter0.n12629\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i7_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49777\,
            in2 => \N__37986\,
            in3 => \N__29842\,
            lcout => encoder0_position_7,
            ltout => OPEN,
            carryin => \quad_counter0.n12629\,
            carryout => \quad_counter0.n12630\,
            clk => \N__56040\,
            ce => \N__50436\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i8_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49832\,
            in2 => \N__32800\,
            in3 => \N__29839\,
            lcout => encoder0_position_8,
            ltout => OPEN,
            carryin => \bfn_6_24_0_\,
            carryout => \quad_counter0.n12631\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i9_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37712\,
            in2 => \N__49880\,
            in3 => \N__29836\,
            lcout => encoder0_position_9,
            ltout => OPEN,
            carryin => \quad_counter0.n12631\,
            carryout => \quad_counter0.n12632\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i10_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49836\,
            in2 => \N__37547\,
            in3 => \N__29833\,
            lcout => encoder0_position_10,
            ltout => OPEN,
            carryin => \quad_counter0.n12632\,
            carryout => \quad_counter0.n12633\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i11_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32181\,
            in2 => \N__49881\,
            in3 => \N__29830\,
            lcout => encoder0_position_11,
            ltout => OPEN,
            carryin => \quad_counter0.n12633\,
            carryout => \quad_counter0.n12634\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i12_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49840\,
            in2 => \N__29827\,
            in3 => \N__29803\,
            lcout => encoder0_position_12,
            ltout => OPEN,
            carryin => \quad_counter0.n12634\,
            carryout => \quad_counter0.n12635\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i13_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38297\,
            in2 => \N__49882\,
            in3 => \N__29800\,
            lcout => encoder0_position_13,
            ltout => OPEN,
            carryin => \quad_counter0.n12635\,
            carryout => \quad_counter0.n12636\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i14_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49844\,
            in2 => \N__37632\,
            in3 => \N__29986\,
            lcout => encoder0_position_14,
            ltout => OPEN,
            carryin => \quad_counter0.n12636\,
            carryout => \quad_counter0.n12637\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i15_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32715\,
            in2 => \N__49883\,
            in3 => \N__29983\,
            lcout => encoder0_position_15,
            ltout => OPEN,
            carryin => \quad_counter0.n12637\,
            carryout => \quad_counter0.n12638\,
            clk => \N__56043\,
            ce => \N__50437\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i16_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49848\,
            in2 => \N__30145\,
            in3 => \N__29980\,
            lcout => encoder0_position_16,
            ltout => OPEN,
            carryin => \bfn_6_25_0_\,
            carryout => \quad_counter0.n12639\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i17_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29975\,
            in2 => \N__49884\,
            in3 => \N__29959\,
            lcout => encoder0_position_17,
            ltout => OPEN,
            carryin => \quad_counter0.n12639\,
            carryout => \quad_counter0.n12640\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i18_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49852\,
            in2 => \N__29956\,
            in3 => \N__29932\,
            lcout => encoder0_position_18,
            ltout => OPEN,
            carryin => \quad_counter0.n12640\,
            carryout => \quad_counter0.n12641\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i19_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29922\,
            in2 => \N__49885\,
            in3 => \N__29908\,
            lcout => encoder0_position_19,
            ltout => OPEN,
            carryin => \quad_counter0.n12641\,
            carryout => \quad_counter0.n12642\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i20_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49856\,
            in2 => \N__29901\,
            in3 => \N__29875\,
            lcout => encoder0_position_20,
            ltout => OPEN,
            carryin => \quad_counter0.n12642\,
            carryout => \quad_counter0.n12643\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i21_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29865\,
            in2 => \N__49886\,
            in3 => \N__29851\,
            lcout => encoder0_position_21,
            ltout => OPEN,
            carryin => \quad_counter0.n12643\,
            carryout => \quad_counter0.n12644\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i22_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49860\,
            in2 => \N__30035\,
            in3 => \N__30013\,
            lcout => encoder0_position_22,
            ltout => OPEN,
            carryin => \quad_counter0.n12644\,
            carryout => \quad_counter0.n12645\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i23_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30407\,
            in2 => \N__49887\,
            in3 => \N__30010\,
            lcout => encoder0_position_23,
            ltout => OPEN,
            carryin => \quad_counter0.n12645\,
            carryout => \quad_counter0.n12646\,
            clk => \N__56047\,
            ce => \N__50432\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i24_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30389\,
            in2 => \N__49888\,
            in3 => \N__30007\,
            lcout => encoder0_position_24,
            ltout => OPEN,
            carryin => \bfn_6_26_0_\,
            carryout => \quad_counter0.n12647\,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i25_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49867\,
            in2 => \N__36297\,
            in3 => \N__30004\,
            lcout => encoder0_position_25,
            ltout => OPEN,
            carryin => \quad_counter0.n12647\,
            carryout => \quad_counter0.n12648\,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i26_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30271\,
            in2 => \N__49889\,
            in3 => \N__30001\,
            lcout => encoder0_position_26,
            ltout => OPEN,
            carryin => \quad_counter0.n12648\,
            carryout => \quad_counter0.n12649\,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i27_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49871\,
            in2 => \N__30120\,
            in3 => \N__29998\,
            lcout => encoder0_position_27,
            ltout => OPEN,
            carryin => \quad_counter0.n12649\,
            carryout => \quad_counter0.n12650\,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i28_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38257\,
            in2 => \N__49890\,
            in3 => \N__29995\,
            lcout => encoder0_position_28,
            ltout => OPEN,
            carryin => \quad_counter0.n12650\,
            carryout => \quad_counter0.n12651\,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i29_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49875\,
            in2 => \N__30075\,
            in3 => \N__29992\,
            lcout => encoder0_position_29,
            ltout => OPEN,
            carryin => \quad_counter0.n12651\,
            carryout => \quad_counter0.n12652\,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i30_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30245\,
            in2 => \N__49891\,
            in3 => \N__29989\,
            lcout => encoder0_position_30,
            ltout => OPEN,
            carryin => \quad_counter0.n12652\,
            carryout => \quad_counter0.n12653\,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_637__i31_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__39467\,
            in1 => \N__49879\,
            in2 => \_gnd_net_\,
            in3 => \N__30148\,
            lcout => encoder0_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56049\,
            ce => \N__50431\,
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30144\,
            lcout => n17_adj_641,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37628\,
            lcout => n19_adj_643,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30239\,
            lcout => n3_adj_627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32716\,
            lcout => n18_adj_642,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32799\,
            lcout => n25_adj_649,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37713\,
            lcout => n24_adj_648,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i28_3_lut_LC_6_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39442\,
            in2 => \N__30116\,
            in3 => \N__33491\,
            lcout => n175,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i1_3_lut_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__39476\,
            in1 => \_gnd_net_\,
            in2 => \N__32539\,
            in3 => \N__32572\,
            lcout => n319,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i30_3_lut_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39471\,
            in2 => \N__30076\,
            in3 => \N__33419\,
            lcout => n404,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_124_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30187\,
            in2 => \N__39529\,
            in3 => \N__33393\,
            lcout => OPEN,
            ltout => \n14170_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i500_4_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__33363\,
            in1 => \N__39475\,
            in2 => \N__30208\,
            in3 => \N__30205\,
            lcout => n828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i27_3_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30276\,
            in2 => \N__39528\,
            in3 => \N__33522\,
            lcout => n293,
            ltout => \n293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_65_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__33492\,
            in1 => \N__33420\,
            in2 => \N__30190\,
            in3 => \N__33462\,
            lcout => n5_adj_697,
            ltout => \n5_adj_697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_66_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33392\,
            in2 => \N__30181\,
            in3 => \N__33362\,
            lcout => n13254,
            ltout => \n13254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10852_3_lut_LC_6_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__33523\,
            in1 => \N__30178\,
            in2 => \N__30172\,
            in3 => \_gnd_net_\,
            lcout => n13263,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10849_3_lut_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38262\,
            in2 => \N__39531\,
            in3 => \N__30169\,
            lcout => n831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12294_3_lut_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39481\,
            in2 => \N__30277\,
            in3 => \N__30163\,
            lcout => n833,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i29_3_lut_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38261\,
            in2 => \N__39530\,
            in3 => \N__33461\,
            lcout => n174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i635_rep_55_3_lut_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34129\,
            in2 => \N__33793\,
            in3 => \N__34018\,
            lcout => n1027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10844_3_lut_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30319\,
            in2 => \N__33394\,
            in3 => \N__30286\,
            lcout => OPEN,
            ltout => \n13255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10845_3_lut_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__30249\,
            in1 => \_gnd_net_\,
            in2 => \N__30280\,
            in3 => \N__39485\,
            lcout => n829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30272\,
            lcout => n7_adj_631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i31_3_lut_LC_6_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39480\,
            in2 => \N__30250\,
            in3 => \N__33388\,
            lcout => n403,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9995_4_lut_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__34082\,
            in1 => \N__34064\,
            in2 => \N__33737\,
            in3 => \N__34034\,
            lcout => n11710,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9997_4_lut_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__36261\,
            in1 => \N__33572\,
            in2 => \N__34250\,
            in3 => \N__33707\,
            lcout => OPEN,
            ltout => \n11712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10107_4_lut_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__33656\,
            in1 => \N__33620\,
            in2 => \N__30214\,
            in3 => \N__33598\,
            lcout => n861,
            ltout => \n861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i573_3_lut_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__36262\,
            in1 => \N__33346\,
            in2 => \N__30211\,
            in3 => \_gnd_net_\,
            lcout => n933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i25_3_lut_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39532\,
            in2 => \N__33118\,
            in3 => \N__30391\,
            lcout => n295,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i569_3_lut_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33657\,
            in2 => \N__33637\,
            in3 => \N__34215\,
            lcout => n929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i568_3_lut_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__33607\,
            in1 => \N__33621\,
            in2 => \N__34224\,
            in3 => \_gnd_net_\,
            lcout => n928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i571_3_lut_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33708\,
            in2 => \N__33679\,
            in3 => \N__34214\,
            lcout => n931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_2_lut_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33947\,
            in2 => \_gnd_net_\,
            in3 => \N__30358\,
            lcout => n1101,
            ltout => OPEN,
            carryin => \bfn_6_31_0_\,
            carryout => n12114,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_3_lut_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55227\,
            in2 => \N__33927\,
            in3 => \N__30349\,
            lcout => n1100,
            ltout => OPEN,
            carryin => n12114,
            carryout => n12115,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_4_lut_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33970\,
            in3 => \N__30346\,
            lcout => n1099,
            ltout => OPEN,
            carryin => n12115,
            carryout => n12116,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_5_lut_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55228\,
            in2 => \N__33897\,
            in3 => \N__30331\,
            lcout => n1098,
            ltout => OPEN,
            carryin => n12116,
            carryout => n12117,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_6_lut_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33849\,
            in3 => \N__30322\,
            lcout => n1097,
            ltout => OPEN,
            carryin => n12117,
            carryout => n12118,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_7_lut_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33874\,
            in3 => \N__30589\,
            lcout => n1096,
            ltout => OPEN,
            carryin => n12118,
            carryout => n12119,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_8_lut_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55229\,
            in2 => \N__30516\,
            in3 => \N__30580\,
            lcout => n1095,
            ltout => OPEN,
            carryin => n12119,
            carryout => n12120,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_9_lut_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30488\,
            in2 => \N__55246\,
            in3 => \N__30571\,
            lcout => n1094,
            ltout => OPEN,
            carryin => n12120,
            carryout => n12121,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_10_lut_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__54598\,
            in1 => \N__33771\,
            in2 => \_gnd_net_\,
            in3 => \N__30568\,
            lcout => n1093,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i636_3_lut_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34171\,
            in2 => \N__33808\,
            in3 => \N__34015\,
            lcout => n1028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i704_3_lut_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33873\,
            in2 => \N__30559\,
            in3 => \N__36951\,
            lcout => n1128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12741_4_lut_LC_6_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30509\,
            in1 => \N__33770\,
            in2 => \N__30492\,
            in3 => \N__33826\,
            lcout => n1059,
            ltout => \n1059_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i707_3_lut_LC_6_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33969\,
            in1 => \_gnd_net_\,
            in2 => \N__30466\,
            in3 => \N__30463\,
            lcout => n1131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i24_3_lut_LC_6_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39533\,
            in2 => \N__33151\,
            in3 => \N__30417\,
            lcout => n296,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1718_3_lut_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30829\,
            in2 => \N__30669\,
            in3 => \N__38900\,
            lcout => n2622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12929_1_lut_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38930\,
            in3 => \_gnd_net_\,
            lcout => n15401,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1720_rep_19_3_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30823\,
            in2 => \N__30814\,
            in3 => \N__38849\,
            lcout => n2624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1712_3_lut_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30784\,
            in1 => \_gnd_net_\,
            in2 => \N__38898\,
            in3 => \N__30760\,
            lcout => n2616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1723_rep_21_3_lut_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30754\,
            in2 => \N__30744\,
            in3 => \N__38850\,
            lcout => n2627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1651_3_lut_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30712\,
            in2 => \N__30706\,
            in3 => \N__35101\,
            lcout => n2523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1711_3_lut_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30640\,
            in2 => \N__31000\,
            in3 => \N__38860\,
            lcout => n2615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1724_3_lut_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30628\,
            in2 => \N__38897\,
            in3 => \N__30618\,
            lcout => n2628,
            ltout => \n2628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_57_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38624\,
            in1 => \N__37425\,
            in2 => \N__31069\,
            in3 => \N__39254\,
            lcout => n14278,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1713_3_lut_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31066\,
            in2 => \N__38899\,
            in3 => \N__31060\,
            lcout => n2617,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1644_3_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31033\,
            in1 => \N__35084\,
            in2 => \_gnd_net_\,
            in3 => \N__31006\,
            lcout => n2516,
            ltout => \n2516_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_123_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30973\,
            in1 => \N__31547\,
            in2 => \N__30946\,
            in3 => \N__30943\,
            lcout => OPEN,
            ltout => \n13816_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12937_4_lut_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31169\,
            in1 => \N__34548\,
            in2 => \N__30934\,
            in3 => \N__30927\,
            lcout => n2544,
            ltout => \n2544_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1710_3_lut_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__30916\,
            in1 => \_gnd_net_\,
            in2 => \N__30907\,
            in3 => \N__31548\,
            lcout => n2614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1707_3_lut_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__31170\,
            in1 => \_gnd_net_\,
            in2 => \N__30904\,
            in3 => \N__38862\,
            lcout => n2611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1652_rep_61_3_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__30892\,
            in1 => \N__30859\,
            in2 => \N__35106\,
            in3 => \_gnd_net_\,
            lcout => n2524,
            ltout => \n2524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12344_3_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31321\,
            in2 => \N__31312\,
            in3 => \N__38861\,
            lcout => n2623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12377_3_lut_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32421\,
            in2 => \N__31309\,
            in3 => \N__34930\,
            lcout => n2423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1729_3_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31270\,
            in1 => \N__32775\,
            in2 => \_gnd_net_\,
            in3 => \N__38869\,
            lcout => n2633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1586_3_lut_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32358\,
            in2 => \N__31258\,
            in3 => \N__34919\,
            lcout => n2426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1640_3_lut_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31207\,
            in2 => \N__31201\,
            in3 => \N__35097\,
            lcout => n2512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1580_3_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32451\,
            in2 => \N__31156\,
            in3 => \N__34920\,
            lcout => n2420,
            ltout => \n2420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1647_3_lut_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31117\,
            in2 => \N__31111\,
            in3 => \N__35093\,
            lcout => n2519,
            ltout => \n2519_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1714_3_lut_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__38870\,
            in1 => \_gnd_net_\,
            in2 => \N__31084\,
            in3 => \N__31081\,
            lcout => n2618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1727_3_lut_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31623\,
            in2 => \N__31603\,
            in3 => \N__38868\,
            lcout => n2631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1643_3_lut_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31588\,
            in2 => \N__35109\,
            in3 => \N__31582\,
            lcout => n2515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_2_lut_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32148\,
            in2 => \_gnd_net_\,
            in3 => \N__31525\,
            lcout => n2301,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => n12276,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_3_lut_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53359\,
            in2 => \N__31522\,
            in3 => \N__31483\,
            lcout => n2300,
            ltout => OPEN,
            carryin => n12276,
            carryout => n12277,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_4_lut_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31480\,
            in3 => \N__31444\,
            lcout => n2299,
            ltout => OPEN,
            carryin => n12277,
            carryout => n12278,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_5_lut_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53360\,
            in2 => \N__31441\,
            in3 => \N__31405\,
            lcout => n2298,
            ltout => OPEN,
            carryin => n12278,
            carryout => n12279,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_6_lut_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31402\,
            in3 => \N__31366\,
            lcout => n2297,
            ltout => OPEN,
            carryin => n12279,
            carryout => n12280,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_7_lut_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31363\,
            in3 => \N__31324\,
            lcout => n2296,
            ltout => OPEN,
            carryin => n12280,
            carryout => n12281,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_8_lut_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53362\,
            in2 => \N__32511\,
            in3 => \N__31843\,
            lcout => n2295,
            ltout => OPEN,
            carryin => n12281,
            carryout => n12282,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_9_lut_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53361\,
            in2 => \N__31840\,
            in3 => \N__31804\,
            lcout => n2294,
            ltout => OPEN,
            carryin => n12282,
            carryout => n12283,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_10_lut_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54678\,
            in2 => \N__31800\,
            in3 => \N__31771\,
            lcout => n2293,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => n12284,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_11_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54240\,
            in2 => \N__31899\,
            in3 => \N__31768\,
            lcout => n2292,
            ltout => OPEN,
            carryin => n12284,
            carryout => n12285,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_12_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54679\,
            in2 => \N__31866\,
            in3 => \N__31765\,
            lcout => n2291,
            ltout => OPEN,
            carryin => n12285,
            carryout => n12286,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_13_lut_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54241\,
            in2 => \N__31762\,
            in3 => \N__31738\,
            lcout => n2290_adj_604,
            ltout => OPEN,
            carryin => n12286,
            carryout => n12287,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_14_lut_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31735\,
            in2 => \N__54727\,
            in3 => \N__31705\,
            lcout => n2289_adj_603,
            ltout => OPEN,
            carryin => n12287,
            carryout => n12288,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_15_lut_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31702\,
            in2 => \N__54996\,
            in3 => \N__31666\,
            lcout => n2288_adj_602,
            ltout => OPEN,
            carryin => n12288,
            carryout => n12289,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_16_lut_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31663\,
            in2 => \N__54728\,
            in3 => \N__32131\,
            lcout => n2287_adj_601,
            ltout => OPEN,
            carryin => n12289,
            carryout => n12290,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_17_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32128\,
            in2 => \N__54997\,
            in3 => \N__32098\,
            lcout => n2286_adj_600,
            ltout => OPEN,
            carryin => n12290,
            carryout => n12291,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_18_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32095\,
            in2 => \N__54077\,
            in3 => \N__32056\,
            lcout => n2285_adj_599,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => n12292,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_19_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53672\,
            in2 => \N__39196\,
            in3 => \N__32053\,
            lcout => n2284,
            ltout => OPEN,
            carryin => n12292,
            carryout => n12293,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_20_lut_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32050\,
            in2 => \N__54078\,
            in3 => \N__32011\,
            lcout => n2283,
            ltout => OPEN,
            carryin => n12293,
            carryout => n12294,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_21_lut_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32007\,
            in2 => \N__55161\,
            in3 => \N__31957\,
            lcout => n2282,
            ltout => OPEN,
            carryin => n12294,
            carryout => n12295,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_22_lut_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__53676\,
            in1 => \N__31954\,
            in2 => \N__34794\,
            in3 => \N__31924\,
            lcout => n2313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12376_3_lut_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31900\,
            in2 => \N__31876\,
            in3 => \N__39139\,
            lcout => n2324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1515_3_lut_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31867\,
            in2 => \N__39150\,
            in3 => \N__31849\,
            lcout => n2323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1519_3_lut_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32521\,
            in2 => \N__32512\,
            in3 => \N__39138\,
            lcout => n2327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32471\,
            lcout => n31_adj_655,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37776\,
            in1 => \N__32845\,
            in2 => \_gnd_net_\,
            in3 => \N__39548\,
            lcout => n313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_108_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32447\,
            in1 => \N__32411\,
            in2 => \N__32395\,
            in3 => \N__32348\,
            lcout => n14008,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32860\,
            in1 => \N__39549\,
            in2 => \_gnd_net_\,
            in3 => \N__32733\,
            lcout => n314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_107_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32318\,
            in1 => \N__32298\,
            in2 => \N__32277\,
            in3 => \N__32225\,
            lcout => n14006,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i4_3_lut_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39550\,
            in1 => \N__32896\,
            in2 => \_gnd_net_\,
            in3 => \N__32201\,
            lcout => n316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i12_3_lut_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33061\,
            in1 => \N__39547\,
            in2 => \_gnd_net_\,
            in3 => \N__32180\,
            lcout => n308,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39518\,
            in1 => \N__32947\,
            in2 => \_gnd_net_\,
            in3 => \N__32586\,
            lcout => n318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32812\,
            in1 => \N__32795\,
            in2 => \_gnd_net_\,
            in3 => \N__39517\,
            lcout => n311,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32732\,
            lcout => n28_adj_652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i16_3_lut_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32992\,
            in1 => \N__39516\,
            in2 => \_gnd_net_\,
            in3 => \N__32714\,
            lcout => n304,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37976\,
            lcout => n26_adj_650,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_109_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32662\,
            in1 => \N__32641\,
            in2 => \N__32620\,
            in3 => \N__32611\,
            lcout => n14014,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32585\,
            lcout => n32_adj_656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32564\,
            lcout => n33_adj_657,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32548\,
            in3 => \N__32524\,
            lcout => n33,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => n12575,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32956\,
            in3 => \N__32941\,
            lcout => n32,
            ltout => OPEN,
            carryin => n12575,
            carryout => n12576,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32938\,
            in2 => \_gnd_net_\,
            in3 => \N__32914\,
            lcout => n31,
            ltout => OPEN,
            carryin => n12576,
            carryout => n12577,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32911\,
            in3 => \N__32887\,
            lcout => n30,
            ltout => OPEN,
            carryin => n12577,
            carryout => n12578,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32884\,
            in3 => \N__32872\,
            lcout => n29,
            ltout => OPEN,
            carryin => n12578,
            carryout => n12579,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32869\,
            in3 => \N__32848\,
            lcout => n28,
            ltout => OPEN,
            carryin => n12579,
            carryout => n12580,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37753\,
            in3 => \N__32836\,
            lcout => n27,
            ltout => OPEN,
            carryin => n12580,
            carryout => n12581,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32833\,
            in3 => \N__32824\,
            lcout => n26,
            ltout => OPEN,
            carryin => n12581,
            carryout => n12582,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32821\,
            in3 => \N__32803\,
            lcout => n25,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => n12583,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33103\,
            in3 => \N__33094\,
            lcout => n24,
            ltout => OPEN,
            carryin => n12583,
            carryout => n12584,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33091\,
            in3 => \N__33076\,
            lcout => n23,
            ltout => OPEN,
            carryin => n12584,
            carryout => n12585,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33073\,
            in3 => \N__33052\,
            lcout => n22,
            ltout => OPEN,
            carryin => n12585,
            carryout => n12586,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33049\,
            in3 => \N__33025\,
            lcout => n21,
            ltout => OPEN,
            carryin => n12586,
            carryout => n12587,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38278\,
            in3 => \N__33013\,
            lcout => n20,
            ltout => OPEN,
            carryin => n12587,
            carryout => n12588,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33010\,
            in2 => \_gnd_net_\,
            in3 => \N__33004\,
            lcout => n19,
            ltout => OPEN,
            carryin => n12588,
            carryout => n12589,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33001\,
            in3 => \N__32983\,
            lcout => n18,
            ltout => OPEN,
            carryin => n12589,
            carryout => n12590,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32980\,
            in3 => \N__32959\,
            lcout => n17,
            ltout => OPEN,
            carryin => \bfn_7_27_0_\,
            carryout => n12591,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33337\,
            in3 => \N__33316\,
            lcout => n16,
            ltout => OPEN,
            carryin => n12591,
            carryout => n12592,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33313\,
            in3 => \N__33286\,
            lcout => n15,
            ltout => OPEN,
            carryin => n12592,
            carryout => n12593,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33283\,
            in3 => \N__33262\,
            lcout => n14,
            ltout => OPEN,
            carryin => n12593,
            carryout => n12594,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33259\,
            in3 => \N__33232\,
            lcout => n13,
            ltout => OPEN,
            carryin => n12594,
            carryout => n12595,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33229\,
            in3 => \N__33202\,
            lcout => n12,
            ltout => OPEN,
            carryin => n12595,
            carryout => n12596,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33199\,
            in3 => \N__33172\,
            lcout => n11,
            ltout => OPEN,
            carryin => n12596,
            carryout => n12597,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33169\,
            in3 => \N__33136\,
            lcout => n10,
            ltout => OPEN,
            carryin => n12597,
            carryout => n12598,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33133\,
            in3 => \N__33106\,
            lcout => n9,
            ltout => OPEN,
            carryin => \bfn_7_28_0_\,
            carryout => n12599,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33550\,
            in3 => \N__33535\,
            lcout => n8,
            ltout => OPEN,
            carryin => n12599,
            carryout => n12600,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33532\,
            in3 => \N__33514\,
            lcout => n7,
            ltout => OPEN,
            carryin => n12600,
            carryout => n12601,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33511\,
            in3 => \N__33475\,
            lcout => n6,
            ltout => OPEN,
            carryin => n12601,
            carryout => n12602,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38233\,
            in3 => \N__33445\,
            lcout => n5,
            ltout => OPEN,
            carryin => n12602,
            carryout => n12603,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33442\,
            in3 => \N__33406\,
            lcout => n4,
            ltout => OPEN,
            carryin => n12603,
            carryout => n12604,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33403\,
            in3 => \N__33373\,
            lcout => n3_adj_567,
            ltout => OPEN,
            carryin => n12604,
            carryout => n12605,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36438\,
            in3 => \N__33370\,
            lcout => n2_adj_568,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_2_lut_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36260\,
            in2 => \_gnd_net_\,
            in3 => \N__33340\,
            lcout => n901,
            ltout => OPEN,
            carryin => \bfn_7_29_0_\,
            carryout => n12101,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_3_lut_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55172\,
            in2 => \N__33573\,
            in3 => \N__33712\,
            lcout => n900,
            ltout => OPEN,
            carryin => n12101,
            carryout => n12102,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_4_lut_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33709\,
            in3 => \N__33670\,
            lcout => n899,
            ltout => OPEN,
            carryin => n12102,
            carryout => n12103,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_5_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55173\,
            in2 => \N__34251\,
            in3 => \N__33667\,
            lcout => n898,
            ltout => OPEN,
            carryin => n12103,
            carryout => n12104,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_6_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33664\,
            in3 => \N__33628\,
            lcout => n897,
            ltout => OPEN,
            carryin => n12104,
            carryout => n12105,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_7_lut_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33625\,
            in3 => \N__33601\,
            lcout => n896,
            ltout => OPEN,
            carryin => n12105,
            carryout => n12106,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_8_lut_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__55174\,
            in1 => \N__33597\,
            in2 => \N__34225\,
            in3 => \N__33583\,
            lcout => n927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i572_3_lut_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33580\,
            in2 => \N__33574\,
            in3 => \N__34219\,
            lcout => n932,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_2_lut_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34065\,
            in2 => \_gnd_net_\,
            in3 => \N__33553\,
            lcout => n1001,
            ltout => OPEN,
            carryin => \bfn_7_30_0_\,
            carryout => n12107,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_3_lut_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54594\,
            in2 => \N__34087\,
            in3 => \N__33820\,
            lcout => n1000,
            ltout => OPEN,
            carryin => n12107,
            carryout => n12108,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_4_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33738\,
            in3 => \N__33817\,
            lcout => n999,
            ltout => OPEN,
            carryin => n12108,
            carryout => n12109,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_5_lut_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54595\,
            in2 => \N__34039\,
            in3 => \N__33814\,
            lcout => n998,
            ltout => OPEN,
            carryin => n12109,
            carryout => n12110,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_6_lut_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34191\,
            in3 => \N__33811\,
            lcout => n997,
            ltout => OPEN,
            carryin => n12110,
            carryout => n12111,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_7_lut_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34170\,
            in3 => \N__33796\,
            lcout => n996,
            ltout => OPEN,
            carryin => n12111,
            carryout => n12112,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_8_lut_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54596\,
            in2 => \N__34128\,
            in3 => \N__33784\,
            lcout => n995,
            ltout => OPEN,
            carryin => n12112,
            carryout => n12113,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_9_lut_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54597\,
            in1 => \N__34014\,
            in2 => \N__34147\,
            in3 => \N__33781\,
            lcout => n1026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i637_3_lut_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33751\,
            in2 => \N__34192\,
            in3 => \N__34004\,
            lcout => n1029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i639_3_lut_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33745\,
            in2 => \N__34016\,
            in3 => \N__33739\,
            lcout => n1031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i570_3_lut_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34264\,
            in2 => \N__34255\,
            in3 => \N__34223\,
            lcout => n930,
            ltout => \n930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34174\,
            in3 => \N__34163\,
            lcout => OPEN,
            ltout => \n13726_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_7_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__34146\,
            in1 => \N__34121\,
            in2 => \N__34105\,
            in3 => \N__34102\,
            lcout => n960,
            ltout => \n960_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i640_3_lut_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34096\,
            in1 => \_gnd_net_\,
            in2 => \N__34090\,
            in3 => \N__34086\,
            lcout => n1032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i641_3_lut_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__34066\,
            in1 => \_gnd_net_\,
            in2 => \N__34048\,
            in3 => \N__34003\,
            lcout => n1033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i638_3_lut_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34038\,
            in2 => \N__34017\,
            in3 => \N__33976\,
            lcout => n1030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9932_3_lut_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33965\,
            in2 => \N__33949\,
            in3 => \N__33920\,
            lcout => OPEN,
            ltout => \n11646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_27_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__33890\,
            in1 => \N__33869\,
            in2 => \N__33853\,
            in3 => \N__33842\,
            lcout => n13323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i1_LC_7_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001100010000"
        )
    port map (
            in0 => \N__38088\,
            in1 => \N__38155\,
            in2 => \N__56353\,
            in3 => \N__38191\,
            lcout => commutation_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1726_3_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34462\,
            in1 => \N__34432\,
            in2 => \_gnd_net_\,
            in3 => \N__38936\,
            lcout => n2630,
            ltout => \n2630_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_60_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__37118\,
            in1 => \N__38674\,
            in2 => \N__34420\,
            in3 => \N__34363\,
            lcout => OPEN,
            ltout => \n14288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_61_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37472\,
            in1 => \N__38603\,
            in2 => \N__34417\,
            in3 => \N__37190\,
            lcout => n14294,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1722_3_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__34413\,
            in1 => \_gnd_net_\,
            in2 => \N__34393\,
            in3 => \N__38935\,
            lcout => n2626,
            ltout => \n2626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_58_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34638\,
            in1 => \N__34715\,
            in2 => \N__34378\,
            in3 => \N__34375\,
            lcout => OPEN,
            ltout => \n14280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_59_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37292\,
            in1 => \N__37019\,
            in2 => \N__34366\,
            in3 => \N__37353\,
            lcout => n14286,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1717_3_lut_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38908\,
            in2 => \N__34357\,
            in3 => \N__34321\,
            lcout => n2621,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1725_3_lut_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34309\,
            in2 => \N__38932\,
            in3 => \N__34296\,
            lcout => n2629,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1715_3_lut_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34608\,
            in2 => \N__34576\,
            in3 => \N__38909\,
            lcout => n2619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1708_3_lut_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34561\,
            in2 => \N__38933\,
            in3 => \N__34549\,
            lcout => n2612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12373_3_lut_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34693\,
            in2 => \N__42429\,
            in3 => \N__34717\,
            lcout => n2721,
            ltout => \n2721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12303_3_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40243\,
            in2 => \N__34522\,
            in3 => \N__47630\,
            lcout => n2820,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1721_rep_13_3_lut_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34519\,
            in2 => \N__34489\,
            in3 => \N__38907\,
            lcout => n2625,
            ltout => \n2625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12348_3_lut_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34627\,
            in2 => \N__34474\,
            in3 => \N__42391\,
            lcout => n2724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_2_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38775\,
            in2 => \_gnd_net_\,
            in3 => \N__34471\,
            lcout => n2701,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => n12362,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_3_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53482\,
            in2 => \N__38736\,
            in3 => \N__34468\,
            lcout => n2700,
            ltout => OPEN,
            carryin => n12362,
            carryout => n12363,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_4_lut_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38794\,
            in3 => \N__34465\,
            lcout => n2699,
            ltout => OPEN,
            carryin => n12363,
            carryout => n12364,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_5_lut_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53483\,
            in2 => \N__38703\,
            in3 => \N__34660\,
            lcout => n2698,
            ltout => OPEN,
            carryin => n12364,
            carryout => n12365,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_6_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37090\,
            in3 => \N__34657\,
            lcout => n2697,
            ltout => OPEN,
            carryin => n12365,
            carryout => n12366,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_7_lut_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37123\,
            in3 => \N__34654\,
            lcout => n2696,
            ltout => OPEN,
            carryin => n12366,
            carryout => n12367,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_8_lut_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53485\,
            in2 => \N__37054\,
            in3 => \N__34651\,
            lcout => n2695,
            ltout => OPEN,
            carryin => n12367,
            carryout => n12368,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_9_lut_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53484\,
            in2 => \N__37441\,
            in3 => \N__34648\,
            lcout => n2694,
            ltout => OPEN,
            carryin => n12368,
            carryout => n12369,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_10_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37144\,
            in2 => \N__53831\,
            in3 => \N__34645\,
            lcout => n2693,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => n12370,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_11_lut_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34642\,
            in2 => \N__53833\,
            in3 => \N__34618\,
            lcout => n2692,
            ltout => OPEN,
            carryin => n12370,
            carryout => n12371,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_12_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53496\,
            in2 => \N__38643\,
            in3 => \N__34615\,
            lcout => n2691,
            ltout => OPEN,
            carryin => n12371,
            carryout => n12372,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_13_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53489\,
            in2 => \N__39268\,
            in3 => \N__34612\,
            lcout => n2690,
            ltout => OPEN,
            carryin => n12372,
            carryout => n12373,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_14_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34716\,
            in2 => \N__53832\,
            in3 => \N__34684\,
            lcout => n2689,
            ltout => OPEN,
            carryin => n12373,
            carryout => n12374,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_15_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37297\,
            in2 => \N__53834\,
            in3 => \N__34681\,
            lcout => n2688,
            ltout => OPEN,
            carryin => n12374,
            carryout => n12375,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_16_lut_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53500\,
            in2 => \N__37360\,
            in3 => \N__34678\,
            lcout => n2687,
            ltout => OPEN,
            carryin => n12375,
            carryout => n12376,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_17_lut_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37026\,
            in2 => \N__53835\,
            in3 => \N__34675\,
            lcout => n2686,
            ltout => OPEN,
            carryin => n12376,
            carryout => n12377,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_18_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37191\,
            in2 => \N__53836\,
            in3 => \N__34672\,
            lcout => n2685,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => n12378,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_19_lut_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38610\,
            in2 => \N__53869\,
            in3 => \N__34669\,
            lcout => n2684,
            ltout => OPEN,
            carryin => n12378,
            carryout => n12379,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_20_lut_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53550\,
            in2 => \N__37483\,
            in3 => \N__34666\,
            lcout => n2683,
            ltout => OPEN,
            carryin => n12379,
            carryout => n12380,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_21_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38470\,
            in2 => \N__53870\,
            in3 => \N__34663\,
            lcout => n2682,
            ltout => OPEN,
            carryin => n12380,
            carryout => n12381,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_22_lut_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37245\,
            in2 => \N__53837\,
            in3 => \N__34732\,
            lcout => n2681,
            ltout => OPEN,
            carryin => n12381,
            carryout => n12382,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_23_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53510\,
            in2 => \N__38557\,
            in3 => \N__34729\,
            lcout => n2680,
            ltout => OPEN,
            carryin => n12382,
            carryout => n12383,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_24_lut_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42474\,
            in2 => \N__53838\,
            in3 => \N__34726\,
            lcout => n2679,
            ltout => OPEN,
            carryin => n12383,
            carryout => n12384,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_25_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38512\,
            in2 => \N__53871\,
            in3 => \N__34723\,
            lcout => n2678,
            ltout => OPEN,
            carryin => n12384,
            carryout => n12385,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_26_lut_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__53523\,
            in1 => \N__37330\,
            in2 => \N__35184\,
            in3 => \N__34720\,
            lcout => n2709,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12965_1_lut_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42443\,
            lcout => n15437,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1841_3_lut_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__47637\,
            in1 => \_gnd_net_\,
            in2 => \N__41572\,
            in3 => \N__40441\,
            lcout => n2809,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2067_3_lut_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44788\,
            in2 => \N__44764\,
            in3 => \N__49063\,
            lcout => n3131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2069_3_lut_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44854\,
            in2 => \N__49082\,
            in3 => \N__44892\,
            lcout => n3133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2042_3_lut_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45543\,
            in2 => \N__45517\,
            in3 => \N__49064\,
            lcout => n3106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2068_3_lut_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__44803\,
            in1 => \_gnd_net_\,
            in2 => \N__49081\,
            in3 => \N__44835\,
            lcout => n3132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10035_4_lut_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__51011\,
            in1 => \N__51176\,
            in2 => \N__51068\,
            in3 => \N__51110\,
            lcout => OPEN,
            ltout => \n11750_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_169_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__50978\,
            in1 => \N__50928\,
            in2 => \N__34750\,
            in3 => \N__39637\,
            lcout => OPEN,
            ltout => \n13900_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_170_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52214\,
            in1 => \N__51588\,
            in2 => \N__34747\,
            in3 => \N__51639\,
            lcout => n13906,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2136_3_lut_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51094\,
            in2 => \N__51117\,
            in3 => \N__50019\,
            lcout => n3232,
            ltout => \n3232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9943_3_lut_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42818\,
            in2 => \N__34744\,
            in3 => \N__42761\,
            lcout => n11658,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2134_3_lut_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__51012\,
            in1 => \N__50998\,
            in2 => \N__50070\,
            in3 => \_gnd_net_\,
            lcout => n3230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2129_3_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51556\,
            in2 => \N__51520\,
            in3 => \N__50013\,
            lcout => n3225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_171_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52174\,
            in1 => \N__52140\,
            in2 => \N__52093\,
            in3 => \N__34741\,
            lcout => OPEN,
            ltout => \n13912_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12689_4_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__52040\,
            in1 => \N__51992\,
            in2 => \N__34735\,
            in3 => \N__51930\,
            lcout => n3138,
            ltout => \n3138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2137_3_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__51181\,
            in1 => \_gnd_net_\,
            in2 => \N__34774\,
            in3 => \N__51139\,
            lcout => n3233,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2135_3_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51069\,
            in2 => \N__51040\,
            in3 => \N__50014\,
            lcout => n3231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2110_3_lut_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__52015\,
            in1 => \_gnd_net_\,
            in2 => \N__50069\,
            in3 => \N__52041\,
            lcout => n3206,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2133_3_lut_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50982\,
            in2 => \N__50950\,
            in3 => \N__50015\,
            lcout => n3229,
            ltout => \n3229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_154_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__42683\,
            in1 => \N__43094\,
            in2 => \N__34771\,
            in3 => \N__34768\,
            lcout => n13470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i0_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37876\,
            in1 => \N__36406\,
            in2 => \N__37924\,
            in3 => \N__34762\,
            lcout => encoder0_position_scaled_0,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => n12552,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i1_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__43587\,
            in1 => \N__49618\,
            in2 => \N__36469\,
            in3 => \N__34759\,
            lcout => encoder0_position_scaled_1,
            ltout => OPEN,
            carryin => n12552,
            carryout => n12553,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i2_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__51951\,
            in1 => \N__50032\,
            in2 => \N__36473\,
            in3 => \N__34756\,
            lcout => encoder0_position_scaled_2,
            ltout => OPEN,
            carryin => n12553,
            carryout => n12554,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i3_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45915\,
            in1 => \N__49080\,
            in2 => \N__36470\,
            in3 => \N__34753\,
            lcout => encoder0_position_scaled_3,
            ltout => OPEN,
            carryin => n12554,
            carryout => n12555,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i4_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39763\,
            in1 => \N__43009\,
            in2 => \N__36474\,
            in3 => \N__35197\,
            lcout => encoder0_position_scaled_4,
            ltout => OPEN,
            carryin => n12555,
            carryout => n12556,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i5_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__49201\,
            in1 => \N__49374\,
            in2 => \N__36471\,
            in3 => \N__35194\,
            lcout => encoder0_position_scaled_5,
            ltout => OPEN,
            carryin => n12556,
            carryout => n12557,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i6_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__42283\,
            in1 => \N__36416\,
            in2 => \N__47644\,
            in3 => \N__35191\,
            lcout => encoder0_position_scaled_6,
            ltout => OPEN,
            carryin => n12557,
            carryout => n12558,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i7_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35188\,
            in1 => \N__42448\,
            in2 => \N__36472\,
            in3 => \N__35167\,
            lcout => encoder0_position_scaled_7,
            ltout => OPEN,
            carryin => n12558,
            carryout => n12559,
            clk => \N__56055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i8_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35164\,
            in1 => \N__38944\,
            in2 => \N__36475\,
            in3 => \N__35140\,
            lcout => encoder0_position_scaled_8,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => n12560,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i9_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35137\,
            in1 => \N__35113\,
            in2 => \N__36479\,
            in3 => \N__34960\,
            lcout => encoder0_position_scaled_9,
            ltout => OPEN,
            carryin => n12560,
            carryout => n12561,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i10_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34957\,
            in1 => \N__34939\,
            in2 => \N__36476\,
            in3 => \N__34801\,
            lcout => encoder0_position_scaled_10,
            ltout => OPEN,
            carryin => n12561,
            carryout => n12562,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i11_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34798\,
            in1 => \N__39151\,
            in2 => \N__36480\,
            in3 => \N__34777\,
            lcout => encoder0_position_scaled_11,
            ltout => OPEN,
            carryin => n12562,
            carryout => n12563,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i12_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36235\,
            in1 => \N__36211\,
            in2 => \N__36477\,
            in3 => \N__36076\,
            lcout => encoder0_position_scaled_12,
            ltout => OPEN,
            carryin => n12563,
            carryout => n12564,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i13_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36073\,
            in1 => \N__36049\,
            in2 => \N__36481\,
            in3 => \N__35923\,
            lcout => encoder0_position_scaled_13,
            ltout => OPEN,
            carryin => n12564,
            carryout => n12565,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i14_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35920\,
            in1 => \N__35899\,
            in2 => \N__36478\,
            in3 => \N__35788\,
            lcout => encoder0_position_scaled_14,
            ltout => OPEN,
            carryin => n12565,
            carryout => n12566,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i15_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35785\,
            in1 => \N__35770\,
            in2 => \N__36482\,
            in3 => \N__35656\,
            lcout => encoder0_position_scaled_15,
            ltout => OPEN,
            carryin => n12566,
            carryout => n12567,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i16_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35653\,
            in1 => \N__35629\,
            in2 => \N__36483\,
            in3 => \N__35530\,
            lcout => encoder0_position_scaled_16,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => n12568,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i17_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__35527\,
            in1 => \N__36454\,
            in2 => \N__35503\,
            in3 => \N__35422\,
            lcout => encoder0_position_scaled_17,
            ltout => OPEN,
            carryin => n12568,
            carryout => n12569,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i18_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35419\,
            in1 => \N__35398\,
            in2 => \N__36484\,
            in3 => \N__35320\,
            lcout => encoder0_position_scaled_18,
            ltout => OPEN,
            carryin => n12569,
            carryout => n12570,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i19_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__35317\,
            in1 => \N__36458\,
            in2 => \N__35293\,
            in3 => \N__35200\,
            lcout => encoder0_position_scaled_19,
            ltout => OPEN,
            carryin => n12570,
            carryout => n12571,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i20_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36766\,
            in1 => \N__36745\,
            in2 => \N__36485\,
            in3 => \N__36673\,
            lcout => encoder0_position_scaled_20,
            ltout => OPEN,
            carryin => n12571,
            carryout => n12572,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i21_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__36670\,
            in1 => \N__36462\,
            in2 => \N__36646\,
            in3 => \N__36577\,
            lcout => encoder0_position_scaled_21,
            ltout => OPEN,
            carryin => n12572,
            carryout => n12573,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i22_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36574\,
            in1 => \N__36550\,
            in2 => \N__36486\,
            in3 => \N__36490\,
            lcout => encoder0_position_scaled_22,
            ltout => OPEN,
            carryin => n12573,
            carryout => n12574,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i23_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__36970\,
            in1 => \N__36904\,
            in2 => \N__36487\,
            in3 => \N__36316\,
            lcout => encoder0_position_scaled_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i18_1_lut_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36313\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n8_adj_562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i21_1_lut_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36307\,
            lcout => n5_adj_565,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i26_3_lut_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39542\,
            in2 => \N__36301\,
            in3 => \N__36271\,
            lcout => n294,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i2_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001100100010"
        )
    port map (
            in0 => \N__38150\,
            in1 => \N__38096\,
            in2 => \N__38203\,
            in3 => \N__56133\,
            lcout => commutation_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56061\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__38199\,
            in1 => \N__38148\,
            in2 => \_gnd_net_\,
            in3 => \N__38095\,
            lcout => \commutation_state_7__N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i24_1_lut_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36991\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_3_lut_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__38192\,
            in1 => \N__38149\,
            in2 => \_gnd_net_\,
            in3 => \N__38097\,
            lcout => n6_adj_592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_new_i0_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36985\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter0.a_new_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i16_3_lut_3_lut_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__40177\,
            in1 => \N__39848\,
            in2 => \_gnd_net_\,
            in3 => \N__52771\,
            lcout => n16_adj_614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i10_4_lut_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40176\,
            in1 => \N__44005\,
            in2 => \N__44035\,
            in3 => \N__40138\,
            lcout => \PWM.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12738_1_lut_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36966\,
            lcout => n15210,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12064_4_lut_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111000"
        )
    port map (
            in0 => \N__36832\,
            in1 => \N__36856\,
            in2 => \N__36793\,
            in3 => \N__36813\,
            lcout => OPEN,
            ltout => \n14536_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12065_3_lut_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__36772\,
            in1 => \_gnd_net_\,
            in2 => \N__36892\,
            in3 => \N__36889\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12063_4_lut_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011000100"
        )
    port map (
            in0 => \N__36855\,
            in1 => \N__36831\,
            in2 => \N__36814\,
            in3 => \N__36789\,
            lcout => n14535,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_62_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37244\,
            in1 => \N__38549\,
            in2 => \N__38468\,
            in3 => \N__37159\,
            lcout => n14300,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1789_3_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37153\,
            in2 => \N__42432\,
            in3 => \N__37143\,
            lcout => n2725,
            ltout => \n2725_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_51_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__42131\,
            in1 => \_gnd_net_\,
            in2 => \N__37129\,
            in3 => \N__44189\,
            lcout => OPEN,
            ltout => \n14040_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_53_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40365\,
            in1 => \N__40341\,
            in2 => \N__37126\,
            in3 => \N__37252\,
            lcout => n14048,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1792_3_lut_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37122\,
            in2 => \N__37102\,
            in3 => \N__42404\,
            lcout => n2728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1793_3_lut_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37086\,
            in2 => \N__42431\,
            in3 => \N__37072\,
            lcout => n2729,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1791_3_lut_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37063\,
            in2 => \N__37053\,
            in3 => \N__42405\,
            lcout => n2727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1782_3_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__42412\,
            in1 => \_gnd_net_\,
            in2 => \N__37027\,
            in3 => \N__37003\,
            lcout => n2718,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12350_3_lut_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__37440\,
            in1 => \_gnd_net_\,
            in2 => \N__37414\,
            in3 => \N__42395\,
            lcout => n2726,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1716_3_lut_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__37405\,
            in1 => \_gnd_net_\,
            in2 => \N__37375\,
            in3 => \N__38934\,
            lcout => n2620,
            ltout => \n2620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1783_3_lut_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37342\,
            in2 => \N__37333\,
            in3 => \N__42396\,
            lcout => n2719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12970_4_lut_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37326\,
            in1 => \N__38504\,
            in2 => \N__37306\,
            in3 => \N__42473\,
            lcout => n2643,
            ltout => \n2643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1784_3_lut_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__37296\,
            in1 => \_gnd_net_\,
            in2 => \N__37276\,
            in3 => \N__37273\,
            lcout => n2720,
            ltout => \n2720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_50_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41666\,
            in1 => \N__42173\,
            in2 => \N__37258\,
            in3 => \N__44486\,
            lcout => OPEN,
            ltout => \n14038_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_52_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40254\,
            in1 => \N__41879\,
            in2 => \N__37255\,
            in3 => \N__41951\,
            lcout => n14042,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1777_3_lut_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37246\,
            in2 => \N__42442\,
            in3 => \N__37213\,
            lcout => n2713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1781_3_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37201\,
            in2 => \N__37192\,
            in3 => \N__42422\,
            lcout => n2717,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37780\,
            lcout => n27_adj_651,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i10_3_lut_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39564\,
            in1 => \N__37735\,
            in2 => \_gnd_net_\,
            in3 => \N__37720\,
            lcout => n310,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i15_3_lut_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37654\,
            in1 => \N__39562\,
            in2 => \_gnd_net_\,
            in3 => \N__37636\,
            lcout => n305,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i11_3_lut_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39563\,
            in1 => \N__37570\,
            in2 => \_gnd_net_\,
            in3 => \N__37555\,
            lcout => n309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1779_3_lut_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37482\,
            in2 => \N__37456\,
            in3 => \N__42423\,
            lcout => n2715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_166_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51498\,
            in1 => \N__50855\,
            in2 => \N__51406\,
            in3 => \N__51548\,
            lcout => OPEN,
            ltout => \n13884_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_167_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51750\,
            in1 => \N__37813\,
            in2 => \N__37444\,
            in3 => \N__37807\,
            lcout => n13894,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2055_3_lut_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45422\,
            in2 => \N__45403\,
            in3 => \N__49069\,
            lcout => n3119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2053_3_lut_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45338\,
            in2 => \N__49084\,
            in3 => \N__45322\,
            lcout => n3117,
            ltout => \n3117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_165_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51842\,
            in1 => \N__50799\,
            in2 => \N__37816\,
            in3 => \N__51273\,
            lcout => n13888,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_164_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51310\,
            in1 => \N__51434\,
            in2 => \N__51348\,
            in3 => \N__51212\,
            lcout => n13886,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_2_lut_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47430\,
            in3 => \N__37801\,
            lcout => n3001,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => n12437,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_3_lut_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54699\,
            in2 => \N__47407\,
            in3 => \N__37798\,
            lcout => n3000,
            ltout => OPEN,
            carryin => n12437,
            carryout => n12438,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_4_lut_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47464\,
            in3 => \N__37795\,
            lcout => n2999,
            ltout => OPEN,
            carryin => n12438,
            carryout => n12439,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_5_lut_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54700\,
            in2 => \N__47350\,
            in3 => \N__37792\,
            lcout => n2998,
            ltout => OPEN,
            carryin => n12439,
            carryout => n12440,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_6_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47377\,
            in3 => \N__37789\,
            lcout => n2997,
            ltout => OPEN,
            carryin => n12440,
            carryout => n12441,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_7_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47314\,
            in3 => \N__37786\,
            lcout => n2996,
            ltout => OPEN,
            carryin => n12441,
            carryout => n12442,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_8_lut_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54702\,
            in2 => \N__44572\,
            in3 => \N__37783\,
            lcout => n2995,
            ltout => OPEN,
            carryin => n12442,
            carryout => n12443,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_9_lut_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54701\,
            in2 => \N__44629\,
            in3 => \N__37843\,
            lcout => n2994,
            ltout => OPEN,
            carryin => n12443,
            carryout => n12444,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_10_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44697\,
            in2 => \N__54321\,
            in3 => \N__37840\,
            lcout => n2993,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => n12445,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_11_lut_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53858\,
            in2 => \N__44950\,
            in3 => \N__37837\,
            lcout => n2992,
            ltout => OPEN,
            carryin => n12445,
            carryout => n12446,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_12_lut_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53860\,
            in2 => \N__44467\,
            in3 => \N__37834\,
            lcout => n2991,
            ltout => OPEN,
            carryin => n12446,
            carryout => n12447,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_13_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53859\,
            in2 => \N__44304\,
            in3 => \N__37831\,
            lcout => n2990,
            ltout => OPEN,
            carryin => n12447,
            carryout => n12448,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_14_lut_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53861\,
            in2 => \N__44545\,
            in3 => \N__37828\,
            lcout => n2989,
            ltout => OPEN,
            carryin => n12448,
            carryout => n12449,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_15_lut_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42117\,
            in2 => \N__54322\,
            in3 => \N__37825\,
            lcout => n2988,
            ltout => OPEN,
            carryin => n12449,
            carryout => n12450,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_16_lut_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53865\,
            in2 => \N__44667\,
            in3 => \N__37822\,
            lcout => n2987,
            ltout => OPEN,
            carryin => n12450,
            carryout => n12451,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_17_lut_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44601\,
            in2 => \N__54323\,
            in3 => \N__37819\,
            lcout => n2986,
            ltout => OPEN,
            carryin => n12451,
            carryout => n12452,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_18_lut_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42064\,
            in2 => \N__55185\,
            in3 => \N__37870\,
            lcout => n2985,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => n12453,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_19_lut_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55034\,
            in2 => \N__42091\,
            in3 => \N__37867\,
            lcout => n2984,
            ltout => OPEN,
            carryin => n12453,
            carryout => n12454,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_20_lut_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42531\,
            in2 => \N__55186\,
            in3 => \N__37864\,
            lcout => n2983,
            ltout => OPEN,
            carryin => n12454,
            carryout => n12455,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_21_lut_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42559\,
            in2 => \N__54603\,
            in3 => \N__37861\,
            lcout => n2982,
            ltout => OPEN,
            carryin => n12455,
            carryout => n12456,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_22_lut_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44919\,
            in2 => \N__55187\,
            in3 => \N__37858\,
            lcout => n2981,
            ltout => OPEN,
            carryin => n12456,
            carryout => n12457,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_23_lut_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42606\,
            in2 => \N__54604\,
            in3 => \N__37855\,
            lcout => n2980,
            ltout => OPEN,
            carryin => n12457,
            carryout => n12458,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_24_lut_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54115\,
            in2 => \N__40522\,
            in3 => \N__37852\,
            lcout => n2979,
            ltout => OPEN,
            carryin => n12458,
            carryout => n12459,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_25_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40545\,
            in2 => \N__54605\,
            in3 => \N__37849\,
            lcout => n2978,
            ltout => OPEN,
            carryin => n12459,
            carryout => n12460,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_26_lut_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47110\,
            in2 => \N__55188\,
            in3 => \N__37846\,
            lcout => n2977,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => n12461,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_27_lut_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42261\,
            in2 => \N__54976\,
            in3 => \N__37885\,
            lcout => n2976,
            ltout => OPEN,
            carryin => n12461,
            carryout => n12462,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_28_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40474\,
            in2 => \N__55189\,
            in3 => \N__37882\,
            lcout => n2975,
            ltout => OPEN,
            carryin => n12462,
            carryout => n12463,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_29_lut_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54593\,
            in1 => \N__39756\,
            in2 => \N__48766\,
            in3 => \N__37879\,
            lcout => n3006,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2111_3_lut_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52063\,
            in2 => \N__50071\,
            in3 => \N__52092\,
            lcout => n3207,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2112_3_lut_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52133\,
            in2 => \N__52114\,
            in3 => \N__50025\,
            lcout => n3208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2109_3_lut_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51970\,
            in2 => \N__50072\,
            in3 => \N__51996\,
            lcout => n3205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2114_3_lut_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__52224\,
            in1 => \_gnd_net_\,
            in2 => \N__52189\,
            in3 => \N__50024\,
            lcout => n3210,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12725_1_lut_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37923\,
            lcout => n15197,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16_4_lut_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__43078\,
            in1 => \N__42687\,
            in2 => \N__49606\,
            in3 => \N__43104\,
            lcout => n5_adj_713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9879_4_lut_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__42849\,
            in1 => \N__42822\,
            in2 => \N__42787\,
            in3 => \N__49569\,
            lcout => OPEN,
            ltout => \n11593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9941_4_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__49573\,
            in1 => \N__42745\,
            in2 => \N__37930\,
            in3 => \N__42765\,
            lcout => n11656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12686_1_lut_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50023\,
            lcout => n15158,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12691_1_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49607\,
            in3 => \_gnd_net_\,
            lcout => n15163,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2177_3_lut_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43642\,
            in1 => \N__43661\,
            in2 => \_gnd_net_\,
            in3 => \N__49577\,
            lcout => OPEN,
            ltout => \n59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12728_4_lut_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39715\,
            in1 => \N__43570\,
            in2 => \N__37927\,
            in3 => \N__39802\,
            lcout => n11838,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i1_1_lut_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37909\,
            lcout => n25_adj_545,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i16_1_lut_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37903\,
            lcout => n10_adj_560,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i13_1_lut_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37897\,
            lcout => n13_adj_557,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i3_1_lut_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37891\,
            lcout => n23_adj_547,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i5_1_lut_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38017\,
            lcout => n21_adj_549,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12457_2_lut_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55495\,
            in2 => \_gnd_net_\,
            in3 => \N__55469\,
            lcout => OPEN,
            ltout => \dti_N_333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101101111"
        )
    port map (
            in0 => \N__41066\,
            in1 => \N__56251\,
            in2 => \N__38011\,
            in3 => \N__41124\,
            lcout => n4828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i23_1_lut_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38008\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i8_3_lut_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38002\,
            in1 => \N__39558\,
            in2 => \_gnd_net_\,
            in3 => \N__37990\,
            lcout => n312,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i20_1_lut_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n6_adj_564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i22_1_lut_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37954\,
            lcout => n4_adj_566,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i14_1_lut_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37948\,
            lcout => n12_adj_558,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_154_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55506\,
            in2 => \_gnd_net_\,
            in3 => \N__55470\,
            lcout => dti,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56062\,
            ce => \N__37942\,
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38304\,
            lcout => n20_adj_644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38263\,
            lcout => n5_adj_629,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i10_1_lut_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38221\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n16_adj_554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i11_1_lut_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38212\,
            lcout => n15_adj_555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i0_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__38198\,
            in1 => \N__38154\,
            in2 => \_gnd_net_\,
            in3 => \N__38098\,
            lcout => commutation_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56065\,
            ce => \N__38041\,
            sr => \N__38029\
        );

    \LessThan_275_i13_2_lut_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41272\,
            in2 => \_gnd_net_\,
            in3 => \N__41164\,
            lcout => n13_adj_612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i23_2_lut_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41007\,
            in2 => \_gnd_net_\,
            in3 => \N__39947\,
            lcout => n23_adj_618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i11_4_lut_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40005\,
            in1 => \N__40974\,
            in2 => \N__39952\,
            in3 => \N__46766\,
            lcout => \PWM.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i41_2_lut_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41202\,
            in2 => \_gnd_net_\,
            in3 => \N__40004\,
            lcout => n41,
            ltout => \n41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12407_3_lut_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41203\,
            in1 => \_gnd_net_\,
            in2 => \N__38329\,
            in3 => \N__41362\,
            lcout => n40,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12243_4_lut_LC_10_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__38326\,
            in1 => \N__41386\,
            in2 => \N__38362\,
            in3 => \N__41743\,
            lcout => OPEN,
            ltout => \n14715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12394_4_lut_LC_10_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__38395\,
            in1 => \N__38371\,
            in2 => \N__38320\,
            in3 => \N__38317\,
            lcout => OPEN,
            ltout => \n14866_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.pwm_out_12_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43855\,
            in2 => \N__38311\,
            in3 => \N__44060\,
            lcout => pwm_out,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56069\,
            ce => 'H',
            sr => \N__41251\
        );

    \LessThan_275_i8_3_lut_3_lut_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__40993\,
            in1 => \N__41531\,
            in2 => \_gnd_net_\,
            in3 => \N__40804\,
            lcout => n8_adj_607,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i17_2_lut_LC_10_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40992\,
            in2 => \_gnd_net_\,
            in3 => \N__41530\,
            lcout => n17_adj_615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_10_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40044\,
            in1 => \N__40107\,
            in2 => \N__40063\,
            in3 => \N__40227\,
            lcout => OPEN,
            ltout => \n12_adj_598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_10_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40077\,
            in1 => \N__40212\,
            in2 => \N__38308\,
            in3 => \N__40092\,
            lcout => n4823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i45_2_lut_LC_10_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43950\,
            in2 => \_gnd_net_\,
            in3 => \N__40130\,
            lcout => n45,
            ltout => \n45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i24_3_lut_LC_10_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__43951\,
            in1 => \_gnd_net_\,
            in2 => \N__38422\,
            in3 => \N__38419\,
            lcout => n24_adj_619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i43_2_lut_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__39849\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40175\,
            lcout => n43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12371_3_lut_LC_10_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41828\,
            in1 => \N__41011\,
            in2 => \_gnd_net_\,
            in3 => \N__40948\,
            lcout => OPEN,
            ltout => \n14843_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12307_3_lut_LC_10_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41731\,
            in2 => \N__38413\,
            in3 => \N__41691\,
            lcout => n14779,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12239_2_lut_4_lut_LC_10_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__39850\,
            in1 => \N__52770\,
            in2 => \N__41350\,
            in3 => \N__40168\,
            lcout => OPEN,
            ltout => \n14711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12354_4_lut_LC_10_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__38410\,
            in1 => \N__38393\,
            in2 => \N__38404\,
            in3 => \N__38401\,
            lcout => OPEN,
            ltout => \n14826_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12392_4_lut_LC_10_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__38394\,
            in1 => \N__38347\,
            in2 => \N__38380\,
            in3 => \N__38377\,
            lcout => n14864,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12241_4_lut_LC_10_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__41692\,
            in1 => \N__41752\,
            in2 => \N__41833\,
            in3 => \N__38358\,
            lcout => n14713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1796_3_lut_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38341\,
            in2 => \N__42427\,
            in3 => \N__38737\,
            lcout => n2732,
            ltout => \n2732_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9951_3_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47678\,
            in2 => \N__38662\,
            in3 => \N__44381\,
            lcout => OPEN,
            ltout => \n11666_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_54_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__41852\,
            in1 => \N__41981\,
            in2 => \N__38659\,
            in3 => \N__44423\,
            lcout => n13403,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12346_3_lut_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38656\,
            in2 => \N__38644\,
            in3 => \N__42382\,
            lcout => n2723,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1780_3_lut_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38611\,
            in2 => \N__42428\,
            in3 => \N__38581\,
            lcout => n2716,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1797_3_lut_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38569\,
            in1 => \N__38776\,
            in2 => \_gnd_net_\,
            in3 => \N__42383\,
            lcout => n2733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1776_3_lut_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38550\,
            in2 => \N__38527\,
            in3 => \N__42390\,
            lcout => n2712,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1774_3_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38511\,
            in1 => \N__38482\,
            in2 => \_gnd_net_\,
            in3 => \N__42403\,
            lcout => n2710,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1848_3_lut_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40340\,
            in2 => \N__40318\,
            in3 => \N__47628\,
            lcout => n2816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1778_3_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38469\,
            in2 => \N__38437\,
            in3 => \N__42402\,
            lcout => n2714,
            ltout => \n2714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1845_3_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40300\,
            in2 => \N__39271\,
            in3 => \N__47627\,
            lcout => n2813,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12345_3_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39264\,
            in2 => \N__39238\,
            in3 => \N__42397\,
            lcout => n2722,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1794_3_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39223\,
            in2 => \N__42430\,
            in3 => \N__38704\,
            lcout => n2730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1795_3_lut_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38790\,
            in2 => \N__39211\,
            in3 => \N__42398\,
            lcout => n2731,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1508_3_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39195\,
            in2 => \N__39166\,
            in3 => \N__39149\,
            lcout => n2316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1728_3_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38989\,
            in2 => \N__38962\,
            in3 => \N__38931\,
            lcout => n2632,
            ltout => \n2632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10045_4_lut_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__38774\,
            in1 => \N__38729\,
            in2 => \N__38707\,
            in3 => \N__38696\,
            lcout => n11760,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1849_3_lut_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40378\,
            in2 => \N__40354\,
            in3 => \N__47629\,
            lcout => n2817,
            ltout => \n2817_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1916_3_lut_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48568\,
            in2 => \N__39601\,
            in3 => \N__49366\,
            lcout => n2916,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2000_3_lut_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__47406\,
            in1 => \N__39598\,
            in2 => \N__42997\,
            in3 => \_gnd_net_\,
            lcout => n3032,
            ltout => \n3032_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9945_3_lut_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__44888\,
            in1 => \_gnd_net_\,
            in2 => \N__39592\,
            in3 => \N__44819\,
            lcout => OPEN,
            ltout => \n11660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_31_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__45221\,
            in1 => \N__44732\,
            in2 => \N__39589\,
            in3 => \N__45180\,
            lcout => n13466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1986_3_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44602\,
            in2 => \N__39586\,
            in3 => \N__42960\,
            lcout => n3018,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1997_3_lut_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47376\,
            in2 => \N__42996\,
            in3 => \N__39574\,
            lcout => n3029,
            ltout => \n3029_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2064_3_lut_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45169\,
            in2 => \N__39568\,
            in3 => \N__49075\,
            lcout => n3128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i5_3_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__39565\,
            in1 => \N__39325\,
            in2 => \_gnd_net_\,
            in3 => \N__39313\,
            lcout => n315,
            ltout => \n315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2001_3_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39280\,
            in2 => \N__39274\,
            in3 => \N__42953\,
            lcout => n3033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1998_3_lut_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39652\,
            in2 => \N__42998\,
            in3 => \N__47346\,
            lcout => n3030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2063_3_lut_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__45150\,
            in1 => \N__45130\,
            in2 => \N__49043\,
            in3 => \_gnd_net_\,
            lcout => n3127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2051_3_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45247\,
            in2 => \N__45273\,
            in3 => \N__49000\,
            lcout => n3115,
            ltout => \n3115_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_168_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51670\,
            in2 => \N__39646\,
            in3 => \N__39643\,
            lcout => n13898,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1988_3_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42118\,
            in2 => \N__42999\,
            in3 => \N__39625\,
            lcout => n3020,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1987_3_lut_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39619\,
            in2 => \N__44668\,
            in3 => \N__42964\,
            lcout => n3019,
            ltout => \n3019_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2054_3_lut_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45364\,
            in2 => \N__39613\,
            in3 => \N__48995\,
            lcout => n3118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2060_3_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__48999\,
            in1 => \N__45028\,
            in2 => \N__45054\,
            in3 => \_gnd_net_\,
            lcout => n3124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1983_3_lut_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42532\,
            in2 => \N__39610\,
            in3 => \N__42971\,
            lcout => n3015,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1981_3_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__44920\,
            in1 => \N__39709\,
            in2 => \N__43001\,
            in3 => \_gnd_net_\,
            lcout => n3013,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2065_3_lut_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45225\,
            in2 => \N__45205\,
            in3 => \N__49019\,
            lcout => n3129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1984_3_lut_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39703\,
            in2 => \N__43000\,
            in3 => \N__42090\,
            lcout => n3016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1912_3_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48429\,
            in2 => \N__49375\,
            in3 => \N__48397\,
            lcout => n2912,
            ltout => \n2912_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1979_3_lut_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__42975\,
            in1 => \_gnd_net_\,
            in2 => \N__39697\,
            in3 => \N__39694\,
            lcout => n3011,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1975_3_lut_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40470\,
            in2 => \N__39688\,
            in3 => \N__42979\,
            lcout => n3007,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1980_3_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42607\,
            in2 => \N__39676\,
            in3 => \N__43003\,
            lcout => n3012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1976_3_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42262\,
            in2 => \N__39667\,
            in3 => \N__43005\,
            lcout => n3008,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2116_3_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51632\,
            in2 => \N__51613\,
            in3 => \N__50086\,
            lcout => n3212,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1978_3_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39658\,
            in2 => \N__40549\,
            in3 => \N__43004\,
            lcout => n3010,
            ltout => \n3010_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2045_3_lut_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45610\,
            in2 => \N__39766\,
            in3 => \N__49020\,
            lcout => n3109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12618_1_lut_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43002\,
            lcout => n15090,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2120_3_lut_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51775\,
            in2 => \N__51805\,
            in3 => \N__50085\,
            lcout => n3216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_157_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43478\,
            in1 => \N__43433\,
            in2 => \N__43401\,
            in3 => \N__39730\,
            lcout => OPEN,
            ltout => \n14392_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_160_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43337\,
            in1 => \N__43298\,
            in2 => \N__39745\,
            in3 => \N__49428\,
            lcout => n14398,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_155_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43199\,
            in1 => \N__43229\,
            in2 => \N__45802\,
            in3 => \N__39742\,
            lcout => OPEN,
            ltout => \n14380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_156_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43167\,
            in1 => \N__43132\,
            in2 => \N__39733\,
            in3 => \N__49930\,
            lcout => n14386,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12724_4_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__51909\,
            in1 => \N__43619\,
            in2 => \N__43668\,
            in3 => \N__39724\,
            lcout => n3237,
            ltout => \n3237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2176_3_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__43620\,
            in1 => \_gnd_net_\,
            in2 => \N__39718\,
            in3 => \N__43606\,
            lcout => n61,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_141_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__43453\,
            in1 => \N__43482\,
            in2 => \N__49608\,
            in3 => \N__40618\,
            lcout => OPEN,
            ltout => \n13856_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_142_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__43417\,
            in1 => \N__43441\,
            in2 => \N__39817\,
            in3 => \N__49581\,
            lcout => OPEN,
            ltout => \n13858_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_143_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__49582\,
            in1 => \N__43375\,
            in2 => \N__39814\,
            in3 => \N__43394\,
            lcout => OPEN,
            ltout => \n13860_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_144_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__43360\,
            in1 => \N__49583\,
            in2 => \N__39811\,
            in3 => \N__49429\,
            lcout => OPEN,
            ltout => \n13862_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_145_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__49584\,
            in1 => \N__43321\,
            in2 => \N__39808\,
            in3 => \N__43341\,
            lcout => OPEN,
            ltout => \n13864_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_146_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__43282\,
            in1 => \N__49585\,
            in2 => \N__39805\,
            in3 => \N__43302\,
            lcout => n13866,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i6_1_lut_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39796\,
            lcout => n20_adj_550,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i9_1_lut_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39784\,
            lcout => n17_adj_553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i12_1_lut_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39775\,
            lcout => n14_adj_556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i8_1_lut_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39877\,
            lcout => n18_adj_552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i22_1_lut_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46347\,
            lcout => n4_adj_570,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i2_1_lut_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39865\,
            lcout => n24_adj_546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_77_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__39892\,
            in1 => \N__56388\,
            in2 => \N__56174\,
            in3 => \N__55729\,
            lcout => n4_adj_698,
            ltout => \n4_adj_698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12245_2_lut_4_lut_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__41055\,
            in1 => \N__56254\,
            in2 => \N__39853\,
            in3 => \N__40722\,
            lcout => n14700,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12282_2_lut_4_lut_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__56252\,
            in1 => \N__41057\,
            in2 => \N__41140\,
            in3 => \N__43546\,
            lcout => n14692,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12293_2_lut_4_lut_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__41059\,
            in1 => \N__41132\,
            in2 => \N__40831\,
            in3 => \N__56256\,
            lcout => n14687,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12283_2_lut_4_lut_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__56253\,
            in1 => \N__41058\,
            in2 => \N__41141\,
            in3 => \N__43527\,
            lcout => n14693,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12281_2_lut_4_lut_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__41056\,
            in1 => \N__41131\,
            in2 => \N__40675\,
            in3 => \N__56255\,
            lcout => n14691,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i21_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55696\,
            in1 => \N__46348\,
            in2 => \_gnd_net_\,
            in3 => \N__43876\,
            lcout => pwm_setpoint_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i15_1_lut_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39928\,
            lcout => n11_adj_559,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i9_2_lut_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40797\,
            in2 => \_gnd_net_\,
            in3 => \N__39984\,
            lcout => n9_adj_608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i17_1_lut_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39916\,
            lcout => n9_adj_561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i0_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56250\,
            lcout => commutation_state_prev_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i19_1_lut_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39904\,
            lcout => n7_adj_563,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i2_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => commutation_state_prev_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.pwm_counter_635__i0_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46524\,
            in2 => \_gnd_net_\,
            in3 => \N__39886\,
            lcout => pwm_counter_0,
            ltout => OPEN,
            carryin => \bfn_11_29_0_\,
            carryout => \PWM.n12686\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i1_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46542\,
            in2 => \_gnd_net_\,
            in3 => \N__39883\,
            lcout => pwm_counter_1,
            ltout => OPEN,
            carryin => \PWM.n12686\,
            carryout => \PWM.n12687\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i2_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40782\,
            in2 => \_gnd_net_\,
            in3 => \N__39880\,
            lcout => pwm_counter_2,
            ltout => OPEN,
            carryin => \PWM.n12687\,
            carryout => \PWM.n12688\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i3_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40768\,
            in2 => \_gnd_net_\,
            in3 => \N__39988\,
            lcout => pwm_counter_3,
            ltout => OPEN,
            carryin => \PWM.n12688\,
            carryout => \PWM.n12689\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i4_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39985\,
            in2 => \_gnd_net_\,
            in3 => \N__39973\,
            lcout => pwm_counter_4,
            ltout => OPEN,
            carryin => \PWM.n12689\,
            carryout => \PWM.n12690\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i5_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41190\,
            in2 => \_gnd_net_\,
            in3 => \N__39970\,
            lcout => pwm_counter_5,
            ltout => OPEN,
            carryin => \PWM.n12690\,
            carryout => \PWM.n12691\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i6_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41169\,
            in2 => \_gnd_net_\,
            in3 => \N__39967\,
            lcout => pwm_counter_6,
            ltout => OPEN,
            carryin => \PWM.n12691\,
            carryout => \PWM.n12692\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i7_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47029\,
            in2 => \_gnd_net_\,
            in3 => \N__39964\,
            lcout => pwm_counter_7,
            ltout => OPEN,
            carryin => \PWM.n12692\,
            carryout => \PWM.n12693\,
            clk => \N__56070\,
            ce => 'H',
            sr => \N__41423\
        );

    \PWM.pwm_counter_635__i8_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41533\,
            in2 => \_gnd_net_\,
            in3 => \N__39961\,
            lcout => pwm_counter_8,
            ltout => OPEN,
            carryin => \bfn_11_30_0_\,
            carryout => \PWM.n12694\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i9_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41341\,
            in2 => \_gnd_net_\,
            in3 => \N__39958\,
            lcout => pwm_counter_9,
            ltout => OPEN,
            carryin => \PWM.n12694\,
            carryout => \PWM.n12695\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i10_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40975\,
            in2 => \_gnd_net_\,
            in3 => \N__39955\,
            lcout => pwm_counter_10,
            ltout => OPEN,
            carryin => \PWM.n12695\,
            carryout => \PWM.n12696\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i11_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39951\,
            in2 => \_gnd_net_\,
            in3 => \N__39931\,
            lcout => pwm_counter_11,
            ltout => OPEN,
            carryin => \PWM.n12696\,
            carryout => \PWM.n12697\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i12_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41712\,
            in2 => \_gnd_net_\,
            in3 => \N__40030\,
            lcout => pwm_counter_12,
            ltout => OPEN,
            carryin => \PWM.n12697\,
            carryout => \PWM.n12698\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i13_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46742\,
            in2 => \_gnd_net_\,
            in3 => \N__40027\,
            lcout => pwm_counter_13,
            ltout => OPEN,
            carryin => \PWM.n12698\,
            carryout => \PWM.n12699\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i14_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46767\,
            in2 => \_gnd_net_\,
            in3 => \N__40024\,
            lcout => pwm_counter_14,
            ltout => OPEN,
            carryin => \PWM.n12699\,
            carryout => \PWM.n12700\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i15_LC_11_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44030\,
            in2 => \_gnd_net_\,
            in3 => \N__40021\,
            lcout => pwm_counter_15,
            ltout => OPEN,
            carryin => \PWM.n12700\,
            carryout => \PWM.n12701\,
            clk => \N__56074\,
            ce => 'H',
            sr => \N__41440\
        );

    \PWM.pwm_counter_635__i16_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46828\,
            in2 => \_gnd_net_\,
            in3 => \N__40018\,
            lcout => pwm_counter_16,
            ltout => OPEN,
            carryin => \bfn_11_31_0_\,
            carryout => \PWM.n12702\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i17_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44270\,
            in2 => \_gnd_net_\,
            in3 => \N__40015\,
            lcout => pwm_counter_17,
            ltout => OPEN,
            carryin => \PWM.n12702\,
            carryout => \PWM.n12703\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i18_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44004\,
            in2 => \_gnd_net_\,
            in3 => \N__40012\,
            lcout => pwm_counter_18,
            ltout => OPEN,
            carryin => \PWM.n12703\,
            carryout => \PWM.n12704\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i19_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41401\,
            in2 => \_gnd_net_\,
            in3 => \N__40009\,
            lcout => pwm_counter_19,
            ltout => OPEN,
            carryin => \PWM.n12704\,
            carryout => \PWM.n12705\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i20_LC_11_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40006\,
            in2 => \_gnd_net_\,
            in3 => \N__39991\,
            lcout => pwm_counter_20,
            ltout => OPEN,
            carryin => \PWM.n12705\,
            carryout => \PWM.n12706\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i21_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40169\,
            in2 => \_gnd_net_\,
            in3 => \N__40141\,
            lcout => pwm_counter_21,
            ltout => OPEN,
            carryin => \PWM.n12706\,
            carryout => \PWM.n12707\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i22_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40134\,
            in2 => \_gnd_net_\,
            in3 => \N__40114\,
            lcout => pwm_counter_22,
            ltout => OPEN,
            carryin => \PWM.n12707\,
            carryout => \PWM.n12708\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i23_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44062\,
            in2 => \_gnd_net_\,
            in3 => \N__40111\,
            lcout => pwm_counter_23,
            ltout => OPEN,
            carryin => \PWM.n12708\,
            carryout => \PWM.n12709\,
            clk => \N__56077\,
            ce => 'H',
            sr => \N__41429\
        );

    \PWM.pwm_counter_635__i24_LC_11_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40108\,
            in2 => \_gnd_net_\,
            in3 => \N__40096\,
            lcout => pwm_counter_24,
            ltout => OPEN,
            carryin => \bfn_11_32_0_\,
            carryout => \PWM.n12710\,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \PWM.pwm_counter_635__i25_LC_11_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40093\,
            in2 => \_gnd_net_\,
            in3 => \N__40081\,
            lcout => pwm_counter_25,
            ltout => OPEN,
            carryin => \PWM.n12710\,
            carryout => \PWM.n12711\,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \PWM.pwm_counter_635__i26_LC_11_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40078\,
            in2 => \_gnd_net_\,
            in3 => \N__40066\,
            lcout => pwm_counter_26,
            ltout => OPEN,
            carryin => \PWM.n12711\,
            carryout => \PWM.n12712\,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \PWM.pwm_counter_635__i27_LC_11_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40062\,
            in2 => \_gnd_net_\,
            in3 => \N__40048\,
            lcout => pwm_counter_27,
            ltout => OPEN,
            carryin => \PWM.n12712\,
            carryout => \PWM.n12713\,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \PWM.pwm_counter_635__i28_LC_11_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40045\,
            in2 => \_gnd_net_\,
            in3 => \N__40033\,
            lcout => pwm_counter_28,
            ltout => OPEN,
            carryin => \PWM.n12713\,
            carryout => \PWM.n12714\,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \PWM.pwm_counter_635__i29_LC_11_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40228\,
            in2 => \_gnd_net_\,
            in3 => \N__40216\,
            lcout => pwm_counter_29,
            ltout => OPEN,
            carryin => \PWM.n12714\,
            carryout => \PWM.n12715\,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \PWM.pwm_counter_635__i30_LC_11_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40213\,
            in2 => \_gnd_net_\,
            in3 => \N__40201\,
            lcout => pwm_counter_30,
            ltout => OPEN,
            carryin => \PWM.n12715\,
            carryout => \PWM.n12716\,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \PWM.pwm_counter_635__i31_LC_11_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41475\,
            in2 => \_gnd_net_\,
            in3 => \N__40198\,
            lcout => pwm_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56081\,
            ce => 'H',
            sr => \N__41436\
        );

    \encoder0_position_31__I_0_add_1838_2_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47683\,
            in2 => \_gnd_net_\,
            in3 => \N__40195\,
            lcout => n2801,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => n12386,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_3_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53560\,
            in2 => \N__44385\,
            in3 => \N__40192\,
            lcout => n2800,
            ltout => OPEN,
            carryin => n12386,
            carryout => n12387,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_4_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44346\,
            in3 => \N__40189\,
            lcout => n2799,
            ltout => OPEN,
            carryin => n12387,
            carryout => n12388,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_5_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53561\,
            in2 => \N__41985\,
            in3 => \N__40186\,
            lcout => n2798,
            ltout => OPEN,
            carryin => n12388,
            carryout => n12389,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_6_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41856\,
            in3 => \N__40183\,
            lcout => n2797,
            ltout => OPEN,
            carryin => n12389,
            carryout => n12390,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_7_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44430\,
            in3 => \N__40180\,
            lcout => n2796,
            ltout => OPEN,
            carryin => n12390,
            carryout => n12391,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_8_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53569\,
            in2 => \N__41962\,
            in3 => \N__40282\,
            lcout => n2795,
            ltout => OPEN,
            carryin => n12391,
            carryout => n12392,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_9_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53562\,
            in2 => \N__44193\,
            in3 => \N__40279\,
            lcout => n2794,
            ltout => OPEN,
            carryin => n12392,
            carryout => n12393,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_10_lut_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53839\,
            in2 => \N__44499\,
            in3 => \N__40276\,
            lcout => n2793,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => n12394,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_11_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53563\,
            in2 => \N__41641\,
            in3 => \N__40273\,
            lcout => n2792,
            ltout => OPEN,
            carryin => n12394,
            carryout => n12395,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_12_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53840\,
            in2 => \N__42184\,
            in3 => \N__40270\,
            lcout => n2791,
            ltout => OPEN,
            carryin => n12395,
            carryout => n12396,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_13_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53564\,
            in2 => \N__41673\,
            in3 => \N__40267\,
            lcout => n2790,
            ltout => OPEN,
            carryin => n12396,
            carryout => n12397,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_14_lut_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53841\,
            in2 => \N__41886\,
            in3 => \N__40264\,
            lcout => n2789,
            ltout => OPEN,
            carryin => n12397,
            carryout => n12398,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_15_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53565\,
            in2 => \N__40261\,
            in3 => \N__40234\,
            lcout => n2788,
            ltout => OPEN,
            carryin => n12398,
            carryout => n12399,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_16_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41919\,
            in2 => \N__53877\,
            in3 => \N__40231\,
            lcout => n2787,
            ltout => OPEN,
            carryin => n12399,
            carryout => n12400,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_17_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42138\,
            in2 => \N__54308\,
            in3 => \N__40381\,
            lcout => n2786,
            ltout => OPEN,
            carryin => n12400,
            carryout => n12401,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_18_lut_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40377\,
            in2 => \N__54336\,
            in3 => \N__40345\,
            lcout => n2785,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => n12402,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_19_lut_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40342\,
            in2 => \N__54767\,
            in3 => \N__40309\,
            lcout => n2784,
            ltout => OPEN,
            carryin => n12402,
            carryout => n12403,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_20_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44167\,
            in2 => \N__54337\,
            in3 => \N__40306\,
            lcout => n2783,
            ltout => OPEN,
            carryin => n12403,
            carryout => n12404,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_21_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44111\,
            in2 => \N__54768\,
            in3 => \N__40303\,
            lcout => n2782,
            ltout => OPEN,
            carryin => n12404,
            carryout => n12405,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_22_lut_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41589\,
            in2 => \N__54338\,
            in3 => \N__40294\,
            lcout => n2781,
            ltout => OPEN,
            carryin => n12405,
            carryout => n12406,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_23_lut_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42227\,
            in2 => \N__54769\,
            in3 => \N__40291\,
            lcout => n2780,
            ltout => OPEN,
            carryin => n12406,
            carryout => n12407,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_24_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44250\,
            in2 => \N__54339\,
            in3 => \N__40288\,
            lcout => n2779,
            ltout => OPEN,
            carryin => n12407,
            carryout => n12408,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_25_lut_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53890\,
            in2 => \N__42309\,
            in3 => \N__40285\,
            lcout => n2778,
            ltout => OPEN,
            carryin => n12408,
            carryout => n12409,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_26_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41567\,
            in2 => \N__54770\,
            in3 => \N__40429\,
            lcout => n2777,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => n12410,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_27_lut_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53891\,
            in1 => \N__42273\,
            in2 => \N__42028\,
            in3 => \N__40426\,
            lcout => n2808,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2043_3_lut_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45588\,
            in2 => \N__45562\,
            in3 => \N__49074\,
            lcout => n3107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1911_3_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48377\,
            in2 => \N__48355\,
            in3 => \N__49367\,
            lcout => n2911,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1985_3_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40423\,
            in2 => \N__42063\,
            in3 => \N__42980\,
            lcout => n3017,
            ltout => \n3017_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2052_3_lut_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45289\,
            in2 => \N__40411\,
            in3 => \N__49073\,
            lcout => n3116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1977_3_lut_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__47103\,
            in1 => \_gnd_net_\,
            in2 => \N__42993\,
            in3 => \N__40408\,
            lcout => n3009,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1993_3_lut_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__44698\,
            in1 => \_gnd_net_\,
            in2 => \N__40396\,
            in3 => \N__42940\,
            lcout => n3025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_41_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44912\,
            in1 => \N__42594\,
            in2 => \N__47275\,
            in3 => \N__42505\,
            lcout => OPEN,
            ltout => \n13948_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_42_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40533\,
            in1 => \N__40518\,
            in2 => \N__40507\,
            in3 => \N__47102\,
            lcout => OPEN,
            ltout => \n13954_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12622_4_lut_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42248\,
            in1 => \N__48759\,
            in2 => \N__40504\,
            in3 => \N__40466\,
            lcout => n2940,
            ltout => \n2940_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1999_3_lut_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40501\,
            in1 => \_gnd_net_\,
            in2 => \N__40492\,
            in3 => \N__47460\,
            lcout => n3031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1996_3_lut_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47313\,
            in2 => \N__40489\,
            in3 => \N__42941\,
            lcout => n3028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_33_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45705\,
            in1 => \N__49463\,
            in2 => \N__45668\,
            in3 => \N__40561\,
            lcout => OPEN,
            ltout => \n14340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_34_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45621\,
            in1 => \N__49173\,
            in2 => \N__40477\,
            in3 => \N__43015\,
            lcout => n14344,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1908_3_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__48823\,
            in1 => \_gnd_net_\,
            in2 => \N__48863\,
            in3 => \N__49371\,
            lcout => n2908,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12655_4_lut_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45578\,
            in1 => \N__45533\,
            in2 => \N__45940\,
            in3 => \N__40450\,
            lcout => n3039,
            ltout => \n3039_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2059_3_lut_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44992\,
            in2 => \N__40444\,
            in3 => \N__45012\,
            lcout => n3123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_32_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49118\,
            in1 => \N__45303\,
            in2 => \N__42193\,
            in3 => \N__40570\,
            lcout => n14334,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12651_1_lut_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49079\,
            in3 => \_gnd_net_\,
            lcout => n15123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2047_3_lut_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__45670\,
            in1 => \N__45646\,
            in2 => \N__49039\,
            in3 => \_gnd_net_\,
            lcout => n3111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2057_3_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45495\,
            in2 => \N__45475\,
            in3 => \N__48980\,
            lcout => n3121,
            ltout => \n3121_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2124_3_lut_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51289\,
            in2 => \N__40555\,
            in3 => \N__50073\,
            lcout => n3220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2049_3_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45721\,
            in2 => \N__45736\,
            in3 => \N__48981\,
            lcout => n3113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2121_3_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51852\,
            in2 => \N__51826\,
            in3 => \N__50077\,
            lcout => n3217,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2127_3_lut_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__51418\,
            in1 => \_gnd_net_\,
            in2 => \N__50105\,
            in3 => \N__51444\,
            lcout => n3223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2048_3_lut_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45682\,
            in2 => \N__49040\,
            in3 => \N__45704\,
            lcout => n3112,
            ltout => \n3112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2115_3_lut_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50078\,
            in1 => \_gnd_net_\,
            in2 => \N__40552\,
            in3 => \N__51571\,
            lcout => n3211,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2195_3_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45766\,
            in2 => \N__43042\,
            in3 => \N__49563\,
            lcout => OPEN,
            ltout => \n23_adj_707_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_132_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__49565\,
            in1 => \N__43264\,
            in2 => \N__40600\,
            in3 => \N__45871\,
            lcout => n13828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2194_3_lut_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46134\,
            in2 => \N__43030\,
            in3 => \N__49564\,
            lcout => OPEN,
            ltout => \n25_adj_708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_133_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__49566\,
            in1 => \N__45837\,
            in2 => \N__40597\,
            in3 => \N__43249\,
            lcout => n13826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_131_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__40612\,
            in1 => \N__43054\,
            in2 => \N__49402\,
            in3 => \N__49567\,
            lcout => OPEN,
            ltout => \n13832_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_135_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__49568\,
            in1 => \N__43183\,
            in2 => \N__40594\,
            in3 => \N__43203\,
            lcout => OPEN,
            ltout => \n13840_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_136_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40591\,
            in1 => \N__40585\,
            in2 => \N__40579\,
            in3 => \N__48652\,
            lcout => n13846,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i5_1_lut_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46002\,
            lcout => n21_adj_587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_137_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__43171\,
            in1 => \N__43141\,
            in2 => \N__49605\,
            in3 => \N__40576\,
            lcout => OPEN,
            ltout => \n13848_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_138_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__43501\,
            in1 => \N__43131\,
            in2 => \N__40645\,
            in3 => \N__49561\,
            lcout => OPEN,
            ltout => \n13850_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_139_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__40606\,
            in1 => \N__40642\,
            in2 => \N__40633\,
            in3 => \N__40630\,
            lcout => OPEN,
            ltout => \n13852_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_140_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__49929\,
            in1 => \N__43492\,
            in2 => \N__40621\,
            in3 => \N__49562\,
            lcout => n13854,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2126_3_lut_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51395\,
            in2 => \N__51367\,
            in3 => \N__50106\,
            lcout => n3222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2188_3_lut_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43216\,
            in2 => \N__43240\,
            in3 => \N__49554\,
            lcout => n37_adj_710,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2203_3_lut_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42706\,
            in2 => \N__49604\,
            in3 => \N__42727\,
            lcout => n7_adj_703,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2118_3_lut_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__50107\,
            in1 => \N__51685\,
            in2 => \N__51715\,
            in3 => \_gnd_net_\,
            lcout => n3214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12280_2_lut_4_lut_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000100"
        )
    port map (
            in0 => \N__56277\,
            in1 => \N__40925\,
            in2 => \N__41143\,
            in3 => \N__41068\,
            lcout => n14690,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9490_2_lut_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55447\,
            lcout => n11202,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12268_2_lut_4_lut_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000100"
        )
    port map (
            in0 => \N__56276\,
            in1 => \N__40893\,
            in2 => \N__41142\,
            in3 => \N__41067\,
            lcout => n14688,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i12_1_lut_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46197\,
            lcout => n14_adj_580,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_76_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41084\,
            in1 => \N__40892\,
            in2 => \N__40927\,
            in3 => \N__40820\,
            lcout => OPEN,
            ltout => \n14_adj_679_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40664\,
            in1 => \N__40718\,
            in2 => \N__40741\,
            in3 => \N__43507\,
            lcout => n4781,
            ltout => \n4781_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9491_1_lut_2_lut_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40738\,
            in3 => \N__55507\,
            lcout => n1259,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i0_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__40735\,
            in1 => \N__40729\,
            in2 => \N__40723\,
            in3 => \N__40702\,
            lcout => dti_counter_0,
            ltout => OPEN,
            carryin => \bfn_12_27_0_\,
            carryout => n12742,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i1_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__40699\,
            in1 => \N__40855\,
            in2 => \N__43528\,
            in3 => \N__40693\,
            lcout => dti_counter_1,
            ltout => OPEN,
            carryin => n12742,
            carryout => n12743,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i2_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__40690\,
            in1 => \N__43545\,
            in2 => \N__40868\,
            in3 => \N__40684\,
            lcout => dti_counter_2,
            ltout => OPEN,
            carryin => n12743,
            carryout => n12744,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i3_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__40681\,
            in1 => \N__40859\,
            in2 => \N__40674\,
            in3 => \N__40648\,
            lcout => dti_counter_3,
            ltout => OPEN,
            carryin => n12744,
            carryout => n12745,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i4_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__40936\,
            in1 => \N__40926\,
            in2 => \N__40869\,
            in3 => \N__40906\,
            lcout => dti_counter_4,
            ltout => OPEN,
            carryin => n12745,
            carryout => n12746,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i5_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__41026\,
            in1 => \N__40863\,
            in2 => \N__41094\,
            in3 => \N__40903\,
            lcout => dti_counter_5,
            ltout => OPEN,
            carryin => n12746,
            carryout => n12747,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i6_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__40900\,
            in1 => \N__40894\,
            in2 => \N__40870\,
            in3 => \N__40879\,
            lcout => dti_counter_6,
            ltout => OPEN,
            carryin => n12747,
            carryout => n12748,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_633__i7_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__40876\,
            in1 => \N__40867\,
            in2 => \N__40830\,
            in3 => \N__40834\,
            lcout => dti_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i4_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55711\,
            in1 => \N__43714\,
            in2 => \_gnd_net_\,
            in3 => \N__46003\,
            lcout => pwm_setpoint_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12273_3_lut_4_lut_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__41019\,
            in1 => \N__40749\,
            in2 => \N__40786\,
            in3 => \N__40766\,
            lcout => n14745,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i6_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55712\,
            in1 => \N__43681\,
            in2 => \_gnd_net_\,
            in3 => \N__46321\,
            lcout => pwm_setpoint_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i3_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43735\,
            in1 => \N__50197\,
            in2 => \_gnd_net_\,
            in3 => \N__55713\,
            lcout => pwm_setpoint_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i6_3_lut_3_lut_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101010000"
        )
    port map (
            in0 => \N__40767\,
            in1 => \_gnd_net_\,
            in2 => \N__40753\,
            in3 => \N__41020\,
            lcout => n6_adj_606,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12279_2_lut_4_lut_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__56275\,
            in1 => \N__41139\,
            in2 => \N__41095\,
            in3 => \N__41060\,
            lcout => n14689,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i2_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55710\,
            in1 => \N__43744\,
            in2 => \_gnd_net_\,
            in3 => \N__46048\,
            lcout => pwm_setpoint_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i5_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55698\,
            in1 => \N__43699\,
            in2 => \_gnd_net_\,
            in3 => \N__45961\,
            lcout => pwm_setpoint_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i11_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__46198\,
            in1 => \N__55700\,
            in2 => \_gnd_net_\,
            in3 => \N__43798\,
            lcout => pwm_setpoint_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i12_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__55697\,
            in1 => \_gnd_net_\,
            in2 => \N__43789\,
            in3 => \N__46795\,
            lcout => pwm_setpoint_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i8_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52732\,
            in1 => \N__43837\,
            in2 => \_gnd_net_\,
            in3 => \N__55701\,
            lcout => pwm_setpoint_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i8_1_lut_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46948\,
            lcout => n18_adj_584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i21_2_lut_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41292\,
            in2 => \_gnd_net_\,
            in3 => \N__40973\,
            lcout => n21_adj_617,
            ltout => \n21_adj_617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12370_3_lut_LC_12_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41293\,
            in1 => \_gnd_net_\,
            in2 => \N__40957\,
            in3 => \N__40954\,
            lcout => n14842,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i10_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43816\,
            in1 => \N__55699\,
            in2 => \_gnd_net_\,
            in3 => \N__46234\,
            lcout => pwm_setpoint_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i11_2_lut_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41280\,
            in2 => \_gnd_net_\,
            in3 => \N__41186\,
            lcout => n11_adj_610,
            ltout => \n11_adj_610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12256_4_lut_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__41235\,
            in1 => \N__41304\,
            in2 => \N__41284\,
            in3 => \N__46713\,
            lcout => n14728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i19_LC_12_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__50281\,
            in1 => \N__55702\,
            in2 => \_gnd_net_\,
            in3 => \N__43906\,
            lcout => pwm_setpoint_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56078\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i10_3_lut_3_lut_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__41281\,
            in1 => \N__41271\,
            in2 => \_gnd_net_\,
            in3 => \N__41165\,
            lcout => n10_adj_609,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_67_LC_12_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41476\,
            in2 => \_gnd_net_\,
            in3 => \N__41500\,
            lcout => n4825,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12332_4_lut_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__41778\,
            in1 => \N__41236\,
            in2 => \N__41221\,
            in3 => \N__41212\,
            lcout => n14804,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i20_LC_12_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__47065\,
            in1 => \_gnd_net_\,
            in2 => \N__55714\,
            in3 => \N__43897\,
            lcout => pwm_setpoint_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56078\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i2_3_lut_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__41191\,
            in1 => \N__41170\,
            in2 => \_gnd_net_\,
            in3 => \N__47031\,
            lcout => OPEN,
            ltout => \PWM.n13596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i1_4_lut_LC_12_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__41400\,
            in1 => \N__41342\,
            in2 => \N__41536\,
            in3 => \N__41532\,
            lcout => OPEN,
            ltout => \PWM.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i13_4_lut_LC_12_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41512\,
            in1 => \N__41496\,
            in2 => \N__41479\,
            in3 => \N__41711\,
            lcout => OPEN,
            ltout => \PWM.n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i9623_4_lut_LC_12_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__41474\,
            in1 => \N__44041\,
            in2 => \N__41455\,
            in3 => \N__41452\,
            lcout => \PWM.pwm_counter_31__N_401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i15_2_lut_LC_12_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47030\,
            in2 => \_gnd_net_\,
            in3 => \N__46927\,
            lcout => n15_adj_613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i39_2_lut_LC_12_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41373\,
            in2 => \_gnd_net_\,
            in3 => \N__41399\,
            lcout => n39,
            ltout => \n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12411_3_lut_LC_12_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41374\,
            in1 => \_gnd_net_\,
            in2 => \N__41365\,
            in3 => \N__43963\,
            lcout => n14883,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i19_2_lut_LC_12_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52763\,
            in2 => \_gnd_net_\,
            in3 => \N__41343\,
            lcout => n19_adj_616,
            ltout => \n19_adj_616_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12328_4_lut_LC_12_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__41317\,
            in1 => \N__41799\,
            in2 => \N__41308\,
            in3 => \N__41305\,
            lcout => OPEN,
            ltout => \n14800_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12398_4_lut_LC_12_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41763\,
            in1 => \N__41832\,
            in2 => \N__41809\,
            in3 => \N__41685\,
            lcout => n14870,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12262_4_lut_LC_12_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__41806\,
            in1 => \N__41800\,
            in2 => \N__41785\,
            in3 => \N__41764\,
            lcout => n14734,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12402_4_lut_LC_12_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43981\,
            in1 => \N__43924\,
            in2 => \N__46891\,
            in3 => \N__46804\,
            lcout => n14874,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i25_2_lut_LC_12_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41713\,
            lcout => n25_adj_620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12347_3_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41674\,
            in2 => \N__41650\,
            in3 => \N__47568\,
            lcout => n2822,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1856_3_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41637\,
            in1 => \_gnd_net_\,
            in2 => \N__47605\,
            in3 => \N__41617\,
            lcout => n2824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_55_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44165\,
            in1 => \N__41611\,
            in2 => \N__44116\,
            in3 => \N__41602\,
            lcout => OPEN,
            ltout => \n14054_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_56_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42231\,
            in1 => \N__41593\,
            in2 => \N__41575\,
            in3 => \N__44246\,
            lcout => OPEN,
            ltout => \n14060_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13000_4_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42305\,
            in1 => \N__41568\,
            in2 => \N__41539\,
            in3 => \N__42027\,
            lcout => n2742,
            ltout => \n2742_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1862_3_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41998\,
            in2 => \N__41992\,
            in3 => \N__41989\,
            lcout => n2830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1859_3_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41961\,
            in2 => \N__41938\,
            in3 => \N__47567\,
            lcout => n2827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_44_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47762\,
            in1 => \N__48128\,
            in2 => \N__48224\,
            in3 => \N__47726\,
            lcout => OPEN,
            ltout => \n14238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_45_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48176\,
            in2 => \N__41929\,
            in3 => \N__48303\,
            lcout => OPEN,
            ltout => \n14240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_46_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48038\,
            in1 => \N__47999\,
            in2 => \N__41926\,
            in3 => \N__48080\,
            lcout => n14246,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1851_3_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__47577\,
            in1 => \_gnd_net_\,
            in2 => \N__41923\,
            in3 => \N__41905\,
            lcout => n2819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1853_3_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41896\,
            in1 => \_gnd_net_\,
            in2 => \N__41890\,
            in3 => \N__47572\,
            lcout => n2821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1861_3_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41863\,
            in2 => \N__47606\,
            in3 => \N__41857\,
            lcout => n2829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12349_3_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42183\,
            in2 => \N__42160\,
            in3 => \N__47573\,
            lcout => n2823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1850_3_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42148\,
            in2 => \N__47607\,
            in3 => \N__42142\,
            lcout => n2818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1921_3_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__48186\,
            in1 => \_gnd_net_\,
            in2 => \N__48160\,
            in3 => \N__49312\,
            lcout => n2921,
            ltout => \n2921_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_36_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42100\,
            in3 => \N__44528\,
            lcout => n13926,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1915_3_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48553\,
            in2 => \N__48523\,
            in3 => \N__49316\,
            lcout => n2915,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1918_3_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48042\,
            in2 => \N__49353\,
            in3 => \N__48022\,
            lcout => n2918,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1842_3_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42097\,
            in2 => \N__42310\,
            in3 => \N__47594\,
            lcout => n2810,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1917_3_lut_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48604\,
            in2 => \N__49354\,
            in3 => \N__48003\,
            lcout => n2917,
            ltout => \n2917_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_38_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42053\,
            in1 => \N__42037\,
            in2 => \N__42031\,
            in3 => \N__44456\,
            lcout => OPEN,
            ltout => \n13934_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_39_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42548\,
            in1 => \N__42524\,
            in2 => \N__42508\,
            in3 => \N__44704\,
            lcout => n13942,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1775_3_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42496\,
            in2 => \N__42484\,
            in3 => \N__42444\,
            lcout => n2711,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12995_1_lut_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47625\,
            in3 => \_gnd_net_\,
            lcout => n15467,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1909_3_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49336\,
            in2 => \N__48906\,
            in3 => \N__48880\,
            lcout => n2909,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2119_3_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51730\,
            in2 => \N__50118\,
            in3 => \N__51749\,
            lcout => n3215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2122_3_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51222\,
            in2 => \N__51199\,
            in3 => \N__50109\,
            lcout => n3218,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1844_3_lut_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42232\,
            in2 => \N__47626\,
            in3 => \N__42202\,
            lcout => n2812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_29_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45491\,
            in1 => \N__45146\,
            in2 => \N__45456\,
            in3 => \N__45113\,
            lcout => OPEN,
            ltout => \n14322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_30_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45423\,
            in1 => \N__45378\,
            in2 => \N__42196\,
            in3 => \N__42637\,
            lcout => n14328,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1992_3_lut_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42664\,
            in1 => \N__44943\,
            in2 => \_gnd_net_\,
            in3 => \N__42946\,
            lcout => n3024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1991_3_lut_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44460\,
            in1 => \_gnd_net_\,
            in2 => \N__42994\,
            in3 => \N__42652\,
            lcout => n3023,
            ltout => \n3023_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_28_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45044\,
            in1 => \N__45008\,
            in2 => \N__42640\,
            in3 => \N__45083\,
            lcout => n14320,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1995_3_lut_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42631\,
            in2 => \N__42995\,
            in3 => \N__44571\,
            lcout => n3027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1994_3_lut_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44625\,
            in2 => \N__42622\,
            in3 => \N__42945\,
            lcout => n3026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1913_3_lut_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48442\,
            in2 => \N__48469\,
            in3 => \N__49359\,
            lcout => n2913,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2061_3_lut_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45067\,
            in2 => \N__49041\,
            in3 => \N__45087\,
            lcout => n3125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1990_3_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42583\,
            in2 => \N__44308\,
            in3 => \N__42961\,
            lcout => n3022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1982_3_lut_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__42963\,
            in1 => \_gnd_net_\,
            in2 => \N__42574\,
            in3 => \N__42558\,
            lcout => n3014,
            ltout => \n3014_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__45345\,
            in1 => \_gnd_net_\,
            in2 => \N__43018\,
            in3 => \N__45269\,
            lcout => n14408,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1989_3_lut_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__42962\,
            in1 => \N__42862\,
            in2 => \N__44544\,
            in3 => \_gnd_net_\,
            lcout => n3021,
            ltout => \n3021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2056_3_lut_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45439\,
            in2 => \N__42853\,
            in3 => \N__48988\,
            lcout => n3120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2066_3_lut_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44716\,
            in2 => \N__49042\,
            in3 => \N__44742\,
            lcout => n3130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_2_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42850\,
            in2 => \N__54865\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => n12521,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_3_lut_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42823\,
            in2 => \_gnd_net_\,
            in3 => \N__42772\,
            lcout => n3301,
            ltout => OPEN,
            carryin => n12521,
            carryout => n12522,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_4_lut_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42769\,
            in2 => \N__54866\,
            in3 => \N__42730\,
            lcout => n3300,
            ltout => OPEN,
            carryin => n12522,
            carryout => n12523,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_5_lut_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42723\,
            in2 => \_gnd_net_\,
            in3 => \N__42694\,
            lcout => n3299,
            ltout => OPEN,
            carryin => n12523,
            carryout => n12524,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_6_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42691\,
            in2 => \N__54867\,
            in3 => \N__42667\,
            lcout => n3298,
            ltout => OPEN,
            carryin => n12524,
            carryout => n12525,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_7_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__43111\,
            in1 => \_gnd_net_\,
            in2 => \N__43105\,
            in3 => \N__43066\,
            lcout => n14697,
            ltout => OPEN,
            carryin => n12525,
            carryout => n12526,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_8_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48682\,
            in2 => \_gnd_net_\,
            in3 => \N__43063\,
            lcout => n3296,
            ltout => OPEN,
            carryin => n12526,
            carryout => n12527,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_9_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54403\,
            in2 => \N__45787\,
            in3 => \N__43060\,
            lcout => n3295,
            ltout => OPEN,
            carryin => n12527,
            carryout => n12528,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_10_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46107\,
            in2 => \N__54868\,
            in3 => \N__43057\,
            lcout => n3294,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => n12529,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_11_lut_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49398\,
            in2 => \N__54872\,
            in3 => \N__43048\,
            lcout => n3293,
            ltout => OPEN,
            carryin => n12529,
            carryout => n12530,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_12_lut_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49656\,
            in2 => \N__54869\,
            in3 => \N__43045\,
            lcout => n3292,
            ltout => OPEN,
            carryin => n12530,
            carryout => n12531,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_13_lut_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45765\,
            in2 => \N__54873\,
            in3 => \N__43033\,
            lcout => n3291,
            ltout => OPEN,
            carryin => n12531,
            carryout => n12532,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_14_lut_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46133\,
            in2 => \N__54870\,
            in3 => \N__43021\,
            lcout => n3290,
            ltout => OPEN,
            carryin => n12532,
            carryout => n12533,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_15_lut_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48635\,
            in2 => \N__54874\,
            in3 => \N__43267\,
            lcout => n3289,
            ltout => OPEN,
            carryin => n12533,
            carryout => n12534,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_16_lut_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45870\,
            in2 => \N__54871\,
            in3 => \N__43258\,
            lcout => n3288,
            ltout => OPEN,
            carryin => n12534,
            carryout => n12535,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_17_lut_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48734\,
            in2 => \N__54875\,
            in3 => \N__43255\,
            lcout => n3287,
            ltout => OPEN,
            carryin => n12535,
            carryout => n12536,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_18_lut_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49689\,
            in2 => \N__54876\,
            in3 => \N__43252\,
            lcout => n3286,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => n12537,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_19_lut_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54431\,
            in2 => \N__45838\,
            in3 => \N__43243\,
            lcout => n3285,
            ltout => OPEN,
            carryin => n12537,
            carryout => n12538,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_20_lut_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43236\,
            in2 => \N__54877\,
            in3 => \N__43210\,
            lcout => n3284,
            ltout => OPEN,
            carryin => n12538,
            carryout => n12539,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_21_lut_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43207\,
            in2 => \N__54880\,
            in3 => \N__43174\,
            lcout => n3283,
            ltout => OPEN,
            carryin => n12539,
            carryout => n12540,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_22_lut_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43166\,
            in2 => \N__54878\,
            in3 => \N__43135\,
            lcout => n3282,
            ltout => OPEN,
            carryin => n12540,
            carryout => n12541,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_23_lut_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43130\,
            in2 => \N__54881\,
            in3 => \N__43495\,
            lcout => n3281,
            ltout => OPEN,
            carryin => n12541,
            carryout => n12542,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_24_lut_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49928\,
            in2 => \N__54879\,
            in3 => \N__43486\,
            lcout => n3280,
            ltout => OPEN,
            carryin => n12542,
            carryout => n12543,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_25_lut_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43483\,
            in2 => \N__54882\,
            in3 => \N__43444\,
            lcout => n3279,
            ltout => OPEN,
            carryin => n12543,
            carryout => n12544,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_26_lut_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43440\,
            in2 => \N__54883\,
            in3 => \N__43405\,
            lcout => n3278,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => n12545,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_27_lut_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43402\,
            in2 => \N__54887\,
            in3 => \N__43363\,
            lcout => n3277,
            ltout => OPEN,
            carryin => n12545,
            carryout => n12546,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_28_lut_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49427\,
            in2 => \N__54884\,
            in3 => \N__43348\,
            lcout => n3276,
            ltout => OPEN,
            carryin => n12546,
            carryout => n12547,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_29_lut_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43345\,
            in2 => \N__54888\,
            in3 => \N__43309\,
            lcout => n3275,
            ltout => OPEN,
            carryin => n12547,
            carryout => n12548,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_30_lut_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43306\,
            in2 => \N__54885\,
            in3 => \N__43270\,
            lcout => n3274,
            ltout => OPEN,
            carryin => n12548,
            carryout => n12549,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_31_lut_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43672\,
            in2 => \N__54889\,
            in3 => \N__43630\,
            lcout => n3273,
            ltout => OPEN,
            carryin => n12549,
            carryout => n12550,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_32_lut_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43627\,
            in2 => \N__54886\,
            in3 => \N__43594\,
            lcout => n3272,
            ltout => OPEN,
            carryin => n12550,
            carryout => n12551,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_33_lut_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54471\,
            in1 => \N__43591\,
            in2 => \N__51910\,
            in3 => \N__43573\,
            lcout => n14461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i7_1_lut_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46314\,
            lcout => n19_adj_585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i3_1_lut_LC_13_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46041\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n23_adj_589,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i11_1_lut_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46227\,
            lcout => n15_adj_581,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i6_1_lut_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45954\,
            lcout => n20_adj_586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i4_1_lut_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43558\,
            lcout => n22_adj_548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43544\,
            in2 => \_gnd_net_\,
            in3 => \N__43523\,
            lcout => n10_adj_680,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i1_1_lut_LC_13_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46473\,
            lcout => n25_adj_591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i15_1_lut_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46560\,
            lcout => n11_adj_577,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_2_lut_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43762\,
            in2 => \_gnd_net_\,
            in3 => \N__43756\,
            lcout => \pwm_setpoint_23_N_171_0\,
            ltout => OPEN,
            carryin => \bfn_13_28_0_\,
            carryout => n12050,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_3_lut_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50206\,
            in2 => \_gnd_net_\,
            in3 => \N__43753\,
            lcout => \pwm_setpoint_23_N_171_1\,
            ltout => OPEN,
            carryin => n12050,
            carryout => n12051,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_4_lut_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43750\,
            in2 => \_gnd_net_\,
            in3 => \N__43738\,
            lcout => \pwm_setpoint_23_N_171_2\,
            ltout => OPEN,
            carryin => n12051,
            carryout => n12052,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_5_lut_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50173\,
            in2 => \_gnd_net_\,
            in3 => \N__43729\,
            lcout => \pwm_setpoint_23_N_171_3\,
            ltout => OPEN,
            carryin => n12052,
            carryout => n12053,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_6_lut_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43726\,
            in2 => \_gnd_net_\,
            in3 => \N__43708\,
            lcout => \pwm_setpoint_23_N_171_4\,
            ltout => OPEN,
            carryin => n12053,
            carryout => n12054,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_7_lut_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43705\,
            in2 => \_gnd_net_\,
            in3 => \N__43690\,
            lcout => \pwm_setpoint_23_N_171_5\,
            ltout => OPEN,
            carryin => n12054,
            carryout => n12055,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_8_lut_LC_13_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43687\,
            in2 => \_gnd_net_\,
            in3 => \N__43675\,
            lcout => \pwm_setpoint_23_N_171_6\,
            ltout => OPEN,
            carryin => n12055,
            carryout => n12056,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_9_lut_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43846\,
            in2 => \_gnd_net_\,
            in3 => \N__43840\,
            lcout => \pwm_setpoint_23_N_171_7\,
            ltout => OPEN,
            carryin => n12056,
            carryout => n12057,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_10_lut_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52711\,
            in2 => \_gnd_net_\,
            in3 => \N__43831\,
            lcout => \pwm_setpoint_23_N_171_8\,
            ltout => OPEN,
            carryin => \bfn_13_29_0_\,
            carryout => n12058,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_11_lut_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46510\,
            in2 => \_gnd_net_\,
            in3 => \N__43828\,
            lcout => \pwm_setpoint_23_N_171_9\,
            ltout => OPEN,
            carryin => n12058,
            carryout => n12059,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_12_lut_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43825\,
            in2 => \_gnd_net_\,
            in3 => \N__43810\,
            lcout => \pwm_setpoint_23_N_171_10\,
            ltout => OPEN,
            carryin => n12059,
            carryout => n12060,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_13_lut_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43807\,
            in2 => \_gnd_net_\,
            in3 => \N__43792\,
            lcout => \pwm_setpoint_23_N_171_11\,
            ltout => OPEN,
            carryin => n12060,
            carryout => n12061,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_14_lut_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46774\,
            in2 => \_gnd_net_\,
            in3 => \N__43780\,
            lcout => \pwm_setpoint_23_N_171_12\,
            ltout => OPEN,
            carryin => n12061,
            carryout => n12062,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_15_lut_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46489\,
            in2 => \_gnd_net_\,
            in3 => \N__43777\,
            lcout => \pwm_setpoint_23_N_171_13\,
            ltout => OPEN,
            carryin => n12062,
            carryout => n12063,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_16_lut_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43774\,
            in2 => \_gnd_net_\,
            in3 => \N__43765\,
            lcout => \pwm_setpoint_23_N_171_14\,
            ltout => OPEN,
            carryin => n12063,
            carryout => n12064,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_17_lut_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46570\,
            in2 => \_gnd_net_\,
            in3 => \N__43918\,
            lcout => \pwm_setpoint_23_N_171_15\,
            ltout => OPEN,
            carryin => n12064,
            carryout => n12065,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_18_lut_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46645\,
            in2 => \_gnd_net_\,
            in3 => \N__43915\,
            lcout => \pwm_setpoint_23_N_171_16\,
            ltout => OPEN,
            carryin => \bfn_13_30_0_\,
            carryout => n12066,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_19_lut_LC_13_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47134\,
            in2 => \_gnd_net_\,
            in3 => \N__43912\,
            lcout => \pwm_setpoint_23_N_171_17\,
            ltout => OPEN,
            carryin => n12066,
            carryout => n12067,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_20_lut_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50233\,
            in2 => \_gnd_net_\,
            in3 => \N__43909\,
            lcout => \pwm_setpoint_23_N_171_18\,
            ltout => OPEN,
            carryin => n12067,
            carryout => n12068,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_21_lut_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50260\,
            in2 => \_gnd_net_\,
            in3 => \N__43900\,
            lcout => \pwm_setpoint_23_N_171_19\,
            ltout => OPEN,
            carryin => n12068,
            carryout => n12069,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_22_lut_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47044\,
            in2 => \_gnd_net_\,
            in3 => \N__43891\,
            lcout => \pwm_setpoint_23_N_171_20\,
            ltout => OPEN,
            carryin => n12069,
            carryout => n12070,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_23_lut_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43888\,
            in2 => \_gnd_net_\,
            in3 => \N__43864\,
            lcout => \pwm_setpoint_23_N_171_21\,
            ltout => OPEN,
            carryin => n12070,
            carryout => n12071,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_24_lut_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46651\,
            in2 => \_gnd_net_\,
            in3 => \N__43861\,
            lcout => \pwm_setpoint_23_N_171_22\,
            ltout => OPEN,
            carryin => n12071,
            carryout => n12072,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i23_LC_13_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55563\,
            in2 => \_gnd_net_\,
            in3 => \N__43858\,
            lcout => pwm_setpoint_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56082\,
            ce => 'H',
            sr => \N__55567\
        );

    \pwm_setpoint_i15_LC_13_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44077\,
            in1 => \N__55656\,
            in2 => \_gnd_net_\,
            in3 => \N__46588\,
            lcout => pwm_setpoint_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i18_LC_13_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55655\,
            in1 => \N__50251\,
            in2 => \_gnd_net_\,
            in3 => \N__44068\,
            lcout => pwm_setpoint_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i12_4_lut_LC_13_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44061\,
            in1 => \N__44274\,
            in2 => \N__46843\,
            in3 => \N__46747\,
            lcout => \PWM.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i31_2_lut_LC_13_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46980\,
            in2 => \_gnd_net_\,
            in3 => \N__44031\,
            lcout => n31_adj_624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i37_2_lut_LC_13_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43974\,
            in2 => \_gnd_net_\,
            in3 => \N__44000\,
            lcout => n37,
            ltout => \n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12415_3_lut_LC_13_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__43975\,
            in1 => \_gnd_net_\,
            in2 => \N__43966\,
            in3 => \N__46987\,
            lcout => n14887,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i22_LC_13_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55709\,
            in1 => \N__46666\,
            in2 => \_gnd_net_\,
            in3 => \N__43957\,
            lcout => pwm_setpoint_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i17_LC_13_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47152\,
            in1 => \N__55708\,
            in2 => \_gnd_net_\,
            in3 => \N__43939\,
            lcout => pwm_setpoint_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56090\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12360_4_lut_LC_13_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__43930\,
            in1 => \N__47179\,
            in2 => \N__46720\,
            in3 => \N__47212\,
            lcout => n14832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i35_2_lut_LC_13_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46905\,
            in2 => \_gnd_net_\,
            in3 => \N__44275\,
            lcout => n35,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1843_3_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44251\,
            in2 => \N__44224\,
            in3 => \N__47562\,
            lcout => n2811,
            ltout => \n2811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_48_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48384\,
            in1 => \N__44083\,
            in2 => \N__44209\,
            in3 => \N__48425\,
            lcout => n14266,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1858_3_lut_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44206\,
            in2 => \N__44197\,
            in3 => \N__47554\,
            lcout => n2826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1933_3_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47227\,
            in1 => \N__47260\,
            in2 => \_gnd_net_\,
            in3 => \N__49273\,
            lcout => n2933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1847_3_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44166\,
            in2 => \N__44143\,
            in3 => \N__47558\,
            lcout => n2815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1846_3_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44128\,
            in2 => \N__47603\,
            in3 => \N__44115\,
            lcout => n2814,
            ltout => \n2814_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_43_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47810\,
            in1 => \N__48263\,
            in2 => \N__44086\,
            in3 => \N__48494\,
            lcout => n14260,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1860_3_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__44440\,
            in1 => \_gnd_net_\,
            in2 => \N__47602\,
            in3 => \N__44431\,
            lcout => n2828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1864_3_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44404\,
            in2 => \N__44392\,
            in3 => \N__47563\,
            lcout => n2832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1863_3_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44362\,
            in2 => \N__47604\,
            in3 => \N__44350\,
            lcout => n2831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1929_3_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__47866\,
            in1 => \_gnd_net_\,
            in2 => \N__47889\,
            in3 => \N__49320\,
            lcout => n2929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_47_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__47470\,
            in1 => \N__47882\,
            in2 => \N__47850\,
            in3 => \N__44329\,
            lcout => OPEN,
            ltout => \n14248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_49_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48545\,
            in1 => \N__48585\,
            in2 => \N__44323\,
            in3 => \N__48864\,
            lcout => OPEN,
            ltout => \n14254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12452_4_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48800\,
            in1 => \N__48896\,
            in2 => \N__44320\,
            in3 => \N__44317\,
            lcout => n2841,
            ltout => \n2841_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1923_3_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__48247\,
            in1 => \_gnd_net_\,
            in2 => \N__44311\,
            in3 => \N__48273\,
            lcout => n2923,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_35_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44556\,
            in1 => \N__44286\,
            in2 => \N__44654\,
            in3 => \N__44939\,
            lcout => OPEN,
            ltout => \n13932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_37_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44615\,
            in1 => \N__44684\,
            in2 => \N__44707\,
            in3 => \N__44588\,
            lcout => n13936,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1926_3_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47746\,
            in2 => \N__47782\,
            in3 => \N__49296\,
            lcout => n2926,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1920_3_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49293\,
            in1 => \_gnd_net_\,
            in2 => \N__48138\,
            in3 => \N__48112\,
            lcout => n2920,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1927_3_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47814\,
            in1 => \N__47791\,
            in2 => \_gnd_net_\,
            in3 => \N__49295\,
            lcout => n2927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1919_3_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__49297\,
            in1 => \N__48061\,
            in2 => \N__48100\,
            in3 => \_gnd_net_\,
            lcout => n2919,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1928_3_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47824\,
            in1 => \N__47846\,
            in2 => \_gnd_net_\,
            in3 => \N__49292\,
            lcout => n2928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1922_3_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49294\,
            in1 => \_gnd_net_\,
            in2 => \N__48234\,
            in3 => \N__48202\,
            lcout => n2922,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12351_3_lut_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44515\,
            in2 => \N__44503\,
            in3 => \N__47595\,
            lcout => n2825,
            ltout => \n2825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1924_3_lut_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49326\,
            in1 => \_gnd_net_\,
            in2 => \N__44470\,
            in3 => \N__48286\,
            lcout => n2924,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1925_3_lut_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47736\,
            in2 => \N__47707\,
            in3 => \N__49325\,
            lcout => n2925,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2058_3_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44979\,
            in2 => \N__44965\,
            in3 => \N__49065\,
            lcout => n3122,
            ltout => \n3122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2125_3_lut_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__51325\,
            in1 => \_gnd_net_\,
            in2 => \N__44923\,
            in3 => \N__50108\,
            lcout => n3221,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1914_3_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48504\,
            in2 => \N__49358\,
            in3 => \N__48481\,
            lcout => n2914,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2062_3_lut_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__45097\,
            in1 => \_gnd_net_\,
            in2 => \N__49083\,
            in3 => \N__45117\,
            lcout => n3126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_2_lut_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44893\,
            in2 => \_gnd_net_\,
            in3 => \N__44839\,
            lcout => n3101,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => n12464,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_3_lut_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55190\,
            in2 => \N__44836\,
            in3 => \N__44791\,
            lcout => n3100,
            ltout => OPEN,
            carryin => n12464,
            carryout => n12465,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_4_lut_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44787\,
            in2 => \_gnd_net_\,
            in3 => \N__44746\,
            lcout => n3099,
            ltout => OPEN,
            carryin => n12465,
            carryout => n12466,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_5_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55191\,
            in2 => \N__44743\,
            in3 => \N__44710\,
            lcout => n3098,
            ltout => OPEN,
            carryin => n12466,
            carryout => n12467,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_6_lut_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45229\,
            in3 => \N__45190\,
            lcout => n3097,
            ltout => OPEN,
            carryin => n12467,
            carryout => n12468,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_7_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45187\,
            in2 => \_gnd_net_\,
            in3 => \N__45157\,
            lcout => n3096,
            ltout => OPEN,
            carryin => n12468,
            carryout => n12469,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_8_lut_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55060\,
            in2 => \N__45154\,
            in3 => \N__45121\,
            lcout => n3095,
            ltout => OPEN,
            carryin => n12469,
            carryout => n12470,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_9_lut_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55192\,
            in2 => \N__45118\,
            in3 => \N__45091\,
            lcout => n3094,
            ltout => OPEN,
            carryin => n12470,
            carryout => n12471,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_10_lut_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54618\,
            in2 => \N__45088\,
            in3 => \N__45061\,
            lcout => n3093,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => n12472,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_11_lut_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54340\,
            in2 => \N__45058\,
            in3 => \N__45016\,
            lcout => n3092,
            ltout => OPEN,
            carryin => n12472,
            carryout => n12473,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_12_lut_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54619\,
            in2 => \N__45013\,
            in3 => \N__44983\,
            lcout => n3091,
            ltout => OPEN,
            carryin => n12473,
            carryout => n12474,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_13_lut_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54341\,
            in2 => \N__44980\,
            in3 => \N__44953\,
            lcout => n3090,
            ltout => OPEN,
            carryin => n12474,
            carryout => n12475,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_14_lut_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54620\,
            in2 => \N__45496\,
            in3 => \N__45460\,
            lcout => n3089,
            ltout => OPEN,
            carryin => n12475,
            carryout => n12476,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_15_lut_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54342\,
            in2 => \N__45457\,
            in3 => \N__45433\,
            lcout => n3088,
            ltout => OPEN,
            carryin => n12476,
            carryout => n12477,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_16_lut_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54621\,
            in2 => \N__45430\,
            in3 => \N__45385\,
            lcout => n3087,
            ltout => OPEN,
            carryin => n12477,
            carryout => n12478,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_17_lut_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45382\,
            in2 => \N__54979\,
            in3 => \N__45352\,
            lcout => n3086,
            ltout => OPEN,
            carryin => n12478,
            carryout => n12479,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_18_lut_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54649\,
            in2 => \N__45349\,
            in3 => \N__45310\,
            lcout => n3085,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => n12480,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_19_lut_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45307\,
            in2 => \N__54988\,
            in3 => \N__45277\,
            lcout => n3084,
            ltout => OPEN,
            carryin => n12480,
            carryout => n12481,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_20_lut_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45274\,
            in2 => \N__55247\,
            in3 => \N__45235\,
            lcout => n3083,
            ltout => OPEN,
            carryin => n12481,
            carryout => n12482,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_21_lut_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49125\,
            in2 => \N__54989\,
            in3 => \N__45232\,
            lcout => n3082,
            ltout => OPEN,
            carryin => n12482,
            carryout => n12483,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_22_lut_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45732\,
            in2 => \N__55248\,
            in3 => \N__45712\,
            lcout => n3081,
            ltout => OPEN,
            carryin => n12483,
            carryout => n12484,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_23_lut_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45709\,
            in2 => \N__54990\,
            in3 => \N__45673\,
            lcout => n3080,
            ltout => OPEN,
            carryin => n12484,
            carryout => n12485,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_24_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45669\,
            in2 => \N__55249\,
            in3 => \N__45637\,
            lcout => n3079,
            ltout => OPEN,
            carryin => n12485,
            carryout => n12486,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_25_lut_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49470\,
            in2 => \N__54991\,
            in3 => \N__45634\,
            lcout => n3078,
            ltout => OPEN,
            carryin => n12486,
            carryout => n12487,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_26_lut_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54669\,
            in2 => \N__45631\,
            in3 => \N__45595\,
            lcout => n3077,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => n12488,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_27_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49185\,
            in2 => \N__54994\,
            in3 => \N__45592\,
            lcout => n3076,
            ltout => OPEN,
            carryin => n12488,
            carryout => n12489,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_28_lut_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45589\,
            in2 => \N__54978\,
            in3 => \N__45547\,
            lcout => n3075,
            ltout => OPEN,
            carryin => n12489,
            carryout => n12490,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_29_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45544\,
            in2 => \N__54995\,
            in3 => \N__45499\,
            lcout => n3074,
            ltout => OPEN,
            carryin => n12490,
            carryout => n12491,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_30_lut_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54609\,
            in1 => \N__45939\,
            in2 => \N__45916\,
            in3 => \N__45889\,
            lcout => n3105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2128_3_lut_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51497\,
            in2 => \N__51466\,
            in3 => \N__50068\,
            lcout => n3224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2199_3_lut_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45886\,
            in2 => \N__49612\,
            in3 => \N__45783\,
            lcout => n15_adj_704,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2198_3_lut_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46108\,
            in2 => \N__45880\,
            in3 => \N__49589\,
            lcout => n17_adj_705,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_152_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49655\,
            in1 => \N__46106\,
            in2 => \N__45745\,
            in3 => \N__45863\,
            lcout => OPEN,
            ltout => \n14368_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_153_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45833\,
            in1 => \N__49688\,
            in2 => \N__45805\,
            in3 => \N__46114\,
            lcout => n14374,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2132_3_lut_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50929\,
            in2 => \N__50896\,
            in3 => \N__50113\,
            lcout => n3228,
            ltout => \n3228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_150_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45769\,
            in3 => \N__45758\,
            lcout => n14362,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_151_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49386\,
            in1 => \N__48741\,
            in2 => \N__46141\,
            in3 => \N__48639\,
            lcout => n14366,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2131_3_lut_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__50877\,
            in1 => \N__50839\,
            in2 => \N__50119\,
            in3 => \_gnd_net_\,
            lcout => n3227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2123_3_lut_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51272\,
            in2 => \N__51241\,
            in3 => \N__50117\,
            lcout => n3219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i0_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51880\,
            in2 => \N__46090\,
            in3 => \N__46078\,
            lcout => duty_0,
            ltout => OPEN,
            carryin => \bfn_14_26_0_\,
            carryout => n12073,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i1_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52474\,
            in2 => \N__46075\,
            in3 => \N__46063\,
            lcout => duty_1,
            ltout => OPEN,
            carryin => n12073,
            carryout => n12074,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i2_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46060\,
            in2 => \N__52447\,
            in3 => \N__46030\,
            lcout => duty_2,
            ltout => OPEN,
            carryin => n12074,
            carryout => n12075,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i3_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52414\,
            in2 => \N__46027\,
            in3 => \N__46018\,
            lcout => duty_3,
            ltout => OPEN,
            carryin => n12075,
            carryout => n12076,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i4_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52387\,
            in2 => \N__46015\,
            in3 => \N__45979\,
            lcout => duty_4,
            ltout => OPEN,
            carryin => n12076,
            carryout => n12077,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i5_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52357\,
            in2 => \N__45976\,
            in3 => \N__45943\,
            lcout => duty_5,
            ltout => OPEN,
            carryin => n12077,
            carryout => n12078,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i6_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52332\,
            in2 => \N__55531\,
            in3 => \N__46303\,
            lcout => duty_6,
            ltout => OPEN,
            carryin => n12078,
            carryout => n12079,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i7_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52306\,
            in2 => \N__46300\,
            in3 => \N__46288\,
            lcout => duty_7,
            ltout => OPEN,
            carryin => n12079,
            carryout => n12080,
            clk => \N__56072\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i8_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52281\,
            in2 => \N__46285\,
            in3 => \N__46270\,
            lcout => duty_8,
            ltout => OPEN,
            carryin => \bfn_14_27_0_\,
            carryout => n12081,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i9_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52252\,
            in2 => \N__46267\,
            in3 => \N__46252\,
            lcout => duty_9,
            ltout => OPEN,
            carryin => n12081,
            carryout => n12082,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i10_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52701\,
            in2 => \N__46249\,
            in3 => \N__46216\,
            lcout => duty_10,
            ltout => OPEN,
            carryin => n12082,
            carryout => n12083,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i11_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52675\,
            in2 => \N__46213\,
            in3 => \N__46174\,
            lcout => duty_11,
            ltout => OPEN,
            carryin => n12083,
            carryout => n12084,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i12_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46171\,
            in2 => \N__52651\,
            in3 => \N__46159\,
            lcout => duty_12,
            ltout => OPEN,
            carryin => n12084,
            carryout => n12085,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i13_LC_14_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52617\,
            in2 => \N__46156\,
            in3 => \N__46144\,
            lcout => duty_13,
            ltout => OPEN,
            carryin => n12085,
            carryout => n12086,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i14_LC_14_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52591\,
            in2 => \N__46456\,
            in3 => \N__46444\,
            lcout => duty_14,
            ltout => OPEN,
            carryin => n12086,
            carryout => n12087,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i15_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46441\,
            in2 => \N__52558\,
            in3 => \N__46429\,
            lcout => duty_15,
            ltout => OPEN,
            carryin => n12087,
            carryout => n12088,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i16_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52531\,
            in2 => \N__46426\,
            in3 => \N__46414\,
            lcout => duty_16,
            ltout => OPEN,
            carryin => \bfn_14_28_0_\,
            carryout => n12089,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i17_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46411\,
            in2 => \N__52507\,
            in3 => \N__46402\,
            lcout => duty_17,
            ltout => OPEN,
            carryin => n12089,
            carryout => n12090,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i18_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46399\,
            in2 => \N__55396\,
            in3 => \N__46390\,
            lcout => duty_18,
            ltout => OPEN,
            carryin => n12090,
            carryout => n12091,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i19_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46387\,
            in2 => \N__55366\,
            in3 => \N__46375\,
            lcout => duty_19,
            ltout => OPEN,
            carryin => n12091,
            carryout => n12092,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i20_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46372\,
            in2 => \N__55333\,
            in3 => \N__46363\,
            lcout => duty_20,
            ltout => OPEN,
            carryin => n12092,
            carryout => n12093,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i21_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46360\,
            in2 => \N__55306\,
            in3 => \N__46324\,
            lcout => duty_21,
            ltout => OPEN,
            carryin => n12093,
            carryout => n12094,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i22_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46621\,
            in2 => \N__55276\,
            in3 => \N__46609\,
            lcout => duty_22,
            ltout => OPEN,
            carryin => n12094,
            carryout => n12095,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i23_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52918\,
            in1 => \N__46606\,
            in2 => \_gnd_net_\,
            in3 => \N__46597\,
            lcout => duty_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i13_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55652\,
            in1 => \N__46504\,
            in2 => \_gnd_net_\,
            in3 => \N__46594\,
            lcout => pwm_setpoint_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i16_1_lut_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46584\,
            lcout => n10_adj_576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i14_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55653\,
            in1 => \N__46564\,
            in2 => \_gnd_net_\,
            in3 => \N__46549\,
            lcout => pwm_setpoint_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i4_4_lut_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__46543\,
            in1 => \N__50128\,
            in2 => \N__46528\,
            in3 => \N__46462\,
            lcout => n4_adj_605,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i10_1_lut_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52788\,
            lcout => n16_adj_582,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i14_1_lut_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46503\,
            lcout => n12_adj_578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i0_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55651\,
            in1 => \N__46483\,
            in2 => \_gnd_net_\,
            in3 => \N__46477\,
            lcout => pwm_setpoint_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56083\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i13_1_lut_LC_14_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46791\,
            lcout => n13_adj_579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i29_2_lut_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46677\,
            lcout => n29_adj_622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i27_2_lut_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46695\,
            in2 => \_gnd_net_\,
            in3 => \N__46743\,
            lcout => n27_adj_621,
            ltout => \n27_adj_621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12368_3_lut_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__46696\,
            in1 => \_gnd_net_\,
            in2 => \N__46687\,
            in3 => \N__46684\,
            lcout => OPEN,
            ltout => \n14840_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12369_3_lut_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__46678\,
            in1 => \_gnd_net_\,
            in2 => \N__46669\,
            in3 => \N__47171\,
            lcout => n14841,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i23_1_lut_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46665\,
            lcout => n3_adj_569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i17_1_lut_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n9_adj_575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i16_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__55654\,
            in1 => \N__46639\,
            in2 => \_gnd_net_\,
            in3 => \N__46627\,
            lcout => pwm_setpoint_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56087\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i21_1_lut_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47061\,
            lcout => n5_adj_571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12250_2_lut_4_lut_LC_14_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__46842\,
            in1 => \N__46859\,
            in2 => \N__47038\,
            in3 => \N__46926\,
            lcout => OPEN,
            ltout => \n14722_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12404_4_lut_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__47005\,
            in1 => \N__46886\,
            in2 => \N__46993\,
            in3 => \N__46867\,
            lcout => OPEN,
            ltout => \n14876_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12414_4_lut_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__46887\,
            in1 => \N__47158\,
            in2 => \N__46990\,
            in3 => \N__46963\,
            lcout => n14886,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12309_3_lut_LC_14_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47210\,
            in1 => \N__46981\,
            in2 => \_gnd_net_\,
            in3 => \N__46969\,
            lcout => n14781,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i7_LC_14_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55694\,
            in1 => \N__46957\,
            in2 => \_gnd_net_\,
            in3 => \N__46947\,
            lcout => pwm_setpoint_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56091\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i12_3_lut_3_lut_LC_14_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__46840\,
            in1 => \N__46860\,
            in2 => \_gnd_net_\,
            in3 => \N__46922\,
            lcout => OPEN,
            ltout => \n12_adj_611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i30_3_lut_LC_14_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46906\,
            in2 => \N__46894\,
            in3 => \N__46885\,
            lcout => n30_adj_623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_275_i33_2_lut_LC_14_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46841\,
            lcout => n33_adj_625,
            ltout => \n33_adj_625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12252_4_lut_LC_14_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__47211\,
            in1 => \N__47194\,
            in2 => \N__47182\,
            in3 => \N__47178\,
            lcout => n14724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i18_1_lut_LC_14_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47148\,
            lcout => n8_adj_574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_162_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__50535\,
            in1 => \N__50220\,
            in2 => \N__50572\,
            in3 => \N__50601\,
            lcout => n28_adj_597,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__50649\,
            in1 => \N__50745\,
            in2 => \N__50716\,
            in3 => \N__50586\,
            lcout => n31_adj_594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_3_lut_adj_163_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__50661\,
            in1 => \N__47125\,
            in2 => \_gnd_net_\,
            in3 => \N__50730\,
            lcout => OPEN,
            ltout => \n32_adj_593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12759_4_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47119\,
            in1 => \N__47077\,
            in2 => \N__47113\,
            in3 => \N__47071\,
            lcout => n4856,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1910_3_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48316\,
            in2 => \N__48336\,
            in3 => \N__49324\,
            lcout => n2910,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50616\,
            in1 => \N__50520\,
            in2 => \N__50635\,
            in3 => \N__50760\,
            lcout => n30_adj_595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50679\,
            in1 => \N__50775\,
            in2 => \N__50698\,
            in3 => \N__50550\,
            lcout => n29_adj_596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1865_3_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47695\,
            in1 => \N__47682\,
            in2 => \_gnd_net_\,
            in3 => \N__47616\,
            lcout => n2833,
            ltout => \n2833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10041_4_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__47921\,
            in1 => \N__47256\,
            in2 => \N__47473\,
            in3 => \N__47951\,
            lcout => n11756,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1931_3_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__47952\,
            in1 => \_gnd_net_\,
            in2 => \N__49340\,
            in3 => \N__47935\,
            lcout => n2931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1932_3_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47982\,
            in2 => \N__47968\,
            in3 => \N__49298\,
            lcout => n2932,
            ltout => \n2932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9947_3_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47434\,
            in2 => \N__47410\,
            in3 => \N__47396\,
            lcout => n11662,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1930_3_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47922\,
            in1 => \_gnd_net_\,
            in2 => \N__47905\,
            in3 => \N__49302\,
            lcout => n2930,
            ltout => \n2930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_40_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__47333\,
            in1 => \N__47303\,
            in2 => \N__47284\,
            in3 => \N__47281\,
            lcout => n13417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_2_lut_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47249\,
            in2 => \_gnd_net_\,
            in3 => \N__47215\,
            lcout => n2901,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => n12411,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_3_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54610\,
            in2 => \N__47983\,
            in3 => \N__47959\,
            lcout => n2900,
            ltout => OPEN,
            carryin => n12411,
            carryout => n12412,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_4_lut_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47956\,
            in3 => \N__47929\,
            lcout => n2899,
            ltout => OPEN,
            carryin => n12412,
            carryout => n12413,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_5_lut_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54611\,
            in2 => \N__47926\,
            in3 => \N__47896\,
            lcout => n2898,
            ltout => OPEN,
            carryin => n12413,
            carryout => n12414,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_6_lut_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47893\,
            in3 => \N__47857\,
            lcout => n2897,
            ltout => OPEN,
            carryin => n12414,
            carryout => n12415,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_7_lut_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47854\,
            in3 => \N__47818\,
            lcout => n2896,
            ltout => OPEN,
            carryin => n12415,
            carryout => n12416,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_8_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54613\,
            in2 => \N__47815\,
            in3 => \N__47785\,
            lcout => n2895,
            ltout => OPEN,
            carryin => n12416,
            carryout => n12417,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_9_lut_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54612\,
            in2 => \N__47781\,
            in3 => \N__47740\,
            lcout => n2894,
            ltout => OPEN,
            carryin => n12417,
            carryout => n12418,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_10_lut_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55233\,
            in2 => \N__47737\,
            in3 => \N__47698\,
            lcout => n2893,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => n12419,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_11_lut_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54614\,
            in2 => \N__48304\,
            in3 => \N__48280\,
            lcout => n2892,
            ltout => OPEN,
            carryin => n12419,
            carryout => n12420,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_12_lut_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55234\,
            in2 => \N__48277\,
            in3 => \N__48238\,
            lcout => n2891,
            ltout => OPEN,
            carryin => n12420,
            carryout => n12421,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_13_lut_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54615\,
            in2 => \N__48235\,
            in3 => \N__48193\,
            lcout => n2890,
            ltout => OPEN,
            carryin => n12421,
            carryout => n12422,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_14_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55235\,
            in2 => \N__48190\,
            in3 => \N__48145\,
            lcout => n2889,
            ltout => OPEN,
            carryin => n12422,
            carryout => n12423,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_15_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54616\,
            in2 => \N__48142\,
            in3 => \N__48103\,
            lcout => n2888,
            ltout => OPEN,
            carryin => n12423,
            carryout => n12424,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_16_lut_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55236\,
            in2 => \N__48099\,
            in3 => \N__48052\,
            lcout => n2887,
            ltout => OPEN,
            carryin => n12424,
            carryout => n12425,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_17_lut_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54617\,
            in2 => \N__48049\,
            in3 => \N__48010\,
            lcout => n2886,
            ltout => OPEN,
            carryin => n12425,
            carryout => n12426,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_18_lut_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48007\,
            in2 => \N__54980\,
            in3 => \N__48592\,
            lcout => n2885,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => n12427,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_19_lut_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48589\,
            in2 => \N__54984\,
            in3 => \N__48556\,
            lcout => n2884,
            ltout => OPEN,
            carryin => n12427,
            carryout => n12428,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_20_lut_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48552\,
            in2 => \N__54981\,
            in3 => \N__48508\,
            lcout => n2883,
            ltout => OPEN,
            carryin => n12428,
            carryout => n12429,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_21_lut_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48505\,
            in2 => \N__54985\,
            in3 => \N__48472\,
            lcout => n2882,
            ltout => OPEN,
            carryin => n12429,
            carryout => n12430,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_22_lut_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48465\,
            in2 => \N__54982\,
            in3 => \N__48433\,
            lcout => n2881,
            ltout => OPEN,
            carryin => n12430,
            carryout => n12431,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_23_lut_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48430\,
            in2 => \N__54986\,
            in3 => \N__48388\,
            lcout => n2880,
            ltout => OPEN,
            carryin => n12431,
            carryout => n12432,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_24_lut_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48385\,
            in2 => \N__54983\,
            in3 => \N__48340\,
            lcout => n2879,
            ltout => OPEN,
            carryin => n12432,
            carryout => n12433,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_25_lut_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48337\,
            in2 => \N__54987\,
            in3 => \N__48307\,
            lcout => n2878,
            ltout => OPEN,
            carryin => n12433,
            carryout => n12434,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_26_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48907\,
            in2 => \N__54992\,
            in3 => \N__48868\,
            lcout => n2877,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => n12435,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_27_lut_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48865\,
            in2 => \N__54993\,
            in3 => \N__48811\,
            lcout => n2876,
            ltout => OPEN,
            carryin => n12435,
            carryout => n12436,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_28_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54668\,
            in2 => \N__48805\,
            in3 => \N__48808\,
            lcout => n2875,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1907_3_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__48804\,
            in1 => \_gnd_net_\,
            in2 => \N__48775\,
            in3 => \N__49372\,
            lcout => n2907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_128_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__48742\,
            in1 => \N__49616\,
            in2 => \N__48718\,
            in3 => \N__48706\,
            lcout => OPEN,
            ltout => \n13822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_130_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__49617\,
            in1 => \N__48700\,
            in2 => \N__48685\,
            in3 => \N__48681\,
            lcout => OPEN,
            ltout => \n13834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_134_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48661\,
            in1 => \N__49477\,
            in2 => \N__48655\,
            in3 => \N__49672\,
            lcout => n13842,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2193_3_lut_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48643\,
            in2 => \N__48616\,
            in3 => \N__49613\,
            lcout => OPEN,
            ltout => \n27_adj_709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_129_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__49615\,
            in1 => \N__49705\,
            in2 => \N__49693\,
            in3 => \N__49690\,
            lcout => n13830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2196_3_lut_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49666\,
            in2 => \N__49657\,
            in3 => \N__49614\,
            lcout => n21_adj_706,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2046_3_lut_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__49471\,
            in1 => \_gnd_net_\,
            in2 => \N__49447\,
            in3 => \N__49077\,
            lcout => n3110,
            ltout => \n3110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2113_3_lut_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50097\,
            in1 => \_gnd_net_\,
            in2 => \N__49432\,
            in3 => \N__52153\,
            lcout => n3209,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2130_3_lut_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50788\,
            in2 => \N__50824\,
            in3 => \N__50095\,
            lcout => n3226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12449_1_lut_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49373\,
            lcout => n14921,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2044_3_lut_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49189\,
            in2 => \N__49162\,
            in3 => \N__49078\,
            lcout => n3108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_new_i0_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49153\,
            lcout => \quad_counter0.b_new_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2050_3_lut_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49129\,
            in2 => \N__49096\,
            in3 => \N__49076\,
            lcout => n3114,
            ltout => \n3114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2117_3_lut_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50096\,
            in1 => \_gnd_net_\,
            in2 => \N__49933\,
            in3 => \N__51649\,
            lcout => n3213,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_158_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51875\,
            in2 => \_gnd_net_\,
            in3 => \N__52406\,
            lcout => OPEN,
            ltout => \n7_adj_712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__52352\,
            in1 => \N__52325\,
            in2 => \N__49900\,
            in3 => \N__49897\,
            lcout => n13676,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_3_lut_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__52376\,
            in1 => \N__52433\,
            in2 => \_gnd_net_\,
            in3 => \N__52466\,
            lcout => n8_adj_711,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_I_0_63_2_lut_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50316\,
            in2 => \_gnd_net_\,
            in3 => \N__50376\,
            lcout => \quad_counter0.direction_N_530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__52694\,
            in1 => \N__52244\,
            in2 => \N__52280\,
            in3 => \N__49723\,
            lcout => OPEN,
            ltout => \n10_adj_714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_159_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__55352\,
            in1 => \N__52301\,
            in2 => \N__49717\,
            in3 => \N__52670\,
            lcout => OPEN,
            ltout => \n16_adj_702_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52640\,
            in1 => \N__55295\,
            in2 => \N__49714\,
            in3 => \N__49711\,
            lcout => n22_adj_699,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_161_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52493\,
            in1 => \N__55382\,
            in2 => \N__52586\,
            in3 => \N__52550\,
            lcout => n19_adj_701,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_new_i1_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50469\,
            lcout => \quad_counter0.b_new_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i2_1_lut_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50154\,
            lcout => n24_adj_590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i4_1_lut_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50190\,
            lcout => n22_adj_588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__55325\,
            in1 => \N__52526\,
            in2 => \N__52621\,
            in3 => \N__55268\,
            lcout => OPEN,
            ltout => \n21_adj_700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12460_4_lut_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__52913\,
            in1 => \N__52865\,
            in2 => \N__50164\,
            in3 => \N__50161\,
            lcout => n4890,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i1_LC_15_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50155\,
            in1 => \N__50137\,
            in2 => \_gnd_net_\,
            in3 => \N__55644\,
            lcout => pwm_setpoint_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56084\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12421_4_lut_LC_15_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__50333\,
            in1 => \N__50483\,
            in2 => \N__50317\,
            in3 => \N__50465\,
            lcout => \quad_counter0.a_prev_N_537\,
            ltout => \quad_counter0.a_prev_N_537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_52_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__50484\,
            in1 => \N__50372\,
            in2 => \N__50122\,
            in3 => \N__50449\,
            lcout => b_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_I_0_65_2_lut_LC_15_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50482\,
            in2 => \_gnd_net_\,
            in3 => \N__50371\,
            lcout => OPEN,
            ltout => \quad_counter0.direction_N_534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.debounce_cnt_I_0_4_lut_LC_15_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011000000000"
        )
    port map (
            in0 => \N__50309\,
            in1 => \N__50493\,
            in2 => \N__50506\,
            in3 => \N__50447\,
            lcout => \direction_N_531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_prev_51_LC_15_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__50448\,
            in1 => \N__50503\,
            in2 => \N__50497\,
            in3 => \N__50310\,
            lcout => \quad_counter0.a_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.debounce_cnt_50_LC_15_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__50485\,
            in1 => \N__50314\,
            in2 => \N__50470\,
            in3 => \N__50334\,
            lcout => \quad_counter0.debounce_cnt\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.direction_57_LC_15_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110100101000"
        )
    port map (
            in0 => \N__50393\,
            in1 => \N__50315\,
            in2 => \N__50377\,
            in3 => \N__50347\,
            lcout => n1185,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_new_i1_LC_15_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50341\,
            lcout => a_new_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i20_1_lut_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50277\,
            lcout => n6_adj_572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i19_1_lut_LC_15_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50250\,
            lcout => n7_adj_573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sweep_counter_631_632__i1_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50221\,
            in2 => \_gnd_net_\,
            in3 => \N__50209\,
            lcout => sweep_counter_0,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => n12606,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i2_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50650\,
            in2 => \_gnd_net_\,
            in3 => \N__50638\,
            lcout => sweep_counter_1,
            ltout => OPEN,
            carryin => n12606,
            carryout => n12607,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i3_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50634\,
            in2 => \_gnd_net_\,
            in3 => \N__50620\,
            lcout => sweep_counter_2,
            ltout => OPEN,
            carryin => n12607,
            carryout => n12608,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i4_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50617\,
            in2 => \_gnd_net_\,
            in3 => \N__50605\,
            lcout => sweep_counter_3,
            ltout => OPEN,
            carryin => n12608,
            carryout => n12609,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i5_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50602\,
            in2 => \_gnd_net_\,
            in3 => \N__50590\,
            lcout => sweep_counter_4,
            ltout => OPEN,
            carryin => n12609,
            carryout => n12610,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i6_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50587\,
            in2 => \_gnd_net_\,
            in3 => \N__50575\,
            lcout => sweep_counter_5,
            ltout => OPEN,
            carryin => n12610,
            carryout => n12611,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i7_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50571\,
            in2 => \_gnd_net_\,
            in3 => \N__50554\,
            lcout => sweep_counter_6,
            ltout => OPEN,
            carryin => n12611,
            carryout => n12612,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i8_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50551\,
            in2 => \_gnd_net_\,
            in3 => \N__50539\,
            lcout => sweep_counter_7,
            ltout => OPEN,
            carryin => n12612,
            carryout => n12613,
            clk => \N__56050\,
            ce => 'H',
            sr => \N__52882\
        );

    \sweep_counter_631_632__i9_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50536\,
            in2 => \_gnd_net_\,
            in3 => \N__50524\,
            lcout => sweep_counter_8,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => n12614,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i10_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50521\,
            in2 => \_gnd_net_\,
            in3 => \N__50509\,
            lcout => sweep_counter_9,
            ltout => OPEN,
            carryin => n12614,
            carryout => n12615,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i11_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50776\,
            in2 => \_gnd_net_\,
            in3 => \N__50764\,
            lcout => sweep_counter_10,
            ltout => OPEN,
            carryin => n12615,
            carryout => n12616,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i12_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50761\,
            in2 => \_gnd_net_\,
            in3 => \N__50749\,
            lcout => sweep_counter_11,
            ltout => OPEN,
            carryin => n12616,
            carryout => n12617,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i13_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50746\,
            in2 => \_gnd_net_\,
            in3 => \N__50734\,
            lcout => sweep_counter_12,
            ltout => OPEN,
            carryin => n12617,
            carryout => n12618,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i14_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50731\,
            in2 => \_gnd_net_\,
            in3 => \N__50719\,
            lcout => sweep_counter_13,
            ltout => OPEN,
            carryin => n12618,
            carryout => n12619,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i15_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50715\,
            in2 => \_gnd_net_\,
            in3 => \N__50701\,
            lcout => sweep_counter_14,
            ltout => OPEN,
            carryin => n12619,
            carryout => n12620,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i16_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50697\,
            in2 => \_gnd_net_\,
            in3 => \N__50683\,
            lcout => sweep_counter_15,
            ltout => OPEN,
            carryin => n12620,
            carryout => n12621,
            clk => \N__56052\,
            ce => 'H',
            sr => \N__52869\
        );

    \sweep_counter_631_632__i17_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50680\,
            in2 => \_gnd_net_\,
            in3 => \N__50668\,
            lcout => sweep_counter_16,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => n12622,
            clk => \N__56056\,
            ce => 'H',
            sr => \N__52883\
        );

    \sweep_counter_631_632__i18_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50662\,
            in2 => \_gnd_net_\,
            in3 => \N__50665\,
            lcout => sweep_counter_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56056\,
            ce => 'H',
            sr => \N__52883\
        );

    \encoder0_position_31__I_0_add_2106_2_lut_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51180\,
            in2 => \_gnd_net_\,
            in3 => \N__51121\,
            lcout => n3201,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => n12492,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_3_lut_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54343\,
            in2 => \N__51118\,
            in3 => \N__51079\,
            lcout => n3200,
            ltout => OPEN,
            carryin => n12492,
            carryout => n12493,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_4_lut_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51076\,
            in3 => \N__51022\,
            lcout => n3199,
            ltout => OPEN,
            carryin => n12493,
            carryout => n12494,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_5_lut_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54344\,
            in2 => \N__51019\,
            in3 => \N__50986\,
            lcout => n3198,
            ltout => OPEN,
            carryin => n12494,
            carryout => n12495,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_6_lut_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__50983\,
            in3 => \N__50932\,
            lcout => n3197,
            ltout => OPEN,
            carryin => n12495,
            carryout => n12496,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_7_lut_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50924\,
            in2 => \_gnd_net_\,
            in3 => \N__50881\,
            lcout => n3196,
            ltout => OPEN,
            carryin => n12496,
            carryout => n12497,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_8_lut_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54346\,
            in2 => \N__50878\,
            in3 => \N__50827\,
            lcout => n3195,
            ltout => OPEN,
            carryin => n12497,
            carryout => n12498,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_9_lut_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54345\,
            in2 => \N__50820\,
            in3 => \N__50779\,
            lcout => n3194,
            ltout => OPEN,
            carryin => n12498,
            carryout => n12499,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_10_lut_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54784\,
            in2 => \N__51555\,
            in3 => \N__51502\,
            lcout => n3193,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => n12500,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_11_lut_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51499\,
            in2 => \N__55076\,
            in3 => \N__51451\,
            lcout => n3192,
            ltout => OPEN,
            carryin => n12500,
            carryout => n12501,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_12_lut_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51448\,
            in2 => \N__55122\,
            in3 => \N__51409\,
            lcout => n3191,
            ltout => OPEN,
            carryin => n12501,
            carryout => n12502,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_13_lut_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51405\,
            in2 => \N__55077\,
            in3 => \N__51352\,
            lcout => n3190,
            ltout => OPEN,
            carryin => n12502,
            carryout => n12503,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_14_lut_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51349\,
            in2 => \N__55123\,
            in3 => \N__51313\,
            lcout => n3189,
            ltout => OPEN,
            carryin => n12503,
            carryout => n12504,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_15_lut_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51309\,
            in2 => \N__55078\,
            in3 => \N__51277\,
            lcout => n3188,
            ltout => OPEN,
            carryin => n12504,
            carryout => n12505,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_16_lut_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51274\,
            in2 => \N__55124\,
            in3 => \N__51226\,
            lcout => n3187,
            ltout => OPEN,
            carryin => n12505,
            carryout => n12506,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_17_lut_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51223\,
            in2 => \N__55079\,
            in3 => \N__51184\,
            lcout => n3186,
            ltout => OPEN,
            carryin => n12506,
            carryout => n12507,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_18_lut_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51856\,
            in2 => \N__55080\,
            in3 => \N__51808\,
            lcout => n3185,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => n12508,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_19_lut_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51804\,
            in2 => \N__55125\,
            in3 => \N__51760\,
            lcout => n3184,
            ltout => OPEN,
            carryin => n12508,
            carryout => n12509,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_20_lut_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51757\,
            in2 => \N__55081\,
            in3 => \N__51718\,
            lcout => n3183,
            ltout => OPEN,
            carryin => n12509,
            carryout => n12510,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_21_lut_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51711\,
            in2 => \N__55126\,
            in3 => \N__51673\,
            lcout => n3182,
            ltout => OPEN,
            carryin => n12510,
            carryout => n12511,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_22_lut_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51663\,
            in2 => \N__55082\,
            in3 => \N__51643\,
            lcout => n3181,
            ltout => OPEN,
            carryin => n12511,
            carryout => n12512,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_23_lut_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51640\,
            in2 => \N__55127\,
            in3 => \N__51595\,
            lcout => n3180,
            ltout => OPEN,
            carryin => n12512,
            carryout => n12513,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_24_lut_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51592\,
            in2 => \N__55083\,
            in3 => \N__51559\,
            lcout => n3179,
            ltout => OPEN,
            carryin => n12513,
            carryout => n12514,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_25_lut_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52225\,
            in2 => \N__55128\,
            in3 => \N__52177\,
            lcout => n3178,
            ltout => OPEN,
            carryin => n12514,
            carryout => n12515,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_26_lut_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52167\,
            in2 => \N__55129\,
            in3 => \N__52147\,
            lcout => n3177,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => n12516,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_27_lut_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52144\,
            in2 => \N__55084\,
            in3 => \N__52096\,
            lcout => n3176,
            ltout => OPEN,
            carryin => n12516,
            carryout => n12517,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_28_lut_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52077\,
            in2 => \N__55130\,
            in3 => \N__52048\,
            lcout => n3175,
            ltout => OPEN,
            carryin => n12517,
            carryout => n12518,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_29_lut_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52045\,
            in2 => \N__55085\,
            in3 => \N__52003\,
            lcout => n3174,
            ltout => OPEN,
            carryin => n12518,
            carryout => n12519,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_30_lut_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52000\,
            in2 => \N__55131\,
            in3 => \N__51955\,
            lcout => n3173,
            ltout => OPEN,
            carryin => n12519,
            carryout => n12520,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_31_lut_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54815\,
            in1 => \N__51952\,
            in2 => \N__51937\,
            in3 => \N__51913\,
            lcout => n3204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_630__i0_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51879\,
            in2 => \_gnd_net_\,
            in3 => \N__51859\,
            lcout => encoder0_position_target_0,
            ltout => OPEN,
            carryin => \bfn_16_26_0_\,
            carryout => n12663,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i1_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52470\,
            in2 => \N__55086\,
            in3 => \N__52450\,
            lcout => encoder0_position_target_1,
            ltout => OPEN,
            carryin => n12663,
            carryout => n12664,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i2_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54819\,
            in2 => \N__52443\,
            in3 => \N__52417\,
            lcout => encoder0_position_target_2,
            ltout => OPEN,
            carryin => n12664,
            carryout => n12665,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i3_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52410\,
            in2 => \N__55087\,
            in3 => \N__52390\,
            lcout => encoder0_position_target_3,
            ltout => OPEN,
            carryin => n12665,
            carryout => n12666,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i4_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54823\,
            in2 => \N__52386\,
            in3 => \N__52360\,
            lcout => encoder0_position_target_4,
            ltout => OPEN,
            carryin => n12666,
            carryout => n12667,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i5_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52356\,
            in2 => \N__55088\,
            in3 => \N__52336\,
            lcout => encoder0_position_target_5,
            ltout => OPEN,
            carryin => n12667,
            carryout => n12668,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i6_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54827\,
            in2 => \N__52333\,
            in3 => \N__52309\,
            lcout => encoder0_position_target_6,
            ltout => OPEN,
            carryin => n12668,
            carryout => n12669,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i7_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52305\,
            in2 => \N__55089\,
            in3 => \N__52285\,
            lcout => encoder0_position_target_7,
            ltout => OPEN,
            carryin => n12669,
            carryout => n12670,
            clk => \N__56080\,
            ce => \N__52896\,
            sr => \N__52827\
        );

    \encoder0_position_target_630__i8_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55102\,
            in2 => \N__52282\,
            in3 => \N__52255\,
            lcout => encoder0_position_target_8,
            ltout => OPEN,
            carryin => \bfn_16_27_0_\,
            carryout => n12671,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i9_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52248\,
            in2 => \N__55213\,
            in3 => \N__52228\,
            lcout => encoder0_position_target_9,
            ltout => OPEN,
            carryin => n12671,
            carryout => n12672,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i10_LC_16_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55090\,
            in2 => \N__52702\,
            in3 => \N__52678\,
            lcout => encoder0_position_target_10,
            ltout => OPEN,
            carryin => n12672,
            carryout => n12673,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i11_LC_16_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52674\,
            in2 => \N__55210\,
            in3 => \N__52654\,
            lcout => encoder0_position_target_11,
            ltout => OPEN,
            carryin => n12673,
            carryout => n12674,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i12_LC_16_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55094\,
            in2 => \N__52650\,
            in3 => \N__52624\,
            lcout => encoder0_position_target_12,
            ltout => OPEN,
            carryin => n12674,
            carryout => n12675,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i13_LC_16_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52616\,
            in2 => \N__55211\,
            in3 => \N__52594\,
            lcout => encoder0_position_target_13,
            ltout => OPEN,
            carryin => n12675,
            carryout => n12676,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i14_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55098\,
            in2 => \N__52590\,
            in3 => \N__52561\,
            lcout => encoder0_position_target_14,
            ltout => OPEN,
            carryin => n12676,
            carryout => n12677,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i15_LC_16_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52554\,
            in2 => \N__55212\,
            in3 => \N__52534\,
            lcout => encoder0_position_target_15,
            ltout => OPEN,
            carryin => n12677,
            carryout => n12678,
            clk => \N__56085\,
            ce => \N__52897\,
            sr => \N__52828\
        );

    \encoder0_position_target_630__i16_LC_16_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52530\,
            in2 => \N__55214\,
            in3 => \N__52510\,
            lcout => encoder0_position_target_16,
            ltout => OPEN,
            carryin => \bfn_16_28_0_\,
            carryout => n12679,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \encoder0_position_target_630__i17_LC_16_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55109\,
            in2 => \N__52503\,
            in3 => \N__52477\,
            lcout => encoder0_position_target_17,
            ltout => OPEN,
            carryin => n12679,
            carryout => n12680,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \encoder0_position_target_630__i18_LC_16_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55392\,
            in2 => \N__55215\,
            in3 => \N__55369\,
            lcout => encoder0_position_target_18,
            ltout => OPEN,
            carryin => n12680,
            carryout => n12681,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \encoder0_position_target_630__i19_LC_16_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55113\,
            in2 => \N__55362\,
            in3 => \N__55336\,
            lcout => encoder0_position_target_19,
            ltout => OPEN,
            carryin => n12681,
            carryout => n12682,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \encoder0_position_target_630__i20_LC_16_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55329\,
            in2 => \N__55216\,
            in3 => \N__55309\,
            lcout => encoder0_position_target_20,
            ltout => OPEN,
            carryin => n12682,
            carryout => n12683,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \encoder0_position_target_630__i21_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55117\,
            in2 => \N__55305\,
            in3 => \N__55279\,
            lcout => encoder0_position_target_21,
            ltout => OPEN,
            carryin => n12683,
            carryout => n12684,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \encoder0_position_target_630__i22_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55272\,
            in2 => \N__55217\,
            in3 => \N__55252\,
            lcout => encoder0_position_target_22,
            ltout => OPEN,
            carryin => n12684,
            carryout => n12685,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \encoder0_position_target_630__i23_LC_16_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__52917\,
            in1 => \N__55121\,
            in2 => \_gnd_net_\,
            in3 => \N__52921\,
            lcout => encoder0_position_target_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56089\,
            ce => \N__52881\,
            sr => \N__52823\
        );

    \pwm_setpoint_i9_LC_16_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55706\,
            in1 => \N__52801\,
            in2 => \_gnd_net_\,
            in3 => \N__52792\,
            lcout => pwm_setpoint_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i9_1_lut_LC_16_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52731\,
            lcout => n17_adj_583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i1_LC_16_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56382\,
            lcout => commutation_state_prev_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dir_151_LC_16_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55707\,
            lcout => dir,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2137_1_lut_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55695\,
            lcout => \pwm_setpoint_23__N_195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_inv_0_i7_1_lut_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55546\,
            lcout => n19_adj_551,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3168_2_lut_LC_17_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55887\,
            in2 => \_gnd_net_\,
            in3 => \N__55516\,
            lcout => n4886,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12416_4_lut_LC_17_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100010011"
        )
    port map (
            in0 => \N__56374\,
            in1 => \N__55515\,
            in2 => \N__56180\,
            in3 => \N__55471\,
            lcout => n4842,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GLC_165_LC_17_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000101100"
        )
    port map (
            in0 => \N__56301\,
            in1 => \N__56165\,
            in2 => \N__56434\,
            in3 => \N__56375\,
            lcout => \INLC_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56095\,
            ce => \N__55900\,
            sr => \N__55855\
        );

    \GLA_161_LC_18_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100000000011"
        )
    port map (
            in0 => \N__56296\,
            in1 => \N__56376\,
            in2 => \N__56194\,
            in3 => \N__56437\,
            lcout => \INLA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56096\,
            ce => \N__55901\,
            sr => \N__55859\
        );

    \GHB_162_LC_19_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000100001"
        )
    port map (
            in0 => \N__56294\,
            in1 => \N__56389\,
            in2 => \N__56196\,
            in3 => \N__56429\,
            lcout => \GHB\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56097\,
            ce => \N__55912\,
            sr => \N__55864\
        );

    \GHC_164_LC_19_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000110"
        )
    port map (
            in0 => \N__56295\,
            in1 => \N__56390\,
            in2 => \N__56197\,
            in3 => \N__56430\,
            lcout => \GHC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56097\,
            ce => \N__55912\,
            sr => \N__55864\
        );

    \GLB_163_LC_19_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001000100110"
        )
    port map (
            in0 => \N__56391\,
            in1 => \N__56436\,
            in2 => \N__56195\,
            in3 => \N__56300\,
            lcout => \INLB_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56098\,
            ce => \N__55908\,
            sr => \N__55860\
        );

    \GHA_160_LC_19_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101100010"
        )
    port map (
            in0 => \N__56435\,
            in1 => \N__56392\,
            in2 => \N__56302\,
            in3 => \N__56187\,
            lcout => \GHA\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56098\,
            ce => \N__55908\,
            sr => \N__55860\
        );

    \i9555_2_lut_LC_19_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55771\,
            lcout => \INHA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9489_2_lut_LC_20_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55767\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55795\,
            lcout => \INHC_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9488_2_lut_LC_20_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55777\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55766\,
            lcout => \INHB_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
